`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ic+e2vwK5Q7PgjSgvwMH2WoojQ4BbTVuQzxkOMVjPI/VZ5NZbfo+pDZV2xAqhpQmyQ9GvI+HXb1j
HmlK88vB0Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EhYQ5ehP63YE16bz7Bs+Jp6XRtGGK+uBxpAwDXHwR28I2BtSgb9ncXucOpIeu0UTEMLqbvoLfbxU
MKaMrYPMo8RM/a2HDSBr9m9kqrCswhqrsj7+l6YpDAYmcCTq9T3FOkfhQRKFn0OQ/XIIbTvvITnM
Im9Df+3DnhnBsRIa6b8=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h0YJz7QAV8KNys9f0Mxlf+pNNU8LPo3hH7TmUMyrhw3lSO+kM5IGhIhrK6tA/vHS9HjpGQeWP4CV
hUv0PJuDbFRDQozJGwYt7sEJSKD17mUe+oi8D93Qmbv3URq5Gi+VGUtURDK7m9vfm75L8tyy5ql9
qECsNvUIWukIEumtJEY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pP+6eQFqDiaeKP3BC0Vnjvzv+UaX8yu0QFcUAsHG6nA3D6UEozm0SxdJ2iFfFcGPTkGK1rJp3wQa
XKLNY1k0r+8h6/HdEgYrEoLQxiu0rGTrMwFGkm5IpBA5qyUQJ9BOMA3RodmPZroFnpuOiQG9fXXi
E9pTQFAqbQwJUIKn68iPFrjVm+q4qLqQgrHvjKnf6JEciMX/HO234NTOg6COPSv7Uyo3FXOOpRHp
TCTyJBrP+6/0PD1dPLxzogieQ1fECqhCHlBWg5ARc7Wy8Nrvyugiw7tyWe9OCXkF34mphNHjHAfM
kre/l/mYmZh4jzXcx586HHX8Gny5RYaZ4KoAiA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DtRivEEQldRL8LC1umq+yZAExH6mDpzyWG1k5T3n0AafinwOAShYDeN3xJBVTROrx8yaZtcjOIVo
RTz2YCioii4y47KGQkU7qOYGP1IL16aZBaLHN0ikiASZGuT2wIZ7vBOHDkXuyg7SHEzSut20MVdH
yT522lI1hnAfDXEZagb5qrrQxGlsFJtLUxTUFbZ7CLxKt7IYJNSHgoLTaurt9KNyJHnk2Oa9efJx
cG8KJwFEfS1eHTBu0rJX6eoLGEyPSJx4qXZ3eGjOwHDiGelueO/b4BZB7QA7g7zVJz86kqUZqX1s
SpXZOqr7kFUwCnN2dJO5bhUtoF+y3GgfGerZaQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pemFOX3XLyQdy4vtMYjiFXTZP+XlsBGKuE92WyWU4tr/zi/kdVNH1ODTNxNJ5DXwFjsQE3XaQKcO
QVG3dkRqyxkufPvrynU460117JgXGW15a8rem6Dsd8qn7VgNRECRRwFEFLE3bFhFjG5aqlEDnd56
Jtv/dX2cI0okyfMCEOBuMBd48KhjQsDycf7KtJc5LpL06fv+nYIvBQGKfMIkl6F4N9MkpkCF18HN
sm252Xem8SRCkTNQW6+o1yOVN45d9b+5a9+kx3Hc+5oEfCtymCxxbWIPnLnMAGhORy7lTFlrznDF
KTRSVyP9INWg2r5KEz1jo7u/eNIyiLfueJeDjg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
+93ue+0K+V+pjfzqa5MG7PcsuqUtaSJlJ1C3g+5PmNsF0k+K0SWg9dc6HZ3SEW0oUBUAZuZ4NQMC
pwKE7jI1z3e+v2BVU3pviQRu4Lz6ZpHq47DbmsjJdPNuAvCy1lXKhMAl5RUHAAHsTEnDAIcKmUIe
zpCTr6bjbDtmeEybza0diDN9DQV9/JCh0uLlsyyFtykb1pM9XZDildiNJTRP8zqycJ5uYSLDBF39
21yy/chK+5M/3/tLMfmc+tB0LMwnHYAPCoq4kodMpfuNoMhoUiBRch8eOQ+VzntKQ7Z9lOthUbnd
LmP/8OFkzFfeOTg44p0nQ4bYLfoPbMPrp9h4blR+tRklvt8gXwVxAET3VCDwre5pUCp9Y0skYyaJ
F5tjc+frCA5szZBHY1dIhrEAdMFCErWNZzrKRaEmlMjff4Zc52Kk7TdmaH2oX+E5CBLfAorgZrSt
UixYqC+TrDLFCih2Bq3/Ba4K+JqnfbE6C0fGdPfPkDFSanezeQf9vY3TLEEiDtwg8yL8qbZxFXo3
tW/ATQ1Miwn1NLtITQteDtpLohgBo/6S4oICSlW7KdZnruZR35QWSI5CoFlOBqO4yq+K2MADgpS/
8+qPal9KpNccavBukh3kf4bxXkoFp5zLRIlL4DIMlvCO+WW1SAUjdQt/a9agUrdkNSeA+DWgoOft
WeWypClsQXlPAxfzD/TavnizJ4RuSadVZDJA2hxpgBYYYcgt+rXmCnElSHQHnoRo26w1sLNtUtsA
GXxG3C9aXZSEV6opM8YeXGrwZY7+HufHcjGzy9ti2NLlFOSuPGwYqvd/yJ8p63z7O2JOQkjg2M77
N39M6nTpt2WsycjvpTDrcQhSiK0j6t33hzRb8Pw5zJOgnzCPDQwqEysMuk8T5tsiWOkYC4Kb/ceN
Rb/v/eEc0CcsZh6/QgQLz2U0hFBeXK00H/E+FWTnRrUTUbJxuIy9/6LWNwVDROGKJ1TI/YcQPLJc
ND1ZwMm+EtA9/RZecsjy4CDictn4mtwjCoUF42TGiszYBTbHx/9Oi+MTujfsSVBzFnBEqXvrsXl1
fHme0y3mVR4bVZRMf+0AvjpRZ5va0zTH6UhYF+NHq8Dhe7b+XVxlG4XNFtwznlUOd4v2z1QLw8Nq
VqAXC2ReB+eGewr1IdQSGO+2zJsyxdWSYQk1w7VLR/D3i+B3JaKqJAbkLtuOU9fKRWiac5Eu6uRx
uhoWqjuEUDGOuqXjTEgJmsaoQKMCy9hDHZuSa33vcXAYEG2+p9GUxCNcqAD/UOK2od6HBlJoVw6a
YqNkWukJVSWkzig3F0Crq//WA8Ts4UKkh7vh7J6iIDmfAOm6m/pvI7Np8NVE2UD+Ot8l3sVxeURn
0BgpUjUb0zEGsDiuNWaj4J/xOye3EzFHEaQTlZ4erF2usSFQkFq4yrOMddoKKkASRHneiCyaHGY3
Hw4/EsbC83Wb6L/sWu3TOi1e1DV7WHW99nkmh+Jsyaxk9yKy1CB9e15EHgL077WdGQh97gcFFenF
9h2dlNrm2cz+Yzr/HTQ9Hk0md/Vp4xnTZLcM2yf6yQCD51l+hS3TM6PFD7DKBoKLeU3ctcp3Psoy
Fvh6q8EQAGW3YFXab0159QibO5/JiMC8hDwCA0Df2+2w1n14g0dldwsoSs9z2WpxQl4+juLxsGq6
uFKLG+oNJxaN+IaLSdgqJIwPA9YOZcI7jGlkGbuthz5rGBPj47zcGAdoC4OI783kvYDbSODLtneF
yN1pLAJuWHe4cSJVfJGvxNgr9A2UCbM0GiCsjas91qJHj1JKPJWh3xECalex0S94B8UTDfkRGCfm
63E9LKoNb7Uwxg2U2CYeDkB65cN+ugPsGpPuxnV3Q2AOZOqCZDsFJHKDcy5lAU8APQBQjVExUb8T
a4reAxSmUYvxBfSLKehWriM0ZdT1ONlUjAwOt7VFJuxbT74vYF9Vi/Mw7+vy9KZ0jJ29uWSRBrWo
K1UqlmXMm6jvygRVfVHmN6Cz4H5jqvU02YBF17DEhy4gE6xmJrJOx9xCrfnqdF/2QZkJYuUx1o4g
qfX/Fvv+PlcwcnZFeu1kNSyn5auxjjjcrtI6GRiRSE47vZBRCMTWxn7Um+yTduDYPhT3zrclKvXI
+DdshLfKajag/ppQwykcswpcUCF3ZGhmzyFSI5WthzTG801M/wWmg2cGxWcFTw9jjo1Xr5cnc4GO
43IQMv9+qcReubLMVsttcjq0hR1k+wPSHu5rnqc73TpJxCI+SBBI5WCTv8W1WNeQzh6XflcwuzMd
9NGsu8WsSu6WpeWDiE8m282QNCzl+UwULYWuY1zUh3dNXiZr6qvTxKQjfXfGFFOA/z3uvllhDvP/
8vEU5tEFH+1HTq+uSwlSib8Dtgob2lGF2JPSJDVWwAuYT2A6RknHgEXMO2WZFgwVDcJj2+qnCZvV
35IPGw6mFAJ2HnnKGFnoMUeoEuzoUVMIo3lPiKZYtWGgmunoD7f5C62wjzrGCop5tqMJS3OshEjW
W8vmnngblDvHjNJ290dpmNUmnYZ87iMyrrECjBVd0F2D6vVuKdUNaK6mv6THC7GkE+umX4gNk8Qf
SWqpYjEgSalFMbIbgwbo75MTFbrL1fLKH7ne6cyJWh80OXiXQ1D4cbSCvnDtQJQ5f/poD4paaZA0
SR5bBcUrDKalzBgh8LxyK0rkC2pI+0nFsEvRxsLwco89w0cBIDZKmT9Ek5GLD606jwe+zjrDIdxI
z35WQr0WHKcUcSjcgsfGLjR/6YQx8umByifnBECcbTuZ9abgWyfXmUW0bB5MHjBBu8wXum/BwC1J
8kN6X9bNdcXlUkjuwnE+M2cJTpTPVf/V/vuMIUj8dsliqwYa27ksC5etzWjWdK0uw+xuBAFDt5kF
nCwzj7Yyw89YzautEurk8mNi3f0OZbW6n10kGw/7OVvnWJIfB+8Gfq+YHWUOIMCtNhqVbPp0bEja
gW9cKOrZsOznOR8k1HkC8pHlkq3iRRJTq+e5yuZD1iDmp8FELRaFibGmB8hA0WTbwb8GIbnMRVrH
PGgUPho4Eyxa7nq1J+EYb8BI/+dxc4D2GdHH4t14XS9jI8sHnU6aorFlAREvSRzFKybQYS7Lupxh
8ed9YLuAyoLzh3tCWvG1o153Qhi4mi4gT5x6ZH3nO9PLWxX/9JVHlYSUUCfNO0oIVqHHk9KhpSS/
35zjhUhfDl4Eh2cbIoFmfrZ0u4J8qO4M5ap0A1TC0ojdT4IITuykBlJ9zS2rjUAG5jP9yEWo9pHF
qy0mhT73eI/NCyYhYDPiG97oD0Hx22KerLJtYfDtUvZ6AxMBE2mM4kh2abJRxM4xADi6y+n/McNc
x0cDGUhAcLVbt6qujR+PKrbqiDnHU0nGzyRg9zLVZuzhEjhoX21PQTpBfkPIraOnQnUS54RC54GB
RVmIuqZnOBSLG+kfUe86QJLfH55EiZFXMyWuurzGw3leEE3SScPh13PJZ/Tv9C0OqjDHxjc/HSXl
lqhrdrinmgGuz3hYHyk2caEGRAAfXmoAmOFe20Wsuwfwb7q9YoHnfyu34Fek330xKmRa9jUGEUgX
eyU6w67EkJH+IxbcUALMKx8cdXjVAdxfpc72g8UQzZmt8Jk+oPL0nna9RvzGYamwQaLULrEKoKgg
trS3brHErC6I/Bg67DDaRmvrJEV9xFa2B/7jdHc9EIJAA9pbQEGlZ8+l0XJVVC+Z40LxWURgnEzW
eo50E7je8Jf+ZXa6FldlB0BKShYQQIedYeAqC25OcY+IfFQ7TfDUgcUGQWRYRhtpFTQSwnUnMEIH
qSXDNI1HOraveLjYfPYlRYubIs8q55ibymXfj0PtoRHrKvHmreaV+dh/WXfc7IEg5hqtnHDZcqEz
WbHrjMHx+mW89bVolRAwoyNZvnHd0CcrtPb4kGau9w4NmuzAIXBf18kqATWPGsdFV8Gy3zFhj2mL
zOn9aDDU4HFATr30MBEGdKE5DrsPbhMFE2InAi3n/OxNYZtvccPY2hrAGM/HmiByn/TDIvvEZIss
9xBBI2qhdgJSjjWHS4+aRUNeeXmbtKGU3k7CHYbi7oeqePWf/XLGfSlCU1DVZWna9+wbqQKMAFLe
IFuU7eJVIczR09nGQsPKkN7zCDhOSQtZ+xekit0lHyZh15NOnb1n/6y2Bt0MF2NRy2WwWq76dBbu
5aYChbq0+ryAfVOTpnQGrdk6+tIc4Sa0++tOoM6QvfZfgdkwffrEHhealgTpftw/Rr39dPWmlyIP
epqioMdLShBDEoXPcEGaTZz2K1NRLrwk6bcjk3aF3QGriX4Jzi2zUEcQbGbEvopuMVmL567+rgPP
N55SZNtTUxHjJ1fGF44RNAB+1daXzrp0xk9CV4H/XDszNqOe2hwdL/4ywPAJJEErK7NeMhlRZm4+
5or79YPIU4Zne2UWukwnBGy61IqJnYsdkJhqCdo9cvLj+hYG6g47XqobPcuJvyYa8clruBY8b5eo
wAwg4jQ4YfRApjocn9hAkx9ia1pzuveliSOXBXcFXwW4aP+4xrZQFptPOj5QyXRG8kBDmYiR9jWH
2O75XC4AAp5G6kkJAH5cMH/oPuyfiiEysua1+/rjHfMd0ep2LsO7iZp1aSvzaJTvHepE5RUHUFWI
z2QCD+6i7jejV3Np2F23OGMLYLSaPVkQjbFDd3h2vU9IB9fZPYmX1FeDg4yd31nxg9Wjb824O+nr
A+52xW6dVufVnJpzlUF+RPgp9zJaWLjsZ/BPWO+Knrj/l61T3cCGNY91iOHZMG/4wYeYfXOKahjT
qUwETSQIQZKxCU5x9E5EnJHSeICnI+77bIuzEXg5SvIPewawTviodW0GsgXxNrbIEN1bpjSR5w7e
XA2zQsAdNIPEmRmZrizFuZJ2aZ5qLqyPwQ3+u0+Q1J/z9puHMeUON2knHjFXlT12jfz8C6mHwpQu
oJU5GM7fu2M1yNRfBu24PFoO4x9T7KfWOdX+IBk3ykJHVSRNlOe/aPc8GwZGdZ+8/1nAbUqZznu3
Pw2docIu5c1D4qAj/NYgO020RWcgLu5HDAfPUT0YG2ZaRg2rmURibh0Y0aN5UOjIc/X0/Wse/m5K
urbEJrXSr04ZIAKxit1LTIeH34tXtPaLkTid0VuBwvJBGUVsCaIzT4GtuFso3QN+095SQeWbkzD+
j1TDMCcqhXmXJlyjWRwYYITAWzGD9AaGiZA9BKTJikb0S7xFZNX8x6dWMP6T3vlcphSOdenYa5uy
tVijVIQXiAjm5AwBYLMGSVk77KzBeZoer3NOi3bmtO+6izgmDAhqkOziIG1tXcieYYSQ7zD6jXaa
bcxqb2JtQC3KJRbge8ChDPB6Q43rcAGWZo21Vy+wCxFJwV/jdahXsTZq1ODPgoMcidBHVgD19mWc
BANwdfSM18JaKL5e3RQEqffLA6I3cTu2RXThNWdS98WY6/fQyAID3Noi84wzNylzBb8vBhvsoQ1s
olPXbYvr2JeOqD5XOTsq5lQrughsEPUalMWkGGZGJg1RIwI51N/Nu8mFxM+hc7qYzAqPWNrne/qL
SogeCOjady4QlaDBrT3TB9Ow2nyxGRRFQB3+KGTl56FouuiCS81kKWViXHeG0kjgGEk34FRriWgN
HXEEWJLl09jSaxjT4+/gCfjF5pvl0cp0ZOdD3X1WJoO8xSeQbONahzKUyuMxjCqP/1io+xiCCLok
ptoGWAXmcQIPQ2fzPJQ/zcsK4aYc0VLlnpL0qgpeH0KiMLL18awNCvhOc1c57X8ZQL4v/MnNiSnf
dxZsLEeVVaJu++27bXa8y3b5gEhcR4HqXcGtr+lSGNAgLCaqvWctX++8t2Jn0QFd+5u6ODOO69X/
9rxXMSfIWOFXucTZGeYN96imW79sLMjZXhpbUXt7pJYWbTC+cgW+wP3ZAjnUrN/AyYysDiqx8IaY
Hvb68eC70CGWz+Nvy/yF0LVkeChdMcLoNjUN+FimdZzh3PL2sMQGVAesq7RX/+g+m8e2y1aVV+uM
DvrvDxu//rAJt00uIDX0KyKQuesk2Kystx7nIIhGzzW8kYf5ZId86sUjZIE1ieUR4l6RIeKJ4gm5
BW5Bamm6Y0Hy0oiCxNL4/9JXlffCpdjpODYmXMPWATy7SN8EUwgfrEseTShp7g+7Nl++Nh8iVDPj
ui36qtcF7+Is5Xej0qxrX5xo0LTHPSK6Zma+xewpiBTKCw44iGsxDn+3bIlr9pR1HJpFs5IH6cU2
qMDBLdnCylaX/fzDiHOg5FErmyFh9Pru3E4gwy5QEqSqreEoNDzYrOcjVVu1T3gX9i8ODF8cFitB
lzRA+KTHqNCil9iN3JbQ5y+xtNJcD8m77gMOpR+IMX6WTxlJcDye9iYKZ6EmA8bpTo2+FTW73vmw
JiCCBi7xIIJON1jgSpPnvLaG8yxyp/v1wopmmBAsldglfDcBeBTUF837kS29An1v4u3+bnqoeEfg
DA656FJveNNyWn5GXnj3dcxircOYaxOEf7BgEyE89w4wBCQXfkQOcPow6FWI5Xrg5umTv3ODzcFW
KFLbVw49c0cbAnH1kz5MBhDxDIE+aBrjUGv6z4erEXoWn1tIciENMyRA/7WtxA1tTplxI38c9l/K
3+aRTwuYxFMlvEhKr6ndqvqn/o/MY9mM03ZcuAYcek0pegIHupoaowf4toVkBKcvipiD4S7q7Fvf
JmFT4sy9fzXzdPhtAM7uYQxjOs+tT+bNTq+8bbXf3XFnOPmS/7woHvaySwf+A+v5iRnW0gNrwM/L
HF10Xh+NGl/FLLsd1PyyY0YQwQWVpYFYAqkfqXibmZsHutV1zd8vSURSXjcyOIOlanhPc4M9iViU
lHye3oJHoNZQZi2b5Thpb9OAxuQEOO1wi2fKirahqoM6Ymo6a+r8pN1+h2JiN4HKwod4kmjsV98s
eQQ/YJS/EM84AJr8qoACoJChc7iXtXDzRTV7l6Vat1XIDdLme517RroB5fuoaX8JUBmrUoPodq6/
iUZddqISDdr8A1yHhzH6m4rojdh03TRmk9BxtaIICC5SDwFPvUDScPC/NKHu7EFfhBnH0CEBu37Q
GYyhN7/7GJe/oPM=
`protect end_protected
