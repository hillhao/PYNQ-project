`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iX1WH6lCwGPTfoT4q/xNrK1Aj2reaQarfseiUAS/ifZXhEwoB6oE2D6RZAFaF0LKNSam6Ru10gWw
5pLuKoROIQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bARjz+rQAsd4I8CGYLjXNRkBYuWKzzuB9PMbJDCJ04njXAjtXL/+6vyr+nxazh3VyCYSnkr5TJI7
Ve5ZLr6quqhg31JXTykN7hQnYHCd9kyM7r0OxtPDQ1LBVhMXDkYfsb9It5sObCsIyuqLphQn9OPb
TnXAYHH1Blz3OHUzqJg=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uhPlqy3xo1NihYW65X7CDC709m7cEaomoqflzTMuS/8WBbp6sRi4syCpke34NLfAuO5W2qaz0R6K
WEYPH+EiH235nzNLMA8J24xu5dT9joybYah3TPZ0DYhTF75c6itxyHJIMV1xl+556A7yxyTqF8zi
s7XwcSTxQDJDiuMSoCU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Eb4QcmBeu+Cl8swJPx7VDsvjSfEWrnkHhWG4rWRwsc73fhQAQLplR4cWpWgTSreaLZ4C48JupiM9
B2hgDC4DJky8pusJSDf2FgZJphdDMwHLGDGbvr4ojVfULIp5wq91+a0GQnWhNlTKEmY5lBkY/P4n
7kf1Z9mEwremI8vQ2FD1+UlD5xKMI9lLLJVag6NZ1YkXBsVJcDVAo6BFDwhoEk09WbjqU65vcpB7
TL8fY7vF4lLCxbhnxZdd/P8p5EcddQnV5zhwTDPiVunMZ3hX4XFz2AQeYuapAnELVOwngFw/ukl/
7rL9ZrqYTxZjst53Sx3KBWP8KZxhzQUaTCr+vQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CVMWmA316JheGpWyNHL/MR7hELV6yopB7vREjYADDQToPcmx+apIakfQlTn+lUhbK8TYawVFWrMW
8PVl9nMkWkYU6XADi6k34a09IpJNL/zeeeR9RCXkOOAFO6i0pT+HWPb/mM+mAEusd4sZJFgErDAW
5nJsfDAJaDxrOASWGYFYEhQkMoNA7UNtmA6oAGI4jfWX94mAA3Zr5lTvq25xDQ9oyKTdcZCIpiiC
Olb288Irph+QJBryAyW6n8zFiZg9eG8BRH7elDSTqTNXP1pu2v2r6L/uBeSc84gGz+5wZijOYm5p
fh3s11Kcsikk8/7ECM//T89z/v2tqdQKtlsxmA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mTHmFURTiwMZxNH+DQsg+aX9Oa+gLa+goHbf9Wxe/MlyJHwoCuP3Q5v/Q77VpR/j1dlxGRKVGWYa
yxG6QgffcjhepHu/PcrwyyCoKhWjCNM5zi+Ot4+wTUhVBVdEJiP6WaXp4cnaIemA+otZGCMu2sX3
qnsAP9E78Xd/i7bWf42AAREfamnrdHKEIM0h7CWavLUaIZNnqa4lk91Uu7RPd225C5Psd9JD95vP
eu4FnUKLoOlr5PEsChnJwV4j2zhf9hh3PLsVUF/pW0oC6mECK5kHdByNct7cUUWMPn5vvIYimb3+
5AT2S53HD36AKdsgk5tHDf9csmg0fD3RLMSzNw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16112)
`protect data_block
/szp2oV7ktTa9Pb86zLCM0ZDlKzMFirSNU21tttYguylq2VXx/5JCDpUYzpABaSAe40JztxsckAC
RzVWAjri3IKixOxDqXWXhTty87LEJvU+XH2oL73j7S6TgEb+zibk3z1qus+ESRaW4cTF16GdqZ5M
+PjNgj0ecvqiQvEs6g25GmshopXYTEenhsEyqotTc4jn1CTqs06OuxzKFAlGlNGjWiSwL2vH37Ci
MisgSjtJZExYW8GrUL3tDU6Pj51vGKhe7O9gtO9LsUFsdRHb7vb25Qdo6gAdMPuyEVYgTbkIOyBI
ZGby9e65qifZqk6ph+4BRNz0XZ6RliHyqdYWN93PCFXxtBtrsoYus1wngBUH1VSWw7IwwI5PUo++
ed1eQYBhSwKgFk4BG93wSXCJ7P/l3XaLR/6h21A8UJEXs37TqSF5u1DinHdfEzjBuYP5OeKhX+Ry
QTF3yWOTVSZ+cPr/O59ZmiCfB4TpXJe/1fNIWhN98w9QyEpWGJ3vdbDxmN3mPEzLvLvupzvWE/s6
h66P29/yhg4Qt4x4alVOvab16+PPY/RGdZprYl38/rRFYUUG5A/ANSjRWtK8zuDXt695gpdfAoru
kek89s+lgE9XyHCODquJNJUL04GKrWIO1Og8R/XmLu9/OPIFuve421GhVz3S9thD8/9d1bGhvG3M
njc2ZeTNiJy0urb2KWaQBCE/8UzbSBIR3U+I21k4lBrQ1R40S9Di7KIayU2guqkF79RNtehMQ7Hl
Ib+UDJU3jnZQ8Vid2tTrItJn2pXnkE40J4xCgC5DkYsXFqVPkUismm+YZt/1VnmvGb3jPYj7LIG0
9b3UrfCE28IbDpIGUd2ydR87OjcGqEMhwOgEk1IvQJwpJBEDG520kwuXZfwzbvlqCCrI9SFHh5DI
HB0OxQAc0xqmhvnDyNyV/05CQ+oQfhQMHEK+NcF28LRghTeggp+SZfKSMvNFGp4ok5AEt4DXEnJM
oz2m55T+KC0vkEalElzXwjOB83GNlmNbKZYxUV4+RNEZ9mefUpU1DWrsTsLFbQcVtYykDjSZUVr2
GJyCk95StRxA1uCVTCjwO4HobxY/PRB/QqQKrNdJQug3rN1QVm+XDSi7M0bPBNLlJACSyjHls/XO
OFi8GEbS4pqibvDAOKP2Z5ZG4qEjvZ9CYj5/c2iQD22a4lDGzEf0adF2dJN5UBR1ljFRduemwzmN
zy59UbYG4bUoEVnpN2Ffo6JgNAS6bWtExdChQGLaxTnly+U9eYnx2/DofCHsmOXxRh548IBwGEPa
u/erIvTC1IjSrNHTwLtIP1sq0xMDGzdak2sTiE+fOYv3tqgo/FyIeZicPajxiKbKX/M+iOEFofeO
tkG5MRNvPsl3v6Xnx65CpSqqL/oKU7nLA5j5vqdH5ZwXN2DyT7WeU4Du78QmZ9c/XIh/xA4rcwxG
2hXWuCTrJdZNI+B0UFAeEzVG9v2Xyn4jcah/YKFUangVGUxxewwRlNhFRIB41ockG4k7Qiz739Ox
6Fvh1FPEfiIj66r2ArVyBBAZMxZZSc10ct4S1lqtMMOU9zYJ9+QMQ4VDSjP3dBwW0mkoqxCs6Ggt
sBa8qSsoZqpOgNWeiFPnFNTAzwv9otTWePrEdWEjHO9ktaT8f0gjyRHvnImGPS7MfO4cPwDazIG8
4NTGkZPs+EhK+Mwi3xAbfnZ0k7A1Zo8JOQ6vmV7cVLUjTcwi1R/NJAi6vIKZpWgfPWvUPl6aqPoQ
aSMBguXgN49bzYtJ2pxBvl0eKNz3gyYGOVLYweS7u61idjIYOnYAtPfhAVjYk7QjU95z7nha7neO
g2jOQKvge7mKh4IGKwvqeF2NYJkaEIFDDQz5NsMlzOGblqWvtPDoW7Eh9uksJscbrZZM1uPM5By3
ceCVeM6U+N8bctRJjJdclIjnlGub5cXWaVGO/DfXKpMHuKXDiE4AB7+0Gw896OhBH4bKRsWngHVE
HiyaaXDDTLXPEHkuh/eJ3iHyQf2LYeBkDY1GEJbEajEQsGN5B+VEBgDvyE3KpNmPOjolfgsUuLDi
RGWBVai2YE9aZhFLcYxmLLiNfQRXnjt9cObkw9eKRa5asJH6m63CH9cdid28AZoxYSIyYZw1U+Es
TYHTlJDnaD/EiTMzEZQZiQe+n11lqkXNLNPRb6kHIHa+v8tkno3Uoj9Mva6y4V8D6JenECZ2HPVL
mNNhggt1tu9+xJanwZ2IECx8A4WsUjk2bRGnkZjiTpUeq2m1fm3kqqNp4RKd6TWpGaO//VluFG1X
6wVvkYCTITKov3XexHs5upMe9UV974URH/OBCPxdM1x7LtlaveiihfGOgZw4dK2yiC8g/muiQYuh
WC4IhwRS9a1kmCqPPEHJGvkNjEOmBP0ZqKxg5dp+1lXyoq50bwx/Ypl7PH+dRc0SDAMLpLxOaDR3
5F3gFdbsT92jKumrhm4b1AJ1ewR5bzeewo0wPxEPOnn8MmbugxiZONq5hm9Ts2oAYOsLK4EQiSbC
j5XHA/guCn6P6oG3aNtWpubTYC6WI/osIJGD3Xy+V+by+q2nkpwXqX+y4WUpWcMnEQKsAXK3MVPL
LcFHA6q5BeuoSg5XjGejEPas67oUDvMTm6/e1U3Nc8qbvkYRgAKo1jyJ3HUQjCTL0uK+y87/QGiw
wL7zl9qdPQaB3k+fKe2Z7uAgZxpswnXBbSt4RajQivqUHyFzsncDun/YMzdzA+NHx2R99uTY339X
Za9PzXuE7oCTCPi9CwZezjRhaPhuRvjw4KSRQ8QUbXxLipPKO8WfuK6egFqMq0sO3zxeYMeB/6Uw
8prKTEz8warBEeCZPo8FlQbj3YuLocqza/A4g7V/Slf2UsYuslESYtOd/2mC29AEpPL1xSZiK2lG
y06pI+nwafl3Wc2W//X1YKvq/tZltWvp13ilU37eM3lyuxCjVBfGXIBrpru1orWckIUS1QSQ00D6
JpDqoSbHTozHo1jIEMcICJXssho589i0E0hiHBXhNBnJeB7hOqrounnM0riMRW3jiWCBNsfVroay
zIwjfMEoZNTT6o0fVJKtgarLXq4dkj8CBwSl/F70Uymb2mb21B+xvK0aV062L+meWFbANbCiFptW
oPHphxyM57mK6Es42pvuWNjgRztJNrYcSO78bS1zkrmUlaKx+eUwhBwCSaF8HDAGu9bVpcmXBMvK
DgblZjOqmbCkY6bZiVxyWZeOhmdzN9XnyUwMtw4lRBStKl80dI7XNX+cKL1Q/qt7DEwz84AthLgr
YoodyOweKDMN/fIz55YJRK6rRkAmYlenWbK2P0Vq/khvTi4iNVMizocuD7uC7bpH801AlDl3QChq
uDm4NFBvtFK/+U4aW8/EJlEbyVlE2gp1Ems5R9na50iOWcFnQBLrJregPeItEnlRuoTAyrgbphJm
0Ltk8nQaagmwv3QQmBWVLoG7dc26AVnuyfYanx/qdPee0hCoPeNusFugDi4LqcJvPX15Wq6mCUKW
X57O0dHUn7o+tfSFD1w5EJK8WSULubKfXEKiqAI9YHpWzFZEY46yg5clejS8AUafCu1GGWTao8PL
Jnx4dGCQynS/tVUzu2LFBsPKVJGNsBDCe2zfRb5huqVPl0vjfoFwTaufIXXYydWCQXWJKxfRZ/BG
lExHNP686rqYEqqZRVeX9iQv14FZ7EL65qjiWB2DssRc2ZGXhi3/PWLJG2OXnAD2OVo8fMyOZ4mF
3SDthEdw2feu9Gc8EPRq9bdXoOpS7WnCKFM6cTpDyqA0+bZPpiPVFV40vDbHPvcI9i2oarfhGoKX
gU53X5lK3ZIn+u0/bXieOyBKcd3lN1C3kVFiyZ4Y4yC/vj2hqYesuOAqzB5jla37cmNWNMnOpO/v
RxtbbHu9GMYdo06O2ZsX0kk+dc6qCsyO4d5V8518ma2q46x0iDHNE51ZFRfXK5bHQuvyA0KzMHvi
Li+s4wafadAyVXDr7JN9O79cm0d425IaMbXOvieGV/KNRP7ShLmRoqWTu8XNm6DyB7WbTvMrmTxF
tKZsl2I+g3NdRFd3mdKThbsLv0/XYsay1inrLzeWMd+D5S28FZW4Zq8Rf4LU3eeIhrNXv6tFezti
CuM43UM2Xbk1RNTlM5rqkJ2IAyMR+bRMovsBAGQmKxBIeLyd9RrjHvhPPZgEugtpjCQiU1mhe9qd
NuCTH+wn4EAJ8/noRb6PeBr5hY/RzUGz9pdgcxEQuX4GA5eGM5IHlDQDOVojR9GaEwDTeZo7QOyZ
a3xGvn/+jovfymHd/ze59DIa6azpMsoZpksuz7PCkArf21E3J7/5ZSX5NbqQGVq5d9JoqqXexIN6
2afJjqJdyjOp6Xe9BzVXh+C3okdPQQnvQ5maO1FgyM3UbELoPTCRI86SnnF57gE+xuvdF5/L6ujj
6lQv+tIIfkPTBNcSXlr9rPWaXyrnfEqdEPpfKuOEzQpTqYl1IqqOR1A7NZw4CIjN/xrnBZGfIt8Y
ZAtSxzvPTDOeMLTqMSDfi2+jdwM7RfYnI2UuUv5Q3L5RVVdZf+V2G2oFdcTr1mzZFL9nBPgbmwhS
ZggdirJ77djw3seACxbKyl5otJHRBIfaBVR4EX4VMdLz0wgyp2bjCiVYu2/Lkb0iNPL3ITycd+Tf
0gx6wjDh4Z4RF3Bq8+3HOjzR4N+cHh9p+SLIlqObK+5ze2sCJ0KZE+wrT6Rn2LoUXlHKwJryTkic
aHHaAR923q3+8tIOKzFN9+2B9aPE1+rFSeGX9Z1eL8tuz/Serbbh1PVlBvE6Ut8aBW4yIpaaK9nd
/lBdlQOpx75z6TIi9x8WdlrqM8/wrUwYPbDdWZtYlT47SeICx1mSRXrqmLu4T+rc0uHu6B7nxUY8
lxQxV/p8VY8O5vj4COVZKYPw77JVCEWMqW4+SzGIUhQursZ3z3jMkXUOTi1OouYakAtelmJ3bHyy
B5GRR2s3WblA5lZSkZ2OWfBZsWAyCUgVL5FZGQX7U/F/0KNFVfrXE4Tl/v5V3bD/TeZS66swrYyz
sOY6ZG7ry1ENW6uRu8Q+SwTEJjtVFnqGj2/KcSZJVPw1Il7XrpfWYblHQuuMlp8IhMpnO+8ZTC9c
JylgwVXMbAsHtrH5Wf7TAEgC+aLAcjCP5XiX3Yam3ZW8ZohVp3m53zX/dKqPeAA5BKvAJ3OfuLnp
E8Cn5vWJ8q+XDI/VxuUH6HNDtqIgSs5fT0Rvj1XL61agptowDp0Dy8/tfWW0bpib5+Jd3YhUrsbb
iMUvQNAH4n8u8ReowfGgYzl9Xkc4MHmKC8py1N3lYyoJom+ykDPnhE/PudeYOJn8bVRRczf8/b1t
eVI5KA4zgtF0ZMREUTxIBCBF/pyQEKvw6luXZMMM3tjCSNNU4aaYwmWQkMrDZJ99nnyRg5jOwhX7
X3t9STWb+f7GDY3d7OUMpKFq2I38ogY6s/BMIsNEu82GsqA7KzmE4vw+GB3N8Kkw/BvVXWOesxiX
89Wyr8+07C9XYLDZ9Xbnnjjr9hvYuwvCimqFN6h2je42V6d5MsWawS+1z+iw15+8bZIO0He6aUkB
vv0QLbKB09y0MRrSHCd97QqKRaBhikuQnz7n2e3GCaNnJMxhx9EWsovk8gwX7NR38nuTtMxWUVIg
KKvdO6+Hmhf4I2EfOdjUd+sI8IW5q/wK7Ao2+mRUWg+3n2mfe0xmQWsrLqAF/+hT3GdwBlp1l0Fu
1k1NBrx4qJhHpI6a2444s7F91oRDJH0lYsoOVvVeUGyUrUK7QYuxWZuYftB0rEPpykTdBkBtubLJ
tBL26H6uE2URkDzJWNHJdKPeU87vBBRJk3oCmq7OkcRhxYrgz76BZU++93kHihupvYYmJ/pnZapJ
v6DpZQG7HRI+IxgXYt5uY5xwUCUyL7H8div/sAvFEBB3e3QCZvmJsn2NdIawqPdIalFb7TRWvc4e
896DMjenAm7eifHSqk/lteerFVacIeDUhMPTm8j2BonOLDXWRNhlovTRrNGXzBx3XYCPCsk1ax5a
iiWZ73lyr9aCzTGO/YULm7xPe+zx51dPoTHx/uy2kOODMxNsZYcs7hlejDWDkEpppvYjTIb6j8Zu
MVjivbjD4v3vOPaBOpfwiqNnrbe3AlvtdiBW8hAaHbZJmj3nM2/AiGJzGQu9Lg7TpbL6Vof+zr8l
Vc9EuKKXwkOB1NPOjcI1gxXCkju30BHzdXa30IrILG+FPueKGJ7Hlspay7AnVaEysT220Xq20xXY
UwLRl0sIK1PzF2XM3ESuBhBHoni6Y+DFnx9hwZ/Qvtvd/6PmiptSelhDBDngXLgBgGAipDkVMHqX
w5goo8EbSplLAK//27ycv1LbPtZy1xNQLh/K5bhxS5AZKvI1YlLNhHt4zmD48Gvh/m4ZE3wiEIMR
4gdjitfb0f8DTLWJz7KN0FPPzx3e3o8odbjcBoAJNOLZs7/rKmb6cfrzVYrwKegPnK96FW5YFCYn
iDP93oDNHad3jwKnfBUWBcddY6jw0T+thDPjfpDW7mUYHBBF+oxmIGexdGresB6VjQO/GWNOmGXG
fE9W1Vuo+M+3JPqCJLrf8x11g1vJTc6b4A7WZdIK6CvIe2W7VdpVSxsGtcditX+e01a2SWcmpBwV
8d8bJnO+4LHzL8qbLIXU5UqI7lKa71BYZVzDKsijUdxjenNjUMyebXlk8y1prHFcFGdtWOJ2zO4W
8KMI0WjR65E8mPCybmfE25e/tUhkugvywwAA8DRRsakbXldkXW9HLNxSgGxD6i0t+YwM52eeRmCe
djjKTVVmI8LIBgqyWbDL1xxgwk75krePswKCgc5ueSRuOUnhTf3ejqOoYSF7royV4bnC7wnsJGua
lLl/+luo9jXSOqdzNTGE4h+RwUohhuttaZ2hpZrsD+TYnUpZTTXhN+7JmdgG/0Db7jtLO9ZgvnCf
lzouw+9KnVX++sJrY+0vTS8/oku0XT3IgxECHwH7yIgqyv9am4yL+NPEzASfyKSw+pwNnF6Fl1D6
tSoQaAYrhU8n3tMJPc5wiCVLVGaHESeYxtlkghUCLYn63GR7GOtBWvTl7DCeY5bT8Gy7DtqUgk/R
irN7rIfLqn0PoaSEzWZ2oGm/wm271WKF0w8DcdkVfZctByiGr8PQtWaF87Xsv/mGQheJKfVvGWZt
tkxTUHKY6DMNE6vfjmlLyw85xLQlYOt7q49wKtCgZOvRiLie8TfWlx01H9cmaEkP2bj3NdjNVWpy
r0lRpWFiUcf42TyOZUPg9iFCN8UK06RR7Zl1T/cyRxCS11Yxm8fdFCx1rAjlkgVg5ugAhwhJYJW2
tyDlPF9LJOBbfSimDTazYEIzE2+pfaLGFJn2qj+BcsnabhO1qLprBxM5S2JOJg7+YUS4BLxELQ/Z
GIo9Exa3Fzvd/EVH3JcS8YXFupzLhPJZfWUi4dUJ5jRNWgW9acTXp8+vRYzcv6qchM994H/Wn6XF
+zLNoa5xToHgeO+4LXn7TG2Qcj1MLYJCNhHoBho5/C+Cy5+O6YVBuGkdTfd7pCt8rTMJfvCnsvoT
RC0EAFhRm+Kd6WSr7SzyC8emf0LUbyU5PesltDLhoNyavCDYtou5ZYNmq9pKY0wsniWP9FQ5Zs6z
UCBok9pRMsa4rT1Ulb+SqrRCYCFK8fTmjWittAexUzLSiO2xEnyecjc0kA5eZ+JGhGOc8BkVDWBb
1+/592nLGOByE5sqUIrddU47dWoOi4S8Wz9yPiq0/zePzR7swNePwr8uIlSF0DrpfeJBf6FOVY9+
fD5xj6tvqdlNN7eloc1HQvnATB1CkIVRJ6bb7n/nx/UtfjfmVUBNN+n8Y8PN4VYDJpHla9Gw/OI1
rChCGdTYt9a4LjEHhX2bWK1idQXPrZWOAwdjUgYY4cUffDHH9l0wJehFULD9Bvc6g0QktL6xcd9Z
QLwJXzwSC5Mfr5sIo4D+KUtnYeV6U0F+9C3HMG+EzJHCQ4lMZegdSz2Sxo3UswdBmIkiCMz29hCi
5PXHpkoL+Rwgj9+zkl0TeogDf9yi6QKJBC/qUU5QMHTGk5tg3s5wkqXNI22ImL2G75i5AQMk9ZRN
g4eYU8oLOmMvaMutyZy2/NqjFMqfbCsjR6DUXWW9Ajy1QXe0RZR0TYU+W3JR6zt+P+79rPoG0XJs
dJZqiyX8pxMhEf1Vpb2zMZIl1LL9DBqfUpD3sSBPAuz727bpEDoZ/+n0+Phy5mxzGN1FpYYCuh0Y
2YW6PIA5LNSkPKOXUsbAMRdfwfoojcBxXUKshhvQrQRlAU+IYvEmDB0nJQ4TL/g6ZfqK7aqbSAdl
DihRouSTm2Q7LJcCReZjt7QpCWipgf62J4x9i6s4039YrvNESVpgjXX5BRzgx/hsCll6yTpL0Pyd
4LZbVb1vImUo317jDeaJBM45+Vw7sXZba75nCH6Ed5a065jxHnnEpEX+Pwht+459cXT8j422LGpQ
DgrQBFu3DJ+WZlzI2jhcP/BNPTh+nn6tN9L1GuluqNnL+1jLIZYo1KbIhY3mxoI3HCzC7D+6+T+t
C04Y53W8n+VrAEvnx4g+h8BxfkySOWI8l/3/LneL/Wb5uA6H65LRWq3vRXIQStu2HItS8jTA8NPf
4QPRESh/YfC/+ummGJlX/IVVIkzhDJXXMZE2PvkruMmJnLT/zJkExrrtiT3bncVLqGIKGJe/Ylll
M2T8046PEm9At+7cVtBiv3ii17nV1RcIEVn/vcv0WZMSLT3/KoX5nO/IKArB3Tgbaq8nnc19cvNR
QNFYDSSYhQdG5jimKMUlvhPjLM07ErmfvL/Bp7YxyUARS1FEf0yXJE77WlNpQhRPezgNWfybjWSl
BtV200i1eDs7p0RWeD1io0zxHeIXkkX4Cpumhg17PN8YP+7ooz+OYcrlE2hU8Vb57hi6ywpinWI6
yOqXEFbG7QDA5AkDIBRV4Ff5vBFlNx9eEpot0zYL82iUIBMgQ9PsqIBtEq8XpIu00ZZ0B9NbBscA
oq4Flzc5km3QcQYCiUgQGNK9gEBu/XGaXDXQgbVicoTYVvAGKwey6XoFDJop76skqhfQn8sUJxlN
E4a0en/WD+F5lzsUESpCpkw2fAlw0Q0yfEyefI2vWA0ciohz6kPDbPIoh2WhPPqbymEYQo8WsiTW
FSRGh/zYhTJ79z8TAMpXw2OIFxCgqoTE/vqJPNGp4aMpXPICistnmpK/a3UIAxB7KHYYNnelH6dS
plcXKN8yKkgO3AVhm9XhBwJ/3jLETZLNXKSUkAp6sxQ4996gOVfN9QXtSyAKJheKAU402EpxeEYu
2S6GSi8tVL9OGaq8cQmV6jTTkM7YBoj50mO5NDdj+e5icJx+WiTlTGxiq/tT3AW6Qf4A9FIdGPiP
3thWc43ykNgGhfMLLYVEex7R3y9h2zpnwZlyfT0q5jYNyZli8kMxzx/SObUXNowu8YNtjyUI8GF9
Y26zTC7gI4zsinkCf6T1rMrZv3dmu705KyVuiEtaBJDBKdnJ8iz6ed6SNynb3sJoLLZhuj1VsNTu
+15M6Mzv5C7uDX4c78YoWhO71DaQShKpnsMb5XsEoCS7MbSsaxqZ4pxoK2WdY4lL735RJ3oYN7Z8
71LlWrLp2oBRep2hlxfgr8XdJ0nFOwiN1M0JE9zF94Nlj4wcy6Vdlzje+5CQDFdvtn1hpdwHF8O3
wyI0DBz34P13EPc2Td61iWVO4BWkuO7Nc9Yeovac/maVoJc1unQgFKrc5XVUKqfcDvZoxhHrD2TA
LLONH+k5wwcpHxjtyAs5dr3wYPnXcQvcpQUYR+2QBXCz+LqylS0YP4yqxj62L3ilML7lQNZQ0TwH
RNr+WfoM3N9nJc7eibb2NhFgahMxiVJsd3hkwrkI9RBjPBl6z1V9kUdVgtoLqpr3SM9X3b0M38k1
HjLFkJb3WcU2PZjOTtIXPv6uHKq4yYT8/zYY3rtbzy9f9JobLaZm1P1HsKPgpjFCJSw7ay3o6j3B
i1bjku2MprbWL4n4nIZXhrz6M1AlwPzAcU0Rg8CMmGkJ9+/Un3XK4tibJXAuVnW89S0yfX1wHnnx
aLM9huRvj329+15qWUft4dhhv07lEK54h653XDHGnXfmVUMpHx0FQ+LEeHwPt0Ja+rXkCUwpVU6B
pk79+Ik85Y3BUanzA8eFoxRApL16Q6zJqcHXjPI5iIqQqwYXvYD5uwG7rndyULCjFAYb9FDVmCxv
b9fLM04+SU4H5ZG/Pn/ZeR5dQoyD4zFGeXViCuCU3wvmZ9QHBHqF3MtIMtD9VuHssQ2od7DjGMw6
ocyB7L4ZlkyHM/jxjpnh2J5m0rD6ldB8UHLenXjIBoGsejZAEi1LK7aF4XvFf6nA0XXv/BUxcTcb
dE3wmeAYKHeCJQEJmX/ZhJYv/r5a5DxCsXL0VRg2q+N9lw3AMbVUviG3zTaqZ+vOkzdQYLwb2h9r
nQnyAbKsMg2fGPYGR9ErQeKpbiitTiEVVRGyRApSOp6ru2q+pbnIGSbOzcFSOGfkBBgPbsP8QLVU
tjylu/skf2f/cQ9rh+3pji7VLPdyIdFGOA9m1A1J4XhmHWAp0mO97XLr+KA9P5X3doDKpuw0GLwQ
WiJhfUdr8qDHVjWRchN5NwU8W+S6CoX36vTOlZJi5ee82DqnA9bgZxmVscSzBYB4nNAxuJbEnSEq
UBlOKMyYg6PlY0JqHtwjS/RXHVwEywSFHETxwrSyvYVibjWd8PjZGsW/fvJIQOWkBF5l7srYypAU
pm0+NwAwfPTKNgfBx4gVfd+tKodTBRv5W/Qr5oahpiO6mkNcH20Z/++PXL1sQ9aQ8wHoTuFurLmY
AtYTQX/Id8oZIXx6Q2CdfQgkr3+LR7Vig9K+dGdCt+60Uh5eelgyT2CW/unTCTDu3WM9KTiUoAh/
kni4dl3qy3YcoWurNzBADXwNKz/4dsXedx5ufqnO8KKn2hEXbSx7jjpWrrdkzi9SgLzDiDJA30D4
6TkuX2dbcwEWnA08cHVn3wAf+goEwlhDeJnvC5LneywH7MZaNkLjU2EwD0dRk34xOAfkN4FWxNZ8
NbTVpBtEydPOQFZgof/0lcC0eGOuWIMp/khktc3KOy9Ny69jCpuo/7ys7k614tfYiXtn2CniB6Qh
wZ04fMBdgPIHfZIsjr2uw5x+OblLwNwzX8Hoan40MYrpuRpOlpHkyB8LSqmz6lx+zXaXTXsye3iq
e35G4HJCuzvw/JwSeC1hFOMRQ+NZJCaJiD9XNMLLBqQma7BJIp0phi6Pj2ArwK/bTlBxC92Rjn6U
sirhVeuN8qCKlW5at8TXrgOofrZf5Xczyw5DUH6YeZF1bUEIckYg8iHQvd06EG5QiaGDQWZb0jsw
NF++q/433itKwO7AQ5r5csp2eW2Ru3hmOqtOmvNZJ7ENsH7Uwf00wnr0zThm844OGtLZI9ck+cAl
9swk0YEMatbOLQWocncHG5s2b6yxRj6JvnR0pF/d0j0AwDlJd9L67G4NX7zi2+wMLl3cvweb4Nqk
n7nfe7YztP3Vt6w/hRsax++KL50w2AO/E+Fi6EwzEja9uB709cYtb5kvWj2zpFQu0Bu+BFhsIupw
MPnyjMk3k9kxlrBOjG/Jg9y5ejvlUGDzE2yQG91umixZVNJ1MCpZVjxIy8s3aCU11n0Mo7arGvf1
6KdfDKs525AZzklvVzUp9MQ3JRwxRRbVxJzVmwVnFh4IA+8EJP+P7vZI03DOSWZGqqFxwMNUILb/
EMEI4ookaviP56utqK72IbrupSZ0tWQLiwDqp3ncg1fdNA0WzOi329H3mQPi3YoXdR3lbhIWq0wt
vwCjVR3qvC05fzsEnDr2uKWLiWDAvDBczm/k/ori5PQkveo8JxBXO8IHtILY9pJ/GEvBbifKRTYi
3LLtoEvnItkLR4iNpFNV+Q4gO9mRM4DmTeLwl7F93vg9aQpnZ7SpIziQCAJc57WCOCEoPk6jKeaS
ikG8PRW7z22BdXBRUF+CG2Aij8rFhb6vMXuezuyUwb3oMWfFIYxkWrNkZPRqXUwQqkdN2ITwO+ow
DQ4vA3nHRio+sFXVePQWYB1LwrxP6DoPLSlIn0ziypzCJtQAUrpi9UWxebwzL6iCfhLZ6rJ5tFKI
SCdKkve55zNCT8DTAlnWIJuQJW8ctqkkMIU/AGGflNCcM/3v9oJoZTydTYTIijRJyaho+SDTmj7b
s9MQz7A5441XsXym0mIxy3/EV6h18COc1z76SD62U45nqxlY1DGG0mMMMpXeWT4Q1iOrdmzW94q/
F4JrUtvX0ZxYw+2tQDlXKXF86o+Buo2dBFyAhHe8hJuu/RwXS7wK8vbTy4tTnuk6CUAW9jgBUb/K
Q5Suo2K2chtJI3ONnJg5WgilhZUAhu/nZfgJpzU8nyLbFYFuYEzAUeQRDhan5Savmo5auU/uDnux
PlCpoI3721v8+4OX09JDOt2A1BO3gkuKlFA9noa2RCM3cgwP1x4pPtpg1QZzDaAdjI+6lAYgl/c1
NTwUKZkqMCL6WpzHFpGWwbNRVgZZbAJ/3TgVI1y9QPAv2tVPZFvORay6ZTyH0rgmkRfTyPmRZkjm
OW1EuY7RO5F2l1GNidIu1cHIE5tHwmMeB1uDWaeyimheF8EcQva7LANFrAt5wPZ6/Yceov6vvofN
r0cTK+aoqwy6dEM92/UJX/MSggfIP+vcMEQOYUSHftg/uLrvIcvXKdMPu/l233udU3Tr3RBHD712
DjpVYqidQuEQuqJ2fCoOw7yrTG8ogM6k7+m0WSYD9o8jVhz5oojsKK3hkeOrvn8Lwom67dMDJunM
ZSWhbMzONjjFroIUZq2ZElvD9GbK1A7SkHw1qdSvd3hguU+BLgxz4I5dQ6AAoFGW56TzX5buuGBt
eD1NbmMvZcQvmFVdW8F5T68197PTBcJNkELKcPg/zFFtGjWuS5vDaNVHidZNQ5REetMGt1g3+Pmm
K/5RaAi5FJKniQ9ZJAPDFuGl0PD/UfVXg8dIo1FMv4pWV4PwFa7ACnPVBRiy+awOptedGWhW+kw1
wSPj1LlJdKMkNJkSHEgCHdE3LYWHfBGIxMa4zPxnodSp/2nqY9ZjIkVy9IW9m4z0L/Es4XOv4Idb
khe9WprJjCH70kbtF0pMSD452Swp6DJNL1/Tyy1yUaXk1CKXGhXfsTZkNk7mCss2k5sOvKOUsOnn
huU0ryGqQWe7INXRlN8x8Xj0eunoX/RvucTzgYMPfdSlje6o8e1TqcTPJipZEFMNm32VIkiLIirP
8v624pEe5pcSUgVIrVCXh1rSyAy7gEdLr/fXOrYxdJ0V3Vm1cQAKILmX2FzLLuYX7ySG21edSYqc
T7mRMpU0wdF5Ews437g2GSarpTlF0d/arASsH2rA7ySkrVjUl/d3//acGJ6MGsIZXnF1ntip9iHl
3torznE+nwrjduEfp7WcqWqBL1Y1Ng32ZY7tw7eRWn+gCioNzqmmicqJZ12hGTzxB7uy2B8JnKcN
F9CZJeB4t0Qk9kSvC4olTjHB0KR9vNhXC3OHzSvR3CuKrX+bSd4i0IhSG20QRhbnx4VjUn02wJ87
88U0m+F/69MeIrJXIHsoU1nZqAiD4flB7y7caZf5AR+qISQDqcfbe6DpsE9HlszeTNQbA61mkxw8
SQHvavsknyGb6vO9VCulMw6EInSEpG2k2rWTew6GYSaFaV8EgKOqHBgcoGTxx3HUKw//Hyq6bsOP
kMbup8RdwbzEW/wL1QcyGMaCBHhdMzh8xK2YBskgw34xUtt1RA425yjdi9/guJI3IWgnqSfrlU1D
2rriMvUFY0O/ekePua2VbP3IJD0j0XyHyT1tZZxEiirvHISwaAJAgnnfCIYiEaEmpaKzIl+NmtsE
NSV/2KAIXRG2XsPFS/DrFmsYbBIxoSYQh/OBzLeYFbjcXyhr1b7ReleAE8kj2xYued1l5L8Wr2FV
eQ9Fx+ga+zL4KsmglAYz2f5i27suNYVazTHDPwiSR8WJ9CEYbbnlhZ9SQn4Jt5MWqwtbYILNFZxl
cBsKQocgVixBkhseLdv4iWOb4aNA7KchEdOKpkzuPQW1b8luBR7Tai6qbrkMkhipfFJxNXidpGwr
i4AfcBV/KHoaIfclP8JF9xFJ7xEqWRtEhyFx0RxWl2FUqN3FtnGkBqmQu+cQL2XvRUlRQXotcWVA
Dm242pr4ZBSGIX70oyDd3NB0hIfL8VWaJoHnZz0pfItO/kKlcXH1og3LiqEiRsOu3kYLmFKOn2N2
clOmSctz4Mzf4eTWAcvS+wiwHADvFt9oKoNUxXPLVB10R425b9mGxWeJ8Bqwz1k4E53xEB7wQsAd
rhhi5e+kkn5Mg6FBzOC/Oj2g9BN9zLOJBrAPvd6pcJeBKQSRzd86fzR/v/Vke/PoHj1QPFrtORhc
ojSZArM1lYPmRE30bO+lTsNf/hOkVNxuoEWCQTfLeQ0pLibNQoAMME1ahO85zLQeMcOH+UAZAp9M
uhrd+bkThXHZJsKkhHwPykDR26yb+LNIq9eKrDFQOP3mKcIZ56jbsVfSeAq5/S4bkSCfjNSAWCna
wZBEsf2vFf4dPWChGRhRbTggUh7KDd9frGBYdwNDeXAA06OEEnanimPrk+qrzFUdElt0qmmVE7xV
A7KXz8NQNy8jl1RvBwvsu1W3ZayICQZsEeDB7Su+peLlJmUeTonuQgox3ruoHzNjX0JUpV4A0EnO
SwClEX7hvytFsJS5LUY3JDtpUONG9f4OOBEmuchguHAXnM37coFRbo6tB/N+KBWlPFOARApnqc8y
H/Nt0AcFG8E0yzPr+ETU8bQ5/jUM/slqlFx18ZQke5DNYg/QOdUYkP5vojGZ73Dr7U/+wAUqknPl
RM2ktRq8eeOCK+N74oa9QVdVL0kboHSOjp+OYO5qQi9S1v0GJXxsos3BSL9xr5gf80/1vrcntdl1
GxD2CvfbNFD5A50Lj6GjNdFvW8gmOPRtkPUSooLJE+zNqpcICw0TsSGTsxDf8TpZa/5T+hJX5XtY
2m6Hj5swl2JKnvdQwCgNi2SQ1MR4NljVMPKWNP1fYxK7uYeyehLnokM7g0zjO+lozPIeWAc95Bie
pCWdmaImDxtA28BBBY/NC2BzSs4a9nU/OOQaSJWbLvSO8FapvOtgEHcza0iUeYNPVuAv55kjkGI7
HR+JBF/a6IGwee5FXusHjy7NuV3gKvaDdlqBNrQiD5vuc+/UJrUzs1UWwob/stqs3oXLmVfMCLYW
pxcXTeTzp0JBeakn7z83L3bBmLAztlqnaHmFXTcunJGhKk5k1IupvnjwaZJ7UaLLA5S5xxHsoz0f
HHDQmEpElNTVqmdCLyGBhqro4G/mcWbEB18Tsw7CUVDohXd7MaSUO1IFpLVD62vnCjGGZEZdbbKa
/sZZJNZjLCEuChy0Y+rDbCrfXROuPLD5OyfIACkvda0PztU1+HAcRAAz8IPGoOJf1Nf1rC4igm8U
EJ4AW2v7o2pSs4HKbzU0A+eeNoI9rLpBSVrPrxxDVZPrh/Rfzz7UeRGVFY5EOrSTqfxzc1in9MQE
aG5N4jwxFiUbMCcdb6rw+PTBZty5tgi3KJ7eHGu+7mMB0zjzvke4S7PYUylGyf5ZCir9Sdm0rvfW
E38LQIhX0io3uP2kyecac1EoxQUsMP8QGPQUMc9WV9Btj2Q7ug6hJ6Dtcb4gUez4n11VUaXXP/de
ilrXlBAt0wN6TQNBvz55w/fb7UQ5BGAnG9twBPisUqmDbq6WONqGLL2Lfsa6PMA/jUhx/cHsZ5LY
zz36pfE98ond2Y0GKMefeAWRMTF6P75ewQfdplEZeZuYyQyviLLLr11zTXAsBysbq6QYZICh5ptR
6R14WhdQNjMiC7IFWckEBX6nSAtMBgRvZj3wemtE+kWXbrlx4GsG9gMxpIyYaK6Ro6PtFt8w/xWc
rATi9fyurCjWDE0NxcTbhnrMjSISa/JPX0DvKMyf47Y3NwFhaPwqv9srjyT+yMgU+8XeSFGsWYmV
KqiiYjTC5LF2nNokzE2VdafFdebYFrx/nvnzROI94Q+OFV0eUiFSgmqU/KoEiZ86pBxEx5frJGgT
fv2b3BC0arIrXpjW9zmo5P+PP/ZdJuNeM+n94jkRAmNWMVM6/IyqddjqHDsSS/z1SxdbdEUH+jx8
mJvQetgBGZae33KuElx4LdmIUwYx5Jv1xE5tm3+6DLn6ZZgRei9u2NUjY6wje9CnDNVSutupRpET
uWP6L6iWK6NV1hQKn6YMtss06YOM6mPsp0mTSd3c1yAZKmVXaoI45oiisH1PfYDgKxmDLMFGvU1f
wCrbLoYa0OcQGuC/bcD7LWQLwVffjlsiogVWmUxQQiVj4MTpTwYV4TEXoI1eIMVafx1W8mvQzP7i
3T8UzHHfgErTQ7b7osBy2bETAS6WQQcVYV/YFD5UvnELn2FqCX49Gl0VA7NtnlBbQFptSAHw77m3
6Sx7VCe+5lIb6mlpTc/QHMWOn8SZcYG7EqpWlbWnYKWhvONLNPi2nICu8cNZEYxAI5eWK6kw0jAI
HXkTrpvQdrfz2Hcle52QZsEc5NsoOlYpvlb1EvO4+i0qKgkmYfJgGYYVmHZ07BBb/S0C8y0roZ5f
m562QKqjaBH7bisoKnY6fJxWa/QD6LWAPdCZRZDPD6S3kU1qRve2e2LdUixxH/yMmEr22KpV60FD
3C6wUrOBTNerxr2ISqh3T6pgM9KMoPe+0jrhgd7MfkijrmD1ZjQAUv1aXuCgyPDGADss/zXJl6x5
yU0U24hHnjtZ074glLnD6E4jpa8sgZYLvgvl214OsWAsEyTeJmKyHFTwI5dwlbiDxl1rN1yWdvl2
awCA8XvLjS2IH7UQ6r1LUs0YbcxLATKFUQG3MY5HwurOq/fVVcpfGs6uS7BaLPZWLbYIiISFDfJB
1Ekk5v5Gu0AGzBw1wfj+hWK1Pljgw+yLn/COzguLhnzoOrUOJzuOZQn8X7cYrZM01NLkMElb8Tpp
ZyZDv+ymoAf+UggjCH7MBj/DUEmBGhFEIM3MXurnmqAm6LGlCKhjILdypKa79/b+XbrFK349g26d
M8YRF+rjrYO+FW58sMzG5bcL2FsGTm65Z9KPkrqG8AHBCikrZXMuFC9x6pzvC+zAkrtPhC5v69ON
uv11oQnuDMmCiDrJsmAD3hdj2DoKlOQoDYip12+ubQyP4Q5ZuZoAmmJXesEtR9Gb5K7yJ22Cr2Q9
TfISlZVIacAdfeow+CgFTPqzZXZXn3dwDXQA5LC5U/VHitqD2lisfXLROf3uoGxp0FIfvbya870D
UGKn62Eb+LME8BDMZruXCJJ8iTkn2tC9RTraJeAOUu1AdOlzM/BDjrtufELoMzPfTo7JIoKK1gCZ
TLJiLcujr9vAXwsE7WR48yKfJ21naUZKl7cj224sRftofjnAy50jiIxPrLsC38kggQeg+F3e+aGp
noDWxtk0ttQcSuTVH3dSHjpfFGM98nxthbrIoR07KDE+RX3U9oKPSN5E7anHb0j5VMLpHfve9HE9
quJvLZ+4aieFXEuiuv+kCtk5yfxK2eMtitrNxY7UWRM0zh6l7qlbm/FlQguXrkZFo93c6wanNHjy
ZGNKvCInE42DPqs/z9njLsE+E95SY8hPNxJ2hwyZqfQivcgoCiaS79opUdryuSQYCGtig7nz8xdB
nO65VCiZSSFfu/cpII5FypZqCiM9JU+96ZbXQbznwkQjUJudtgQTz4ZBiC6nPr2C04vAlOzH5+1a
QvjD6pi6U6XBSJiSAQzhMR6seTghuxV0236Xtt/TpQ1IccxSG2r5uKAkEAFesWN5D0t62eoO8l4P
aqCbFjmBDt17q6bVqGx+NuThJ0duPVapegezSHw1ZvEkkVju2hD7h9lEDJ6MxQoudi4V1mBMq57f
LcsfZ9kQnLnuaIMXcTyghRDat0HYVdbcOjl6YVw/tTXv4YY+LGR/O2hyvpbXRFMbQEjXxzPgoixt
SDY+CUF/9E/UtZ/17oxzZ1pLIaAkGUdlyLToQ5qDoJ7hiMeYsryzFIgAYkuIcaBEFlvXWnGD7XPp
uZOrxO2eQxnC80sByPqUuz1a5+G8R9LAVL5frpfk6n2c94zLwvxNjzxwIaW8qhh/K5qQN1mz03EM
o6RNpuzA87cbVnY83jE7iK5CLhYnzArgL7+EGA3Oeah2NfsFhKLKibsNT2mp5QSvjJtlswex/dKL
4B58+B+nsC5x66N8TE8lD/kpKH4drGWlR2ETETDk/D4wbP4ETXBAgib4KRbnW8HAQ5uYzxouWYsT
nM5fNJjzO25/eGdMPk0UD93dv5k9wp5UjdUKzYKXg+YgG+HzX/cKjD/o/WjdjS8dn1Ch26ftZm1f
ve2epM9Vd2tnRp4AZ7OpjgtUUeBtGBRqksj2UK9kCgQBXcwODJuzXs32w7tojgEAOSffEU9G6S2D
bLDgTVVPiMx/puxbbm1jSq19LRM7NRdEvInsrPoqLFerad7Kdny3iSW0IHkKsuLEON1pZ29HD+ja
YNFTSw8ylvSuEucbN84lsbZ2Q5WAkaYAdKmUe7uo3tv+WmsTPtg9b/5JneB4vTSwaTt3jh5Y6OaQ
sPWorWifZI6CZ+kMq9ObLsyoApTiM+ZFZCEet3I6bU3fxSLJdDZtsHN6pvWVLUy5n3TSdMMErC76
hPRqay1P01jVCmGPVncH9RxVmssrWCoWhl73zGhvOfNSh55FANvwj7TvM8yHVAqv/faQVOjwEllp
0zv5puGWdDlYR1LEEjpE91S8OsdsxE7S/vUXgRGfmofEYQ10VOv4d+qnB9cVCEn+jDGFuO6us4vD
auua846ymn7OvpXMGBMAx8IKeGi725eTRBMzKvsuw0EWoll5bcW2toay0AEAHX5TCaQMFb5Bf7Ri
HUxX4A4AGmjq1O2qJoAWNnGE0XkFxrF+9bg2B/f9iMDrUlX70gF5ztzu45NHXAc1M1C4BIsbwB08
sJhRRmdA/vNFpPrBcjpD88+StTiYdvp+zmGNRHRi+gdjEvwNbRv4Je0Ziu9YTzjjtlnTD83rNSQP
lHDAl16X6LL4JXeKPVL7/krvXjUEDzJyX9tAZA2DNWvDCcdiuqUCH/GEu8W/TbUSoXx5JxpVHOCy
ArhN7qki9R34wR3M5jKKZKbewbtJT9hWn2u9/Bbl/74KxeMHkms922Q1+hglhjcgCqCDMj1/gkLT
Z1FUHcnfqy6cn9VYOAJXOdS4fxZDJKqjLng4w6pRKJ2IcqSzEzuNh0et06PiS7LySqUdgq70ugRt
7Whk1mAb/uZt8vjV9DiSx+9M3e8nv9zWcyYcnySUqeZPpD9geTTBCbVqyea4NOOnaSUJJzwjuf1m
ooER5qh8t02Kcs9dbL+dYODuwCRHbUEbotVQo30frj7dQpZTj9lLFVVddlQAbwEF5sYfnC9fgLs1
Cjq/KeViQgnA3gLCmHr5zAm8Ybo7KzrJpNv/Tb/9cLvXWnvR4moJ/Q4+yoHu3NFQ+R99MNotOkfC
EeU2Q/AJhEr+xxXL8ULA+kYCFHOQIHXBmPPNObGSiATaFbtu50b2Bl1MeYY7BrtP3iNssTDBXpi4
ljMjn4rof0VmzzNqF1CN39W05xZ/qa0SsoSeQWdkAqy9Z7/1O9un7QTkmZmLG8r4T5GPlFhlj8OJ
aCimU5w1ISwbCJS5I54JMKemr/DDT9zFpqpSGo3U62Uf1sPLDUnQrtfQud+sOYHmEzK2RfmvYtK/
ulBzlidEVG57FrOVf8KWJABGqnjq+SJPya5fY2Oh412b4LuenkicR22O9rPZqj8L3km+sy5lVowR
Hs8srqwcaCrCL1My2XLWUQa6n3ESAV43vd6PDIlUeW7KgPhDXGDNcPy8Dv72j7uAB34JJUC639fS
0tgZMYQ6lk2xfRTK5zm2dqgbc7c+wSjGBifAaYV8LiwFt1m37KRb9Rfc7AxGvRr4mjWUvqwhoReh
CT6ax1Jz51qjkwWuJDpAZZk1t7A5gyj4geeVUXNLH7L/j/1GCbXwJJOzBLFoBCpD8XGsmRKtEOkg
W31KjCVKVnWqxrar/iuRvmst1bX7KyKCdy4xaeRLoQHVK52oJKviNGX/eW4guEnBlQaJuDkjB+nI
cIEyi0WMBNQXmfqq5BfP5pFcUv7kIlX7fs5YlLFjxUJCAJg4cL60AJPnVRC1noQ2QYuu+mcYg8pZ
N9aUS8BhISMrUNrq+EP+/Ve7k2yAZ1Ba429v38ABLLJVKLhyauKHMts2PoD27bECQgeGfDH2DQFd
Xhd5kWhZV60fcJeMDYuABlLPNxBtieOgDwx865f+mTABThaLWdfETBtWmdjOlmI/M25RFFhhO1K1
W8n1nUYRP5gWKxqTLa9/0sPNWWEDWvNC2VvvGyq3m1jRMSeKKCF4Pj78Z6zniMt4tV+/gENiaexg
pn1CogFpdAPAfDolKZ4p+5DXQ76ePd7y7+lev1u9vAMMTUc37KAqewd/KOCMuOALl6rZxt+9FHAP
YTvdLsEC64AgMSDguq/1Ff647VCSOky2d5Y2Q02CN/GmFaDtuix3zD/kn/190eepaGVqPz54TkXY
uUSKv7/HIClxcDZqC1+tjCP520NETT+DkrJ237pwKNzxnEDVXMrWn08amMvbhOyons9SMvgImlrQ
OLWRrNTf3TyKcDP3ldfJjPiseXpA97G4mGpmqv9K4sWCZJvoxS+NvIKuD4mQFhDVf2kwfSWYPzuD
aXwKXydmlQ6WAyUIPA83mNq5XE9V+qtrSb0K2CuP12MmMcFPIGbNKW2RqKt4DyC8Oiof+NsAoBaS
RaymBnDabzloJaEGDnYu2Q/PYjmL870cakLzu7fIT5/mqgwuYjesxYtfolBnyk5kxQwEt/vvSlje
5dOFSKrWo/i1U2M8OccTvl7CEIx2dnL/zXMGDP8m6Y5rKucmHDl+ljFmBS/fIT1A2Lzy4NjwTYyh
2zEZzKlRela1REsA1j3kkZlYVG9uHueCEtt4GNZfb5GKpbXBd0rEqJlKypVwhJTo5pwOm3ngAsXf
m5/N6XOndHYqhy4LAgkcspdiUIND1EMvsZF2nAY4XXwfsSdV7RcIBocDG08S+J5T9adao4uiCT3z
fh/dPkmvBTGJWs6ntx891/pAQTycizF/gqoRKd8/TFDk3qvG9wi2p9pAmJSy4itMQWMBZapfACt4
uUqSaghupcIJMslyUM/utsSnqJczruLDCUR83uXFFkJUDB1K1MCvtFU8jwB4+RQ4+3u226QFYOVL
j7EUtQNKdP8h9eJBwUBxt7CDOjuLM/Ir3gL9FtvZ09tczHVlRk3b9WE9QTLO0Ublx6k10PGatbr0
06mgVvd5UzRK83fgMoaU3H1lAnqc48MVZwqgZ7v3UXGcgDAR7hJS9rRlmnZgve06xIKNHWpnb/Wi
bJIHUGG/tRunH0nZ1tMhfraOrQSdH0oN0Gzsd6FE8SEFrHVB4tTCum9Tc+JESafrY1+jX5Ub/vEM
KDD6/SJZuop8t7I3b0+V0t59Eedu6jhYhcDgsdcxlplgFeqR47Q=
`protect end_protected
