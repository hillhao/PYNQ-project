`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ic+e2vwK5Q7PgjSgvwMH2WoojQ4BbTVuQzxkOMVjPI/VZ5NZbfo+pDZV2xAqhpQmyQ9GvI+HXb1j
HmlK88vB0Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EhYQ5ehP63YE16bz7Bs+Jp6XRtGGK+uBxpAwDXHwR28I2BtSgb9ncXucOpIeu0UTEMLqbvoLfbxU
MKaMrYPMo8RM/a2HDSBr9m9kqrCswhqrsj7+l6YpDAYmcCTq9T3FOkfhQRKFn0OQ/XIIbTvvITnM
Im9Df+3DnhnBsRIa6b8=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h0YJz7QAV8KNys9f0Mxlf+pNNU8LPo3hH7TmUMyrhw3lSO+kM5IGhIhrK6tA/vHS9HjpGQeWP4CV
hUv0PJuDbFRDQozJGwYt7sEJSKD17mUe+oi8D93Qmbv3URq5Gi+VGUtURDK7m9vfm75L8tyy5ql9
qECsNvUIWukIEumtJEY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pP+6eQFqDiaeKP3BC0Vnjvzv+UaX8yu0QFcUAsHG6nA3D6UEozm0SxdJ2iFfFcGPTkGK1rJp3wQa
XKLNY1k0r+8h6/HdEgYrEoLQxiu0rGTrMwFGkm5IpBA5qyUQJ9BOMA3RodmPZroFnpuOiQG9fXXi
E9pTQFAqbQwJUIKn68iPFrjVm+q4qLqQgrHvjKnf6JEciMX/HO234NTOg6COPSv7Uyo3FXOOpRHp
TCTyJBrP+6/0PD1dPLxzogieQ1fECqhCHlBWg5ARc7Wy8Nrvyugiw7tyWe9OCXkF34mphNHjHAfM
kre/l/mYmZh4jzXcx586HHX8Gny5RYaZ4KoAiA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DtRivEEQldRL8LC1umq+yZAExH6mDpzyWG1k5T3n0AafinwOAShYDeN3xJBVTROrx8yaZtcjOIVo
RTz2YCioii4y47KGQkU7qOYGP1IL16aZBaLHN0ikiASZGuT2wIZ7vBOHDkXuyg7SHEzSut20MVdH
yT522lI1hnAfDXEZagb5qrrQxGlsFJtLUxTUFbZ7CLxKt7IYJNSHgoLTaurt9KNyJHnk2Oa9efJx
cG8KJwFEfS1eHTBu0rJX6eoLGEyPSJx4qXZ3eGjOwHDiGelueO/b4BZB7QA7g7zVJz86kqUZqX1s
SpXZOqr7kFUwCnN2dJO5bhUtoF+y3GgfGerZaQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pemFOX3XLyQdy4vtMYjiFXTZP+XlsBGKuE92WyWU4tr/zi/kdVNH1ODTNxNJ5DXwFjsQE3XaQKcO
QVG3dkRqyxkufPvrynU460117JgXGW15a8rem6Dsd8qn7VgNRECRRwFEFLE3bFhFjG5aqlEDnd56
Jtv/dX2cI0okyfMCEOBuMBd48KhjQsDycf7KtJc5LpL06fv+nYIvBQGKfMIkl6F4N9MkpkCF18HN
sm252Xem8SRCkTNQW6+o1yOVN45d9b+5a9+kx3Hc+5oEfCtymCxxbWIPnLnMAGhORy7lTFlrznDF
KTRSVyP9INWg2r5KEz1jo7u/eNIyiLfueJeDjg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 962560)
`protect data_block
+93ue+0K+V+pjfzqa5MG7BJrgXiGn4kNdRfDw8+yn7trEE6+JTDP2j1T58WRIxGnjWDV5RmoMP2n
gfd8qKQoEUZqHUifneZsvxz7zylDGpA3dkCdCq+LUil9bj+8YUbj2Bk9B972JPidpTAHBZIPTykz
8KCHUzcyOvqiW9+leCtXkFYQTt0Rn6go6AOk8tl8tbUFBynVWRjXPcShLQv3O52JxspXGH16Gtq3
CE0ca6FK8AFh/no2nhgPI56STKYapVl7a89ubEnYOUAiu4lc5gvXSsD1g6l50JOGobHvopb8TbxY
2UbceEaUUEkPS6QbYXvUqn/x7wI+Kd/hSsgjvBOkcyU5HWHmmLapwnVx/OJG4BeimfTf6diqiSCA
rerdGxgU2ICihm2zfnV+FaN2KXjJEkDdkMsSTfSQh9fOuHB6ATldDnHiziGEBnbtZ3Y7UivsqKRw
mWLL6u8tPFSudv0UNGtAwLTxhtt5WUCZnERNHZLLU70UWrEMCS6ibvlFRPB9l69a1hHcshlLz4LB
abW3c3HUL1ifBHsZtmcrMLOrsEiEOqWFaD7/hnVPEoGJoxzTQ+TtpaLaXEw8vuf9Xll/t7cpI7NI
LgRps9ZrofIkPE+CIRH3ovEzQJKNgvW3OiUURHgBm8XjbbAbNYOcjFsquc2BFif9AU2A/bSoy1a3
GOhyPd9PJfGeL/1SLRPHNFSSTrKGN6oTY+rxecGF2v7T8w0j+xb23Cpc7CSSYu5gU1tjGG+u+ZDU
muZfME34ekYz+03A/KERtKIuO3mtus/GAw87/ajbJnX4gA02KQNCX5HcS1uCpDCMwgywKPWVaqE5
e7O4p4r4nvk2w0FY4fk8eAd98a0F/TzX3DwX3GNSozcvYqiojcptX2RlCVpA5VFXFHlMnQtgi0S2
B9CdMnKkPkCmJI9rTjAJHvpMV4JvFhjuYcCgLTY+fWXIiDICyx/W8Q9TtTrgQGK4mjrmgTImIyVC
/lBPLGLTy7MTWBYZAvgNRZC8sNR+xThcqjdRrOT5u7eBjRVx3OkZ9Kk/MhbIiHBVJ/iSbP5+J1Dl
HVNCarYKwoRtqcdE6TK3D2I9Hz3TxYzMX9mJ6HhYQ153Nn6qIsIpHWD3SKN+3kIESeZUd2jV0ksG
lH4wKraAHT4QRZ6aMXeJ+h36Vb6NtLaJi8uEOoofLGGb+gaWMUSwwqgq5vMv6kP4UJzVPld6jmJk
pIbRdfyBrc19bJfzOp/CktzDF5YiQy4enRquX8PemyxSERhl93xSENM+mOeUvMRzCtOVqKHeO7F+
Rhvz3krhGItsSjc2W9RC+BZIzjHvwXQpWIhXCFjWLWbxvY07g4Wb2bxnP1XHcvxtxZzsD33klvm8
ElfhKej5KQf6uPkWYE6nk+goL7DlBbi4wybYsp4sm7o27Fi3VE70bbgsCSifHIqg2M3GlLreNDbS
wEjKr8SDUG1zeVTzZgr7y332V6pYV1d4RAUGWSkoaf2C86gvLG1aQhDFYZYHiJAWjFBtHOju+2zA
dgho0A3+Tep6KJac16/e4ihuYdbvLfA4fzIXDWer7YHPCGAQNer44KmkgHHLlH/Mm8cTtCQo1Tm5
ncT2KzcbCqlGxBK9nUQuOhonOpLgjIO1gaXJAVwHV7B/CNpxjlVcTSUqBngcyVqGn5vMqLsyDbIT
ek2Mm5Id4DNHMG/sL8UKpZVl6wEiblF+o9Q1NqNcr3q1anJASoC93VYbuIn08ZJCLEn0mP3U8yJO
EbNXRtQYJdDDllEXK1/2Adgp5hPpWjMG8NSyEojnisHpOSYSFA77LefQPNXVUD8l1ASlcIHd1Y/d
Ycg2JID7FYSZCSHbthBHFlpN58xV5wA1J75WLxqav0TlH1iUR8S0aaAiHXL2goF3GbNAyXtPMq+Q
5zCVxcG//ZP7+j4APGV618AO9AJRqHpsLaotZX13qCc/hZwZVqAuA/1hM4oEewK50FuQURtURoJV
tl/1yNoB4ZQCf948tb1EvPx7d5Tw91s7bG/dC1+N5b5tAcUwlevx04YjjuF1H4fcKf17HH+Q0q2b
eV3JcPMH5D0vHwpiii2fkoen3heIlFWbC1aOivkGdRR7PKzO60BHeU4UfOQS6bAzNWqjHwcDgPoE
7f3gBkl0e91xSZY4Ci471c4Zx2awE54jvn9A/qlAFXUwxocjHATPjrTjMdWdTWq44h+fGHKP2KEB
lwBLoSROIL9KP0Y3Y/URsyLAy/jt1EV8qzVKHL4cabzjFmb/bOJfG/qn4ZP050HtevRz5d8hZbIL
HtiZHVqxXRweXLssjRUuZz66jqazeUmCwwHyST8o1JLpaJVg+e4+buo2rUHp25pxzyWjsKw/t1a+
JV3EbPSxM/OrltyCursKJDCGV3rkir/ZO0IXHXPlgxQ6otxriyWZK84qi8TC48CUxqOk7C9AJjdo
8CRNFcmYWPuLmlrhc9EHvzjcaAZ883b401La2VQhLmiuMpTmHxM0MfNJVDz+F1zn65fL0vSoqp8Z
cNUUVbFp9hkU9EuM6BNbEbErpCRoSsUALm2TNMkUxx9VdWSWGiH0ND323lF09Pp8oYtMDiZ+JLny
uOAm6YfQM2yJ5B4RQQPQ/j9xSswWs2yJ5WQJl1BlC1z/E0TcwMUYc7y2Jf6qP/P5Obp5zAQfAWaI
2DWAc2NI9PA6UgTwtprYE10m3vSKc7OlAoaeVEGiZB51sfJpFQ7XdpB+gXX3yZEaSCLnVpC6M6Gq
U+0kpu6eq3zo3WjO4vXsNQWyOV+OAJsfiQeJIC/HvXPIoEd6yUpPqzUGuYtCNXaWDZDXj2jJTbp/
T19UQMwI6sddQb0KReDqsnyKbZyZ+dmQy08hLDMIscymj28pgn4LjZV+egnJyVjrv2nD0tce9uNe
OXlkkrnDIgmOg9I1QRZLLFiBc/n0LB1ZWOF6SkzIfMUD0CH0BuivcVN3EoMsqiOSvlAw7IidLi+E
5ZRXOM7z/LqK7ZQIOoOV9ng2R7T2tJGOMjeOwUu/a5tcKuVKkUHuA94lAMgsZyNEUpGW2yLugCNQ
F93Zaax01KKP+x9E9B2I7mgaCJZdi/xtgxPxrTHJBwg0Vu5IEuWN72FNq2hYwNoeeyEa8UcjE6RG
qVMOoDEG4FZMZqkn8n+4Jzp4k0BgBbSm/6ytQ/UORWU+NQJ7UF/F1LoH6Eqegv6JgehbYmIgrDG1
ExvLwsTV3NhgFcRjMFNJ06iBHdiEfsBg85pzGutjFjgQiyKR+1Ma4mVHhp4ZicSN5nGS0q2zN5v2
okcoaByBL/4Ciyc0IQYCDWbQACoCvsFdLBDGm+mgEgx7g9uOC0iugxbFPFR7i23yvZ0q8QY5k/sS
J70VyWyRLI+iysYvajt0up1rG2K1JlMkxexFEVkxf5UiW610Ri3c6kS9QNejoAWLdt61OyuBGsFa
8rHNiLTyEAQG6Gisvvl1sVTRkBurNmO6knCRQvHyDhd4D3Tw3+qe33Mq0kWSAgFMbXdvsG9S9jaw
yG5VY2kZuBiFwf4kSpmfK+ES+FVkTlb94rCPPCgNCcOc4ScL90a1lfDVmUSjXkOnLsVGnAuxn6nG
nY1YsR6KHtq+h0wao2TWmPzOcq3xOWRyCKll/4ScHIV2OI4fsMZrYC6/SAvXTQa3CvoxCC95NNsL
vD0b8dWP6XM3yhlzskRi+7qCrwPNSB5P6pPi6LqjAHpuYznQ9kzqurXyLXm6z5Xx556LjmekLKCX
rZY2/MACzGt8ojSHQ/f8jASkK0c5QM4XV/FNV0FGoDeIDeE5PiTIwGxnz6IBB93B1SSqXgl/b1nG
PQYZjwQcfkq/ltWGsQxzuEad52T3wgAY8D7JOBZAeqtS10WDUqO4YNVRAWbr/SKQ2Ea1lgLfwtGt
z0Nycdh2pEWdZgXdYwrxX2l1skoq94TMLZukx/GB6d2BPFm44lycaSq4nmmh6R6IlOQ/2wUD0T6Y
BTX0v5itPCddVi/tXF+OhvDZ0c0nsEdkCaZMZDDnMeSQQzfwCuoTP18Rfl00KHrnRseO8nEqp98B
OLHv5ZnfFx3gjN8lxUMnv7ZL2sWIA5Rh/awB0q3vT99+cvk8JLmKG+v+1omJEGVh8lAeGtlXMhhN
W06Jd/3yoni5fWhSbgkMGjBSqcmfMyt+eCwCU7qFZOcsy77PCIUOjeYjfpHctZlg+3GmNkhVGISU
y2VPsaCPD8KhRNMabPm0avn3zda4cEQLq57FaHVrPZs39FAyNGOMIZmDbQ9TPtsNWD0WP68bbW1K
C51yAy1LH4MiXb7YHao3E5+bF670Jyg51CkwAHUSYQyo2C2k1YiHJspIWJ/xKXlJ3vJJeUZAgaor
83Gr9nLr8BncWd7lEz9Iw/wOjvTC5FrR3/f5TOxPM3D3jY1xTWDmYAZQIspAMFTcsiV1zt3WVZN5
ij6QoCbIEsJxgP4lX+g1F9xZuhwVAatEjAMN5WSsLP13aFANtX0xV0M3HuwZl0CVRWBVyxLR9CeL
55vW4RCxdhnT/AgrzEXNUVytZOXesYZ676dB/p2jqmoMy89HWowaCB5C2kUvN3JRqCgIseB3TTwB
kuYvTFU6gc05av6/L7R/KtcZo7+XhQkw3eHRCWxHUOQ7iUUUEU96111hmmEdYDai06XRx2WNn3uA
YvWprX4kDDy99LXeexgulszTBUrqRTnE2INxFNy82AOjBRYrAglFjVj1D3xuPogiG22rg8GjoH6o
akqBC4Bim/3K9yFbA9Wtb7gB4xcO6MhvWwYknBJ+zxY2NdJ5D1QcDSgnoXAnjxSMGooYW07kE0QQ
lxz57H7B/r8O9WyIhREJQCtzA9GPFp1amMIw94/QWx5T+iJZSBM0K59vlIIZYYdnflY/VUP7Jpnn
RUYztKSGvTFtvkJrJilbRa+OQZpZCX3CuQuoXFstQqYJ+crTrrfA5+mQhYgfVdRQkJ53SuZWXgnf
FCD6hROOrRRvUzwAFQ5OeGZ/c/0whiUTvny/7/ZkMWM/eZh4cbUyQ8/xW67U2BbraWrlV47fHiYN
p4JOzTzzaNthmSCBKI2e+TbE6e/moeOQLkd3R7Zy1TxR137SaUfU8PGXMZQQ4pCrj0zDeAELCmJC
ugxQfUkDOQYRFTLUJL5aQG1P/9etinM8vzc035cPBYU473hdx5S/W97o6VzXCa4vkdxZAS1r/q5q
5Oujh2/JpKrP37OVJD1A1u142Gs51aPYfaApjUObNhtk1M52WrjtFuNeDo8mYUDDF94rSt4ky8je
Yvjeje63UhtwtHH6M98NfPlwO6N7v3xBaj5uubGkDyCcCJyqrq71Vc4KLY8yqtktlUgZmimk3pnu
Jqv7CVlSA12XLitUidsiSeEm41M8eRVdWKRODOEg4vW66/OlAmoHgXuNbRdkcucPbkLdRP/4zKNh
UA7mmy36VdKQNXaWNxLgPIjNQTf+lbNaI5NYcEsAbnSrJNXdVjoDIL+xx5CFcsVf6H0+9VhuhxiQ
hegMX8TgOSrWL4did6vSslAl5ySboggRRlszaSdn0XA6OhE5KdNB5xPPOPmESiNUXI79ppVpiFbV
MNJ4kB5rzU3XRH3Hk4aHYavVw6vogF6//aeIjxlVEHpSPTDm/WJx6D45HIZHMmu4BA5FkwKbZPKs
uEDwQvI3waSF34EC5Wsz88PPCqueeVE8Wy2dSeGFqQQXQ40DoRFg11EARQb3cBvhT3R21jJgO9Kl
6w1UPEPBuHmEvB/gJV9YScdJHEjZgsUBP7REK3aFMfWG8REhvdMsaw0VtgCUBDMphxXjgQNAE1O+
/r3eWoearPhsLR7nClSMREyFtkoMsNIOXsjSxUR+O0Irte8g9lgZG9YDEgxMi8ifA0nOShE90U9M
HbDVLY/l3Ma9ZojzlLXVygYFK1VYPasxW9pqqpS4GhJBT2VAkF0RnOQ3LryWtjAoCcMIDe8Vvni1
PxmQzjTvN4pYMtkX125emZLy9eQHEbTv0ZJZ9+YiG7/E+1kRNuIUKkHjtiri39RYXtQB4X4ZiYds
an7EyIK3Upue4aM034wmfWMn0LX+OphvrMSDP8lzrnEd+ETXwopBfuCCe7V6/a7tlz3CsPYXu+dZ
+IlEC6inp6Xh8hoA0ypRjNOgle/cTc/OvUmW64h0MEAysC0iAYYNnBuTQMlSSpq+ndDFXiNtY6cX
8JuRfbAySJGbhEG9AXUm7iRjNvfrkUoHQMATfKFZ9LcIxD2iekisyu6wNTdfqymKps1qTnlef8bK
2Qj3jZLW8Bc9HHmluA4A+9aWlznk9/CYj0lpbxhKd3SsiGibvDQ7hhdtMpK8TCKnGFEwz30JXmNp
R6wCzfIj0UKgZGBO20nKIvXW/g6Dapmnr5gI/3Duefg7N8jUDSWg191etRRPUbSneIwzxHab726b
9xsm3j0x0kzJU42/vBSvtTMph1NCYjoWzSeP5mO/3wB6xE3hF83FIYm+/sJn5QVXkOoTm1T87OtA
cyi26YuAF+2U78dgBQpP404FrT+cP84KxFZMkQ8fK5qPw4KxfB4cWoi7ntd3aVoFcOxUYbtY6lom
HkdO/DBa9qZhmb+Y+1oKL/ueTsWZspD2Ng3lWFEQ5dgODZHjNmliFWqNHi8W9pX7BkDPjxYOqbDi
ZLlNvgZ3XnDgEm78hvJHARCqeo6kPJiMoaLGkgRQtGNei5rBg8DjwxSUqn/AlU+RfDucltONERKv
v7F4+Aar30pGsKEXUZrLwS8jiUuPllrcNvOjYzVMMhhJmsfwywaio0bS8QN1GlQJuAMGoBXHRiVa
3oSDhKiiwbUzUoBI5le3rEwARkJ+9ZREfVefnyGokGMA5e1k1ptGYc+r8gKH9HsDWo6x6MlUDkrT
btpB9DSFU9nCrLBOILlfKrgAK1f12vnJoGkbKhmGrQ5PBPKIgpueOuBnN94jyMtPLOoQD8Cl14O1
DoC0H56T9mG5RQ70mlQwbc+aXDG5pVL1amr6QTGs0ToSMW+WLKUfGsWVF6wx2Q5yf/6GyATFh48Z
15yeLLXaxlUSGIRDeJhmyDaqMiiw9+uClFGsjV2Hn3VfJr24LtOYG3gPc1mfg4NTZ52qX5n9P671
g3a8oUQ+GBf6dPfGEHQPzv6jTJDL2Rs4f4rfIJ0+kV8G6UlAFN52oBp3UxCSGO8FbT0Kgf1wb44Y
OxwQO0Hmr7EjqY/Ca4IXrVBM2jNu7X7aYYL/fYZPhXSmEY2rsTWmMwekpWFsGVVAZJMzHeH+zqkK
xB3EtzUq4vliV1CXc1j5ozHwTP/eRfhdL0Y/EtbqdN+XC40QTD6yZRwlUG0nV0o98djzPPoJgWHh
IElThdrv+IaUknY8spYHMdFrjWzSa4Io0AkPUOjffA+bqpQx2q/T0wzSK1blHajZ2gNWKtnKAykq
ssTgtmhLftGizv8CO3q6SDanXcIZYC15D5VOL5mnBZzkdnGP/pokm1+ZTsztAxxYh5yTncnoNudl
Ugr3FKaBZ6PfGGac5v6aCk/Z8rQ0JL1GIQkA7k1mVAzDJ7rK6GbSV6G0hJrRSXEtX7oJtjopCkAk
HXa6AUoMixeJ5Z22XjdrWobLSO5jfNv3gK4gxocOyb/qwS454WPH9E7f1PUyhLaaBEKG6j+GC+OU
o5tyc/AlNgHexkual2Ja6o60HYIKKp8kVKoguJDVXpoL/cs2MuxmZJjlfFBGx0YBEFjvYWKXfF97
0xkPt5HoVxvdRpKYukEfVwjWeA4XKVudRJISJJk1d6/TEfBH38rO3qSQJSV+8RizxBSQ3XFqWVET
kJp3XSUtH4h+5Gx4OjyygEiGlHt+pfQlnt7vcyjeo7gIHJQMzCo6KzAbhf7AcgdvX+DqSNAk6HHg
Fu6/KFsEjbrVZLItRKYrWyquVtIblrWw4JmbM5d87t9opsM8ejc3rllFbYFXFUz6IHZZE4Fy+Ftw
76Iw4fAtKH0OV7sPVt5cQtzd7IvsFUOWr31qnbs+4iYhVANMXkKzPhJu6ke2snKAWoa6IS/7F4em
bISNa01NHyjVqUCBj4y09SekqJJK7rcDXb9sdzFyfRX74LK2g4zkSVnOziPOppoWTSb5Hb2iXQ1z
Ho65h86vF+HK4gsN2UbhnxtAVdIsifEppBiDciquTwddY/C3PdCNJQiIsGcCGHxPjXzl+phzorYl
HTv/scbUaypiZGY2mIydP7BAGUOzMvt32chNdoNTlD85SvQeKLfA11JVuzorOwcpfs666oSpVW5i
wT/L9CkeuPZ6Lt4A1fuy1g65hfUhdhxhKebV+gbXhKxwik6aql5uo8eUz6ULIeFxFXI/5lc8uXhf
5rGy8rRmxoWsUX4UIdlWVpFL0mAoEL0bwmrtxPHuNv79flVqc7BKWKUnoS2CmZEDK6wF6aap8UEt
jGcYM2ZE6nhnflvw8ltNfkHv1jlHHC02h7Z3AGBq9DnFxXHP1zY0y5teaXq/7jqmNRMx3qvAWhP0
MrrcqE5EDqsdilhwg5jDrsJaQhbrgkdyiWNukPgPi0rflXs4DgyKXmFhXjruoDZvCGldXngu2aWp
nPN9PIcDtw8xX9tGkm1m0g4MhZVViKWUW6ajnCBJg+/fo/qE08yzpxx8uRfWm5Vact6QJ4iF0h+i
SVG9lyIORzUg4WmKZtoiVOvIplyTzFe3eCTcXvdT9w0QTTDs6kR2Nwa5imOT48i216LNcEKCGhSu
oAxil7aRcdeNo5dyFrfF+1FuUYH04B0tL2PV5Gt7D9Lmn2q0VHDpJXtrmBJDHADE/w8TIMyTYrtU
ruQwU1DPx9cpjcHWaE+nd7NMEVCOWGvG5BrBy0ifX+9MP2O7qmKLycC0ZH+Jli4TwFyPYy5qxBTo
vttGsfTi5rdld6d8isTvC2G53K/OMP0PYG3WF9oViBxtA8PoP04fd9zfY9yoiyREfFg+K9Mr79xE
LNMIUnucB5OjkmpOomplxjn6zQyYhW+RlurPgbmDLLWy1wUG6wwpW99VY7l05MaeP0NB1xl88Cr1
+f2lPC5hDMtz+NkXRYJUlvBqkn7L2lM/QZFPW5FAxCWOGCHL57F3JhHXa8Pa9Mprz4neVu0g2gSw
FveDQ1+AQ171ZqiEV1La4TYsYhTWaVMY2mdbBwympMN4Gcl9yusAFL6/EV2KPx/CPqBueXqWplO4
zbGRNjcM1sDwnIa6OUEPYxw4/z8AP1xeXXNFMl/K/D0ee5lyvEnUzOA4IdzR3J3DlJ+6+rHqFtkh
X3mfEQqXN7Y71/dJai0GOP7302dX7p+UgvGsBB6qm6VLjIYzaR6t0zfz8q4c9DYIERSo13ZH5yOj
UulDDiTcMKDcBSG52z02SnHwTEAA4nxXCcVUKSQicnJ/0Eimra0+rDOp8FOeE539JLETUk3uEPDL
3w0deFJuU05KfuBPKDriYOiIATaQ1b17BPKYwBWcmgZ+SycZKv917DhqaAzj7nJP1rOwg2LE2UZx
z8vPY6d0EWwZhDNtk8ANgqUy1QM8z8tUFbPTFZCyQwpwwxtii3BvL/zqcbXtjKkL+m3nKqrbdOlh
FwTALb9SaaOKZ2YuTK2zwYoLX/q9OupiWuAx6Zmwh+MCu1GlU8TS/gbLipjuEDxUct5sMiNsrjae
/9d4kLHud4915kYh7QSc88MMO40H3iowI0UCu22fb4DroVVgcR1vnvX0Vkt/RNlt+t+vXKGM9XPY
gl04j/W4tuLiTPaHwPfx9ln3qOzt+lWHjt3yvzvHs0nLpfmZygem5dvbk+B4qAleBTXg4M5TnY+U
zH+VcNcfionral86Wwcbo9aTcQymwlZMtlP0pQgfauZEAmKFrUUwIFmv9C67/sc8xHhjg7RinHJf
Ie8znnW3E6ZpJyXkH0zv+I4814fbj95YW8nU1Oe47kntv/stZLaUHd2V933Iy+tYQqVNVTiPDkgi
K07cMaJud8YB4QZRWk99F4SchXEtkZ8II5ZJA/pLOUub9HIXbnf4xt4mjk6q02v+xCmRpVFa1o4W
Zj3EDOULXH4qkSML2KPP0tslk1KQNZxcF+yaFs7HlDUq/ZxiTAInTQ5NJjofIZmNh0zfPblt6gjl
ZcmhWTQ9qj0Iy1NEy2PSQK1nnPY7Dzjr4eyEM07xgsiHkrOIjJkopJmh34ZlLaYTqqVEjCVnp7jb
pG9MXmTRCLZGqs+lQ3L67J9KX4LRmAoNAzR1sZcRboTFljC6Ob0EFmjvlZG7g0yOGgDZeH1uEsuA
0cZZwh4zvlTXYQjHLt7nMfJ7iDGqiNqpKrWNlXcOXNsfBjv74iPQiTJyAwDty/BFl2aA/0pUw9NB
lDZ+pxPF78VI5nTLUcn8dNtNxCBrjS0bonftL/ib04c2b/15QQJ4EBTh09SOinVwgaH4bRYE1ULa
m2p7CyE4MFif7m8qlfsx+H8OoDkWS4O6kXy6pGQi2HPzgeXZ2owtSsnQFQSYiYLlYOIAivdnXIW/
vUyF1pQiHNmtEVeBwzYhhGbPfST3MPB+CGXKZk2fkOeMUpXm1dY8tSuv7SEaSQpK3xC/R4McaGJK
CMz0mNkYW6vXH08440sAS7AmwCgKOza+jAwmIJoDyAFL7OlBah1Daco6idWLjRC+Fq80XI0Pu2uk
0EmPfGXCkG8Cs7qEDrX70HFpD5l5mVYCX2cuthJBsRNJlsG1jnmeAWbaW016G3ikyJ6fNlVWMi3G
PXBvEXo7bEQctr4bX/ePjcnIit5R5H/9frEabE2V/214zumiotp7Z+W8/efiWzWZfMOY/8eUv6tD
cPPcdLVENJt6VCGRVFgklYxebSqZ4T49glKLsJiu/LK5+GqUU8er3ptvjSXkTj0qIKs6dxm8YMOH
TDhq6vv7U11nSk8lbCBNXTmaS4irdc0+H3XUttNHcMcErOBSMop8z71mR+5cldCGes0W1EX4Kfmt
DvBeSTKfd0Vb8siwK9+SOKGeqa9w8hx9hi0kF3ks2SHNG0imwRI/A9Uitc/CNPnsmSoDjPwEFqR5
eRhHghMf76VPg2qnr15KYWSFLr5+MvI/Q5KSwwhU0H6lRl9Kpy9MSkGeW38tY2VOz0iAL5TsRg06
Es0iATEFzZayLJ81uw7LNmtZLAlzHvn06D9s3Yjt1UOfJQkXQPk/69sH1kR+RvoW7eUu+kfN/HTh
J/BTAxYORMbjHRxImOg2IV+dGLSy8Oh4+umdxxgn8skxG45lxPOrN3hbkkXPODBH+bJ6bQcKz1Yh
5HP7b757xbKjYmr5SbaCaG1rT2Y5UA3LdqSN2wnXhUBuyh3eDU1QykiUua53hUQluvKvKrPSmpR8
5XOiXnI0FU96HNK6NX5cOPFVWxtFzJ0G9RVgSSp1662fqOoG72RoucYVDES9cQr07yDW8t8r5tJo
cQHHVTLntKdV8BnsOeqtigTv4c6UPCL7T7Dn2aQBCurTqhg3dyd3KjCfkVOBcWCU8iLOFZPSrjE4
6RfRn2Qcun2R8gj3Deo4XAXBCJkyV4mhdsO4T8e4XdXWNufgVbttaHpfVWxmIMVoL56wCrxvBEnK
GQcmYv3Gu2UokVKeN++D2YZ8ASUmmC06S/Tu7YLkJoNsyteKHy+Nxf26Mr38Kk+5aeBdIZkVGUNy
A09s21jam5/1VyvR1k/91NUljhNJYRlsVrdad6DxBgEG+wd0BF6rbGDAhM1qs+fIG5Ya+Ue4w3T1
s9IfagEgY3BkurmN1PSO6IIXkO3b4lzeFESqWiw5tmbT8hMP8OAXIxOboykiHJ2/YjLuTcoFdmhM
NF+12ic7aNTKv88WO0B2Gss404M/wMpLK6d9YI4mm4MKBGq3HN+twW9N4VLyGA5D4JerfaMDbDK2
tzjWCDBUnBLbXmf7TZQQ3T0MOQP3AONinj3CDTMdgxMUUWWVZ8hHE0yuF6I6ghY9CFfBD6PAC928
5vO9cFen4kCewCMkNoXrm2lR7b9tXSFABfRzU/02R4S4cekgUIV1fo5aOoEFz14ln+oBkjwtIiIq
WX4lYxxHITpSXPu1hZb6i8lgqRWlXU1t+m4EFoCfpyc47rAr5FRfdP+DzoKrNtcXWAvgsWU75S71
lg+xYpJCiWMog2dzDv2qfldTmilC9ltbIIdRDsddWVfkxsUQIqGaq0B1Ye+Im3pBwZwfYRGYtlzE
xFcfLkTKctzLWITjcIuq2B9e8fd32bvFgtAlAqfPvAkR8A0PeYAWZ1CDl/lGw6dJ876HCtfvkuhF
drzcudsNy6I/htwrrO4qLHCRQF2jFTRmUS32xpEWD4RBM8ATLm2HWiyAoqDTSdI21U2qDid8UWjH
Tg6c5ejYUiQRUxe8qaT9nPQPAbLP+FVNZ/u9RTuwCLlQb8HcdIGlCt4wkfnyptTkh9TxCKrYrlxB
kl0Eq266wcLCtT4eRrxmd2XoRl5Szm7BGIbR7t4arG3x78EJlZvZMnaX5IieJXkn5frIgrP3pY8y
uMK2ejz9goBrFrj+zn594w89v513NNsBThnxKAwSwetQZA2wzFCNggIJEfitoc8lwpAJXXBbzrp8
UnkWsr3Bw6P752Fj/4hyrs32fQQwGZP3diEDobQ8nv5Glu8zcXkIlCyZClm3BBuMbQSMXgt49wQu
6xPd/kduCtR8FVH2MJCt7Omh3Bydq9lrCrSBBNB4x1+8IQPUajsHlUvpNUptatAPMn9IY+mrO7a2
K1Hyw0ZXxgCQ+2B1R8wZ+YAvGdl5yGMAdwEBX5ioZqQueSrny5NRtO9UsIg49ScAl2mUTtVkBAk8
sjvkkW56k6EXWuss7h9ohBv2jitsGa4VMI/Qtqm8TG9LDswNwdCR8sM/bAK90zxvwDeMne7cv+Dh
0xzg4jWpm338+2cr5rL848kuO5DRS8QJknJrABEoJFry7XW6YUiUkm420XHfIDM0Bc3WgMwytxHD
AImPKsHJjXdVNdRlEzIPqIc/YrT8UPtmCC2ZosP6N/Z95bBDvn9Dt4vs1tdchismVhz6Z1l/81Qz
kEseLPDPwvzaodAxn4NZJj/SrTYEVNbYMODb1r8zQuw7EQAM1hMrdXUgNC1C2SbTDVwSsqEy7Y/v
26pe6j5w7Sv9BZNNrgGoKP1vxWHhdKn1NmRJWC/LWDFEJAo9NE3h+8obUgef5c66Jo2O+mxLic8n
gsGUtPMnMnkjyg+WEe2iOhjJh98APL1q4tM3KR83ANB1cRuZvRShYCBuadTzeC0iPsOJL3gm84WJ
fYPmHhIblrIdV9mFOx+Xmd7rZpkQtOQvvDibsn1mb5VOE1PsqGHk71IoeH9ZB1TTVI99/qlM+A6z
7gXeDUnaqYRV9XQttm8YnFpNfnKOwvAG8SRtbizgGRqlNZ01o/zvvGcBelUQ8koBc5uVT6eXA2BR
6ajfA6kVAg7fvhpbm830E5wgXfHjGiUNJZjwrVd2BhQT3kCedKzw30Z55jzkEIhMOJ2Z41NYZFWn
PatuU15slhK8/m9C8AGnhWeYJSDL6+DHsl80jYsptetQFfSyYHUAS4NmlZS+PZvvTgvY9qKm1kax
uiBBeyG8Us89hTRla+afzilEuWScWvJVd/nDdrtdud3H3WvB1ju87PZNFd6OA7u15V7+aoInOyTr
Ghl5Zy1uZamz1E+y/+09e/Zqi9S6FtxqzQsjA2eL1zi2qlMpbl4c7wLFbHPatT4r7RPtbi9ZdF5n
OQHzEmLLvG3OPn8JgPBA0Lc59PMAViC76jlNe0Uw5qPUR5/24jJqxuS1IbiAN4ejFVmRHjRxVqsN
D3VMV3TONEpqccXU6EaK/uokGylb1wYCQ0lMt3trfTzZxX3MV/eMRecfPCZYuSY/LhYIwn05znyU
lPS/Uu0yi3EdmL0iZXchulQ71jZ1k7nHz+fRjDDAvrGuEppi6Um6Nxdrs6vwIpQSfF8V1sunRLCq
ACznayDkisVozrDIaxuO+ppcj1mfaEUVSSYrSnUOtfTUx6qjDugcAyNR9e4mSe+iga5MbieqV0Vz
aIV4Hu6GoAKNgyUiKjZ1Ky2vHINYtRnwRwCPwvORXr3yfCFcu4WouiLoXfDibKNwplGqyd/vB2bq
9SYz06zxJEiSXRClVbRMcbgHWj3dXWIVi7mZWINDJgKylHWkE1vupYnT1+yQn2qCmMGPxgtFY2gW
hFw1oyiFMfCJDy+MntzUTeDlih6Bn6JmPuRbLVUVquwudB203bYgwU2UaJZ0vwZpW2hA9/zwH5So
Jdbu6FjTesQAu0sdHefMipf2ay/bI/qtxk/us8RjBM1I7qc2tsG4DUEQK95fU56yBRu8Cl/b6krQ
ooZVnPCcAjEJRiTsrnJcVd223SJub7pNtlG3sdPTHssxr9MRyx+HlS1EccZjEIr2ZZ5poiPdpoge
ntV0NSUxWzXh2VCZgQk0WWv6IjPlZsn2PQmDl0oVBYFpS4VMWk2s+OgcKq8roAAhJ6yEVGEQYPPw
EjNkpBPnCNPAbLz0DMZL8jqqqw2+1JCVq/IXzWnZsRIqpcYrhUi4AhIyYTYamTV8a5IrSkMoAshK
+ZfvStUL2yRYLxInwHapiEgCm1Ks6N8ei5UL5Dpr8rzKv2GlENSG/FFTLElkjr0HEWoo4kvqYBli
fnFNsvMEiVQwM/VJMBXZCpwYR5tBoMYYh4AS8AIYkS2aIAKqPSfjPMTkUoOc+GXEMAbY26Mis9mi
kNi6L50gaCrBIXxoadiUvXwruWSIUtuKNWICnOojafSDTd8hUocSOHx48d0mFJvZMBKwF6eTVguW
SHmI7cbNjmV8yn8l7h8SGwjN2j3Shlws3MK86TRomtpc3hDg5WbQ9v2WRSpxNBFGCGPR/n1qkK6x
hkcxst+ycn6+TQRGNJVMNQYa/TjJWouLVupnBQCEpGvUR8Tu7obXkFNZbHBn9HzKmYiP3vlR6/s/
ueAMhGEXzqYqWD00Ab4Lk1Fjnw0NNmSt67n+8fcsa6ga+oYZddu2j1LQFbZeq/QIsPlUQAbybcN/
tSYru7bkmf9EceBzEw7Q77/ry1byVro7/Ly0dv6+qltrnZxCiIImt09XXZfBATk883VqAyVTE8g2
ezBQYzgzUQ6IGf7CNtPQ76Ee/4Mhx7ZdUX5v1a6cOXeEHB0FJuViK0NabcHsBdarsQ0KQhBau3gw
W0Wc+neN8h+dCUAowZcaVdZzVNO/q8GupxEiabweOfKuZxI6eIrTe1xHUPxTLTQFygL458pbF4ER
eRU8wreKS4JVwdVemInz46v4faaXM2dSCqKWIxnKaS0g/FZKZOSIn2k8LvXeB7QDi0yYQgSkc6TU
+5fb8Her2TeizZOZUpVqg1otsNlbdLEqEtf430HoKCf3rwYbqAxPeCeS4Q6yvzj4bpsy1ovKJJF7
4ETcj3bBRnICC4CqZz7j7I36cyVQS3amgEzktFWf3AHziaj+y3BoEb9hj2pJcBy/fYKrrrwks5Be
HJTJ9QkKlJ4JHTi85gbPNpSxwxZFs/3pcgCldZ727Hhxu+NpyCwkQ8Kkzu85fnRAGu5lfL4LvrH3
VYXRu5HL1fnCohPC6tZm2sAyKfhFenaE7N4zSfVsAEJNg+Fvk27MzzoIROIj3cXce2MwU9TCtIrG
sjDAcn6cYRX/E+4++F9GhRmcT4qMw1/Yl+e2eJjOXWSEm8KOGUCcW7qSqpm+PPbfsedC4eGkUZPj
ekZRrk+d2WBplm6tf85MW88u9t/Rl5gf3I2YsyfBLi7dVEOSJaS8p0WP4U75LB6JobLyS4lwwDnk
JnmTNoKed33HCfVtqEOOtHTGoov9vT+Mo7iF0JRby3IdG1BLA4CUNsCfXc14z/wArpPsh8UHBH2h
/q1VfV565nr4Adka4Dfvv7zx2N0LhB1ep/vr171xxZTkKPUsblhilLJ0aO+e6P1oNlCYxWfuGPFF
wKUMceOJp/MskROtcbBq6bg+g+fmud9qQnmFMWIouG0Cacd6sRUXQArZLobC/oed/8lJ3m/hPznG
bSh0a0pOVckN5K5sQu0UUQDpNir98Juljnwfo3I2FmYsLDN5p4BaWJ4DAOmLjZu1QNTvF5oY2upR
QlF7LsJ9vzub51bGonRmDrYcSISrjf4cxX4SykeCktmELwuc+88BWDexh2DiwV2+GgGYjfUx2AuK
CTSSTaeTzV3KHQBGH6Cynn2p/RaX4Mk7MrxgzcpJPE6BVETbCQKn6w7VtMLZRbwxO+AAZ65EIsvr
z9RnWETmhSspOjU6bXnb2zPN0KrZTvnCzYpIGiG+ZZt3AE3+nnzOeVk2NSntOue6lO1Vbp3+cExY
XkgBrJL9GVdPvtqnfTsXJbt/oBhXVE8ERp9zrOMOp3131J0uq6FgQ+FccrL98DcAJyflGvFbpglI
33cNZ/GCKstdVSxmmFsUoIItp76Xv7yslgERJ4y5ZVcM+nq7Yoga1QiuNQL1ppEJeyoHJ6GLohJE
iq9omB7h23xgqh3BWTBfyeEQZMlgqaZWQP79mY6hsSWkGLoiCM1LBgGJVHaykKoX5kPMqgKEhrDe
Zdcg91dXW1/XsL++7YZLAmy/VC0KtQsof/TzukqKk3WOdyrQqF10hiXGmn0KvWj6dKCqiZ+AC6yJ
3DIx6ZSJhSD5frD2ophndDJuLNcN6B4dHu9CzDGoIvEuOme7zYjn+V6LvOMnQKEmFA9xcSiWjWVN
7ocB9m9gouIdawv/OruAZJDMSWLQhDd1TU2umjs61UjrMVBoTOmM+msT9u3/h3KXWtpBT/k48Vtx
Aavi35hHoOok0nof6zTZY675v1o307u3UOwzMFVQMCRAFVVQ1KLS1pB7rfu1FKl1b18aiGboIDTr
o3VZLvgnIlO/d15hFr9t2SnFn1r2dZNRFX29cZaKduAzLsio/wLvXBagaOoE5dmFVAQm7Zc1+4oM
BexwBBw2zeSfHDku3P76E+4fbLQ1d6UW6ixyYKclqQ/mIlRDaIwuwwbXyuAwkixV662RGCXeCWia
2/P0rxhWL7yQkB9RCQs7KfruRa6cvgJEg+cWFxaHnL4scK+KGOOzM3gKR5V6l+ngh7yBYRNgeGAQ
UuTJYL3nl5b1prsdhtMiM94uacrEf+E3J8bF1nEjHl/9NQV/VE3uTbmynx2Nk9/s23mL4x6eKwPP
XYwGKi9GSnE1ajhp9kVuYgFx5RitUyL2ktjBa1K4f4z7xuvw9KVDMLaw3Y0uhBTDMfFW6j5TXzXQ
1jDc7ZR8YgO0e903CrZUn/WIoYSN7EbmvyoaVeq25kjmjjoWAZRtOIBdzmyHzgyf2y4nrvVojckZ
Q0GPotEfclUZ6R5Tf1C47h9jtyQqSP7ZvBQsijZglfl/sVOnnA3uV1rrl/CQw1yUueGQ51ILEZcS
JcPwTVNE1+Y1gyDuL/b2PhwOgF2JQYH7RN3foS2rWC1vWueWfHT9iuMHE10qvLKAjf6UWk9yXuKU
KeeInbprAbA1T5yPDuVlYx0u+KLie34dOCfJs4dtZq1kRNbxUI+VrbY7AoW5frECQWlmIKzjd1Ym
x9Gx0mAK3kumzeIpxGDugfDAa5rMp0Mzn+t2Pq2OVTG3BtyCjZ4BxQKZdMFQ8bpZsFMbh5dT0lBk
uvoXJFOb0EJr0nIO1dlA57gT1NUrFjUaj8GRn5NExS3mLIpTubWub1xHUQR61ILOnkJqS1oc6nRW
MAZNwWrndL8kNYBB3+AbOF25zf6j9fanXu8p92LNFlhksr43FFQEHgqfOtS4Rx2qNw/t/kZ2stsy
enaQZVPUwslHzrUXJTaVfN+WU01dyyjCdkg6sTwdKZgqlIvX1+V//HSBWQY/q+uSYytORpg1B4uP
Rc+yLTNw9G0Gv8KA3jbtV77j/QBoFCEJlfmCfeseqssOMxMVfbq4MwBqpXyzRXoEHtgGGBuU3JTB
K8eza02nLslJedBjfvpLWZ6hH6X0TsC7Fn4JLrwm5XhhNxj3svyTOMPopM75yO97ShuTy5depA25
jVYmOA5MEQ3kEhwFq2Vv45KaTY5UDzQtGOsDu0m9htiETuDpXw9hbEDqu/s81Z3HQY9KjMj9Bfyf
sNQzyDW71jnDTgB1dW+dANkQi0P9NZyHj5dK2Me4uvokggXaAcEigrldXWgd7fx8XHkQSQlZ6Xj0
LsnKRtN2eIsU7805FdHBJgHYGeX5fLUetfBlHoUMoA9rJrRbjQ1IZOfhaEgB+0xEh3RppXPblqTL
TPb+nH0Fj2cRqCrfB8A6Ej/E31aeIrFxDEam/BUGmjTZ3ryDaUgC/WzXtIvr+bfGmzDLs3mQqP3A
jExh1nR7P2gklXs74UrCX+FLSsL41gpR6H/a6dBXXAuKAVYExpeOXaWd9I+FDabqX0Uzs7Vttqdg
2jAv5Tvez8GY7mo8ugnNbEHv7MSAmNqdvOJWjPBGA6SrbAO05VZb7Or0IP58rZPdKdLPgaQnopqH
4knSeQxWXsBA1JckfFrXneoUDAD4QR2wQTRsFryR2qM4e06d/0Cai9dSNr+vkXKpTTInJUBt6ZQ1
zyWYH1iQALdHarlp5t9LjMqiC9FToLT+1786lFy6R7wDcm5m4wlQaphchI4+DzBYxrhmzresg7Tf
0/kc0k+/FMrTuRi92DzvVvQlGC183VNTFc9iX/E6VeWuLsYsWkVUApbhBT5h9dEIyw/SjR7syHfu
2q/zYR0peSXuktSRbOiDzJmJCh0aF6np7LFRp2+uh7j6tCDTi0wX7NF0tBIWBtAconUMdCmUQsuQ
lF92rfo4Ie/BYl51E4Ed0kpT0wSv9VAfsix7Jon7Dq6epJDJ03v0n8HpaK9OehuofuZQ/HLj/opy
+q1ISYDTspNqNoEocD7seVbd59P/O3cJl5rfIl0124XU7bbdBYcSOfEbhPCoFzvk9aXaeZ+2j/af
UNFq/2MBTMfPfTh3dT4o0m2FjsYNi8f1zWCHXANyWltmnvcvqAiGU7eoFuflhEnlvWw2RWPQnEIJ
OsjK/oqYvcaFGC7tET2G6IfEIIyd1+HnF/KfI/d4UvMhjif9F+sj1wBuJBv8oBwRYt+GVD28e9uX
oeYFdf2rADaFCi/kHDrJw/JqtGAqdKdaE4RJW7gSf//pwtcIPIFNjtnbmm0z0IzjMCE2PqetMi5+
EF5TVRE2NkCpNZCjxuv3hc53Ul2xXXkpRf0Ydy8QrBpJBp5IF4/Eq/Rdh1LeO74amFwfqIfXBSWb
GIVVHgk+kAO2YxutIRfmBFG7qe3v62VuDCHzhRot4cR9nsRydk7U+FCnMHPAiYR/JJkG0iZXqazu
TxMrIrSTp9C5RKszOHCvxT/f4ZsEYcjV0I1wg1KkCjIi8x9q9qPU9pnygmXsxcCeyVsUm6dmOm7Z
BD0MhnGWuUszv8PIBMHXhmLkuaTxEmI50LkwGSdBwtPN7rJc5jEQWXKxa9L89K9lPDL/sczXkvHL
CM19nH5Hz92sz8ALOaKYKejl/2mRpkouDYyqCYUUmcxlYytLfRsuttxm/WtxDUfA9DBsp0KtGhgO
AXjjTMsxujR2F28B+GGpvrF2BeDvim8x/4rdZD3XDgcLnml7LCadmKnBxR0Hxaqdztk571mqQ0sz
FOqyBEA9z5I6p4Zchxj4taBt7M3dnOOPbrZCtv+bs6eSTRVHs+vKdGJDNkxjHCvjrASPa/iePX9p
i4uKaMr5HXlaIqOtyWBFrao9FVtgrcKq6vE38jginnZqlNW+vboeUTDGDprMqUcswpbT8RW7z8mZ
2FWjnuZoq6UL1rZh28u+7B1ZLcrIweBlwkbHpvYuAnTMEyUY4BrRdo/vIaMPcvt8OSutTCgB7HCO
ND2U3uxJtwlxWn4mLQ1JQ9YXe8aaLgrodGC5R1ExX7VVk2LkC1PaWIz+xRRq+TFv/TJZzWIG2GD+
bLPt/lKQSVQnpqDyiyNG2nBfBhq1bGni+bTOAbW9wQDzNugl7C5QwDO1ZYeiVSmjGczQUG+7vDFA
aj4SV/0VOPceVA49F+3yuR/JmzD/rHbbZ7M9D/b/MjKheVqpqpJ+PBRIpbMy3gaWUUaHHWO+UtYt
LzH4zVvSUVhYcKOJaudlsimP5Vspjqpxs+R2ceqv6wh3YMj68n87Fw4lTMpLqFD7L5/wIyh37/fw
sAMWPjrJ6ScMX9WyENZQwVGD/JtOVlvClAU2rSkFjdaVvKB87ZX67Z4gzst6o09Kzk03axiXwGkw
0Emsy3l0fp+qNy3Xw6NZYcjiWLmwRU/iW82L89Sfv086igxsJKsIvAw2lFoPSidrEaI/JpuQ9K0m
cxIpOZmtAp7y9HNPE7CdvkqV3Ihiv7Hp/UfMCXql5jO0r3gT2YSl62jkDpqsUmU+5UGYk5ppZJEY
vY8BXSh3Srid7KvX83Yt6iWcf3nNlcn+mpFNKq26pKntVy5rdk5S5Zj5NyyperSBNh7sN9NSRe3c
Y/HSxzIEHqiNLWqGIswp3RPOaMDNxB69cwdpXTNE78vGQ74AZil4sI2+zY43zYLAr51dq677JMI0
fgZ2IATzO4yIimM6IBbluBff7cVmMNRWWOcd/iKZRIeHxXvlY/3RlqIxiQ5xNYfe12hwsldXQU3z
fydu8BpvynWvTxi+qFsW2jLrO4rb+JMF2sziXgeMpAg3Lcbnj4cQwJXz96rhVCHhCaNINOjDiJi3
TsVkQqX4Q1spW71T4MMrKGdDWu5U1343X4sL706vXkCfri+c0ju17Hk2FCQIMKQReuUyvKX0v07R
kE6AB5Y9L3kVgWExIHegMJ22FpwQ3Wa9kM6HYP2MKB1XqhVMiEfPHW/7ckGzPK8p1Seu5cNmIVbA
yQkz9Vz4cGpVBnZAeb29KQLcz+OexNiJlj2Zxra+BPYSbTEQlWYqkgHItQlmZYjSHl5wMC/biUOj
zRhlft7L73nUinexzJML9KFbVDYeyC330wX6a3D35+QmxbgJXOBY+a0NTowUMGSQQNljxZ60Y3Kd
xepBY5OdrGMxxACl7IWiXt3Ezk8EH2LuO1YNOua8UItI+Q9b+nGXuJn3Cweyum7eTlj6gru6HelL
2DWk0o2or5NDt+AhL9KLzBPLQuivvSWxehP2vFiy0eGoTJVE2mB1UXP8kR+PMh+YLmjK9Znl+XsG
+6/ETdwvNUWvV0a9R64DBsqQPmayblO7t9mbdT7Q+dJVeRlDQJ9QCMIBZFHQaD9C3Mig//eGrjdy
nFdsUp6co7ubUOJ2BZivwo90JHgr43ZPKvTfTV94fuLE5UMHE+bYoqNjsfe5R9fWKf2lcnFo9rd8
wezOT8kjAp+OiQd/8Qp2Zuw/DoyzII7tMJ+MMixUzV2W6GYkpgtPXoP0BmcMPaYMqBXDr/GEKxg6
rN7A/gWjYaCXCvAw3blycIxhNexuTCJBRdtx8oj7AkLN7c4ERhGDrXeFTAO+YTIpFsA5jX8XzlZv
ZDAs8w/XSdCjlfKP6jEKJbFiC91RwOHTvUX/C4zQ5uXHb8CCvTZlf2HZ4u8iazFS8llMlRIdwtZ0
XLYwwjcD/TiYHHKzKlEmdwIxk5fw8Fx5dFs6f3Nf345y4GMAQah/WXSTT/Zfp6xawYG5I2o5XKVs
CTEm76ZZsc4xyb+eZzfrMUuGkuiymyY9ia2gfP4DyaFFVgbwBc7T5JJFiULLRTiUQXYayUDMZK3C
oMixyQEP4yr+sn3MW0/cupKyGnj+jYRm7JjodysCEbBmzPjfUcBj4xikcuulZO5QYbSWM5YUDxno
9QlyXw/xbZzpiaMo3F8kJbePVUKfImJAuL/dHLsDlPl8IZxLEPKrHVbWRdyfGRwFASxwcXCLrZCi
tCOGlEJaHhABXJj+Tdyxv43OqpkqKbyDE5Vg3NnQruEAJcuonSUmFqnIQOkyllQvgVh7tiKDJIFj
mTR8/CBfXUYez7QzAZ5/y+x9to0V5av/wVrxP/X5y/0h9YV3CLNO9Zz7d5Bqv4Tdw2hz0pAJRrIi
LN9GZ7PgQiJ3rxq7cc1rv9IFvuqVFKAi+5Kg/ulaKo1Va3RqrnJBQ3QbE4u2hDhbjXFwlmwI41LZ
whDAiM9fpOgSp4hpMk6erbgguaS3e3OAbNelf5E6F2h0nQr+FQnVoOv8Xfk9TOl//hsmZhOwkKEv
WVUphbjWFiCY19WUxi8UHlluSe4ADpnh1VTlw4SioaTYu9dgG1Q/Jamiwm0+qHgPao54K+NJ9u5p
hnkSJTpvDJsOtKmkoUQZVZID8nba8r6InF8L3xFX9bJ4Lcn2tQXfHKjTrH+e1imebGURALnPQ9pz
gH3BzhlQ/92S7r9H+lSdSI5ZiXjYhmN1XE1I+gEWWaLHh+CJLQlKIdQkjeBsXWvgU6qXgHp0l0Tw
Zt6AzOYVkWMFffBwZfLP4/+xZ20CTFsH8ECui0T3xGJ+E31ybOvl+9/je+CoRMXsAyMqN/A1URnz
l+A+mHq06OdZm4TT2wIoMrThFWFJwEKPNa2bjHN2Xf5m5wwIt//27V5mwlkfpZ3mS7uAxiSzxsa9
ENX3Vk/etapHED4lJ3/o+2COriS77HEUh4aryfsZtVLTB5Ia9S/fytO0ca8yfJ0wtU3C8f2W7jyl
U68SV8qQrAute/kDffo3gOVQDyFoffGvJQK2JNZGlU9/MlRRmfCv1d9gtnRnGQy/jL5/LaX8vNO4
MhEyIVf9GvgHQb5oAFSiCy5fOkp30LTkP3oSRaCqebuCtuHJ2sOP5jxqHz9PK6TpH4FytKDiXAxx
HmMARSStqno+xY2QDU82P4Hz3Gf4Q2nc5S4ZfeksCJTTvQp4UcOUNuYPvp7ppdYT3uC1F8YqHeCO
gO2LtbbY/cs8ZzpqzjGe81wF/kBJoJ1RRjwUW1AODugbZHdULa2kG1l1A+uJJKeWgPzja/P/V7HC
KmxHFJv2ekIf5ciYo2pxa0nJPCWDz2u3Nd5v2AsNzGR0nLHPrYpxCB79g0JKKdl7C7KKHYLsl8hb
xgV9uFrwJjeboBuuFMarHGGn75tRis6+9mD/8eIDox1asXh9ocPsLVi2LkY6vnh+YqELUqiKtqwS
j1UZZbuXJ8rbckJHZGY6Rm0K9MH1UUAGsm9LtzW2mxu74IgXAk7bwlNBkgBE+KsJ19cOBu9B6CK2
1/38UuTgaf25gwW3uI2T/p4Ta8EBTf9tZXiqnrAGvsojxo3278mJxA6FmimYFB1c2kRQMNr25+eY
GHjlrR9VOc6QFMBgKRTMc7f1Plw4AajTTJlA3kLhuTsjxvHxhvqDJqAl33PXmPASkzz5g8B/nF/e
AZ9zZbJdp6JmB63Jkn05GBQmVCs4KukVtFubTvwpVZY/crJcp/f69dlAwO44/6XZqtIo/dJ1kuGJ
gglGGgdQyDpeX0DxgapzbwQ8ZkDpLgO9lKZPX/fn/rGbSz5atNx4fSvAC4GzEhVIUH97sSAhpXVl
v9WSN3iEJwvaBV63QeXbR7lkEf1z1F5kcrGDGJ77MgFmnO31vcuyXDYTtyxt1eVzFeLSFqtO/F42
rRXk1fqlGmJLTex8tcfyAEBgEB5LnkHuJghqFUtJVEAJj3C3uxmPWNfDUSr9rJxAnuGn4YLSoVrc
4Gq888B6bCI8yttZMHeHdpavVkK4H7V+WQYG1Tw3xriXT8ZBaBqJSYZvm0MHf+6qb9xmFXnnASgS
eP0eNSQ4LlLRpe8g3iLC73vvQhmxPQcNMd7ZxcNlMT4YFL3F1rpITsEYUgtKVbxZbJvqrRG2bZRi
raeKCIQkfaKils+Tf34zjah1FDZWH9GhfWI89zQUVXM5v6FQk9Kmjs83J27Hei9v33yTmf+yc/c0
43FaiX2qnaq68W7L7h1M5GJGWSMZ/lDiznByPwHoD7q+/5pmm1EIREvTNhb5uyfz2//1jdDcw8Mt
qDaDDtEjEwdIGyn9WmPOyKrEt4ZxC2HE5HtxydhzNMT2dRoDsK/W3d1DrQNnLgrSmeJqBpij6PM1
GIIsodBwZ/FtrLwZEqLs54lH6Mlmf/6wGNOg09Q98lxHm1oRJ7FKylFC2KkBoNt+W0xd7MIBTHdt
E1Esk5xiRfAdQ3JCOBT7++sYBEunwp/yYc7HW2V+TeLqfH/+es1pAFSnUP41K1lxXAgiPCAnqfkj
XiloPdcnltxVazjAkv2WvDC4NVFnz4GUOdZVOz3zl1MzMJQfa/czkW32i+6zO1C8/GKXrbQ3yrad
j1XuWccOz4RXpbiPbV5dNKsZQwvIRqHnSPSbKwf9DguTKIsUz8xXX4oiCIR0zgpTYyIp6+P3pmr0
m3x1wlUMEyIEUAxYhiBeX3Scj63ADzrDrhtPAPx7BKdFIQGIaGD7M+9tw2gTXDxPvwxceL515Jx0
Cdrwr0aAvhR7aFyA/wngQD2bpRCiTJVWpchpEy4lggKXa31PmVmnX55LYMYlVCBVRFUQiXqzRMz+
rc1jaoNurak077+brbZK90jvL3b1iq/N4uJaVNZ9a1f58HSsbUI2TQwWesYEDYJLyFtif7pWwXff
1A95tU4xh5tXWKSRC0x22aIQwsN1O4bHcatj48BmQWcG0rmY4I8vjmOwp3m5CJIMHK8UBeW2Kh0Q
hy/iE7wneez26zaXly/KFTFXLDrRhQPNR8FeSAcMrZ9iBlVvgfbC+8/HYYmT2fm+8TfxFcMt+Jpx
f82qDN8WvizLjiwCGYHHn7V+SBABpHe+CFmqImzAhLmVyEK9wVkU8C3DkQ73pw4C8dUgNnJVM/hr
MvtjbyT+w5zzQThKDp0HKKKs73EABkTo/Vu2VjFHtlL5yn6AAf34yU1cZPUffzK4Chgf+d+dr14k
4PwMHaKhEIK71IkWTPuQH2/meBUUpeFNAAjBBL4UYUkJ8q2+3noCgxWLSQoC7+MId6k4tr415xY3
OvcnGB4H4zLkuxFR789VOh2uYkBb1bTLqWX+sCbAVjM+Xeds9adlutMKrYRI54SPicxg0M5bivNA
He5sIwH3QTI2gDD7mo2KWFWRWFu1uxgCBZ4fXmJVPITJvnXpTsgO6LJXl7qp7Vrf0PsPMYlkQD0t
hoFdO6lirGYav9jEU4N9eiGh0Fsc22KY4xDv9GFH8Lm7oFMKHyilSBpz7Bmx20kJoxIQRKW6ds/c
0OXBLDhyQmd3boLZ0sgjC/TEMqaBJHWf88v0KsJpNtd9lBKx0+mjdobQDZPPTDTUr7n0F2Itzrit
Nsuh/zouDq1Cqdbt1SaF5pSTJxpnnGHHsz008vn/kMRpQLNg83kUMTwKf1LOiNEEiwo3UWncL2Kc
tH2ZdyAgrs9t8VdxG0D1psS4BvPvdEkenJVFrDDow18RwsKy8jQKvU9849oOrjXjlD56kcs475LA
qoNFSH8z0O6RiAiWzfdl/fXAffAYG9YrwqFPWEuxH6N0VaZzVo81iLYMTdqfPyxNmJd476Ioxd5O
ituKvENA4zVrCR0x66XXg4OuLPa0juxHQyJNZLXLx1GanV4FW3vZJ61Mxm6VgtgO/7UEOFMoX6NY
fG+JtihDEGRL5fY2WFDsfFLrJIplPJ3sMxW1Ke/iHDsAL/ZjgRkyZvC3LEBVEHR8Kcltlflt9YSX
BLqcjctNfVRfHcxjMk44gRxuFRclThO7o4cNDet/6AZlHCD6gIa+GYHjIPwYl4ndpEDXuNjXxRDd
nSVmjtQ+vmlD8bViPvWT9T184bU9+l3Z4ZJLr3w4zkDpTI0dCHG08ZrPpUkMBVCy12MkEj/tFQ6V
8CN4YKqeg3EOpw2xm3w4pSWUT/nA6x1QzRfpiqNOY8GBM36n4LvPGFTAeywV26KKTGnJggLj9SSk
B4JVaOrclZU6WZkg261xyj5jqq/YDtriD0vzW5icG5W+ikdg2kLRBPEAehKHA9uhDr5s+i8+icuG
zM4ltF0VxOR5DLwq/trp0u27IbZRgmJVRGzSamPvn91rvzLv8JtNDh/D7Kip0Y5+1p3kLZgirK6I
NsqSu6UHPSU6D6DCSwvTQGnRBeFboUkjj58ebhxtUdckOtNyXC6v17zKN4N5ob8aE7fIb7h7XebE
7uzn8X72gG/r82W32gCYoskm1gd3m14sODPHtBqXDvxo4Yfr18mtZbcn6JTu8Do7d/RMebsD8y+O
1BcE25Rr2r3hulInI4SHZ0hCwia4uTnjFVT/cGMtGIY5CFG9TSkmIXpB6DvcPKboJ89X5jDHOQwv
QT6WEXukOVi9qMF/JCYrJAiJdf9swpK3Gpdt8WcmSjB0HIA+ZqsXypAXDXEoifWtvtu5ux0jsLn4
M7aOu0RP6EodK0z4bEx0elFQADvkntFcO8Cah5G/c3U8Hj/TUidWKvM0zUAxeLLtNUOxbslMuX1K
kymGJqifyWNCwqe6qpF0WTchyRuV2CnIWna80BSMZkXCSAu6rQZ8Y/lk6ydTALknFZyLaeLpikZi
Qm7q2Egtqey3dOj+c37J9e7jVlQYHR1CIn9pH9qX/ELrGh8wjGqSkVI2QmAvDbDYJUbNVHjPwjEA
MZISlzNF/Uebl1y0pYSwQcetyjuse676n2u6Y6jwiQ3Eab7645zvZKeFSYprR11eyPbSv1x9yRA+
a1D8uoXRoj2W3ezuxTgF2UXh7eFApDmsK1g6/dDOLeuxp2+RzOOeL4EqD2H/ZN+4BiMrr9J3epGP
uSxR3AlT6iNd9tqHZnjblD7t8XExZanu0lnQkiaC9kVT+bDaDVxHdEqLdgU8yWo9j1s8qsiTeX4Y
B4d5zO8IlYuuN5Q2DzoKbdCp2mysEnZvF5gwgh3qJMtsJIWEj7DcfgWKt8CM6sWmDQym/D8nk47X
M4dAZ99UC+GveVT/CbuXDKv0c9dpvCAWgi+mKbU2zN8xPZW4/AtlzOVMlzwY6rNYRX0bX7k/XtJZ
SeW/VuWg54UcCHDAIqWMLmNRVRita19jywF265s4dnCG89sose43Wsiwq25ADMjaMLa/ypMkkKgU
PckVQs9JvxmDKWii4DoiD4BK9s1kI9RsDNZanHnhWixfsXD2gEyKGJDINPFIqLKQOsHOdYaDaJhV
zcNflDAMJ4LZ5f4aGPLORqXnr6I0UczZG08x6B9myNmWn+nJlS9yFkjW6/18dPaCzSrUV4M4ltyb
OJzhJ50qCFzhfs+WhrhchM98cJ88wQJD+MPYKg+DPmr43uWCoLeJJ/9XpQt9w4iK8oACnh4DdMnT
sVOWdaFjw0sbhAhFziBYWLR/P6idJHW4pyPArPDmwmoEnctD7Y30SwLnHqnkMtJW9CFJTVUOuKyb
s0pKCBSvHlAsBy12kq6q4YLuH8udLl5nT2Wy23k3PFxwFpMRdjs1k+3TgN2jX/o5eZAnyoWxGMIM
QllXSUKIVQu3krvwmC7UL5S3L4yABrw6+sYaYQkOyClPM/IeZAbbBxSw1pQpOGJwdbD9SGvbIHU+
gn6Kd2JLtAnYRo7nVgEwwOiSh0U5i6zPYOrcCkrbc6Ej9dvgKfaqzP0qB80hGfraLXZRnKCLLPiV
d3EsY7VZpeiZRltt3RR7aaQbnfscK1ocjhU+3LuaMBlGIfu9KboyBALikQ1mT669yaMVHiSv+PHq
DbCpjFilO72THEkgZT6LR6pa6SXIh9Sb108hocdDabHJTcmKDAxw6tNKpCEuYa5Or5pHDl3BIgw8
MrVP+L24JR/8CIK3wI6EVNHp2ODcLX3MUYw8ENlNy83zjJlo+erADhvbr3DRTMJtOnJI4bYPRyV2
5aJH7zCpjqC/T+osVLmbP0xK1kogxxNVfIUbWveftL+vo5Iw20EbD1nWyNWCoUEAlntFbq17Hlw+
WKhbto+2FEHX7aXj0Y2ZtOaf4LfFxuiQ6946XY3hganXItnITlaSIQ0CbnBJthL4aPiI4grUzu2Q
rvrjGutFHYUjehrkF1esbkeZ6ZU1JcHWpF8FHDbEGlzZXn+OvSfzTK9SbJGn3IYQJV7YS+qY5sZH
U9JDjRaav3J6DJRdu+Izqxc8uYz/2lDk2LCmkeqlxtI0goyAVNeNutv9qsWS+/kDWhriKHc2YZAO
7BSGlMKwwFDsORpBW1Y9vm+NmM9ms1HfTLLNfd92NqWhQsc1maEI94vWxBBNpkL5fapyBJn6RFw2
HVfKWpyEgmDi1hiBxEgXh1/0Wh18ZMDmZridLXUol/qtyedj+3YYMqsjFuYokvDu+Z4viSP7Gprp
yNvAVAApMSf/J9TV+/0OgvR8lrYzBmhDplr3b+O/ne6v5VdOQgHFOSQaTW7pY/3Jir2IsloG7rUY
5eqg09ioPjipwWve6BN4WROwhD6rkqXFk9gVwFH5WOZPHSkxutjL9dIV7WztGykDaJdHxlWYkP4C
DzsQkA6tziVSTs5Z+xrtG3mXndAfQRjLCAxVXBZSXkn7r6hT1yJViTVwrhe106D5YE1FmYq2ZOIu
daNoJ2WhiHneCGoXkxu1i4E/+EzdA3ioGNUxesx7Zf/RT73+kqCVF27cs1qa2qpIBAGwduYQ1snu
k6jrP5vcl29cJov181usKH2cP8RYp9wM+DR6UwvX59S0UfYE0/t7qBt6CTQfiN7FZmrcSFmYUOif
buYrUz00sQw6Ka90/UsVmaredhpCTnhve0MkNJNnpN9l9TPL/+gKPDKgie3AaQyMpTxTEcWwYQtH
hasW5mhkofuutttOPcjIqGBN20ot+sKTGpf6BuqOnYECwsgTe3BjxmncaApUWEQV2395sZsUnEBh
3nBeohfpbIlZ4U9pIQwBk/vi3PemWWxyUhXbKDLB+XfyQRhqFXacFOGk7gZeP7dIj+ooQAUZlWGs
O6+cECFgu22GZDBzgvec0+5v08YYqOeKL4pHmC5++JtP+BXSg0SfV9ArVRTXMd96j1p2EqOfbgbJ
mFtsZVcZxEtvwpRsBVBYXWbx3/SrytXGOPPqIFCP3NOorCP04Vq7FluX6j6tafO9wumVVRINLcoI
N1ciEIvv1/Tyxr4lcC46OVDJilsol+WVj84aLjPndhKAjzVwQ8b8u7SOMJC+9Tl8JuFOK5pk2SgM
Iz60MBfuHZK/6NlpdSngrtSNyYHb6qMhMEfglPfH6P2RxekgRNPiMnf6+4SHHeBSl4iQtZqDOwxS
bW6e278Bxx8d0uhDJGwAxzkbQ3w1fASLT9EjJEyfYvxImNbmjo4JM7rbxBeYHvAQfhJQnX7NtTdu
pu2QV9rt6EMiGQco57x3sPSd4bsWj6aV5L10+dRJOtgp27RSqU65MqowETadn3gecyV5K/yIjN0f
U5D/ro2sEYTZpSxOGZrgQr63Xd5zprBW9wDvZ9mMgbMU6m8ITjsJ14RHHEJrdLZggOo9ed+DUnF2
MWHj2BMiou6Wfo/EG6NaO5mfOGWZ5xS/G0VW3LjCkzMLwMQRxN58CPgD6ehsDw0FwDwVSCbW00qy
nZrzShERGv1GooXcH3Wsn1bnxaAPAVqTDiKBF0GA/kjkpKUAgrzcsbDvKcHt9Wnd1rbViqe/sqYV
VLgIlnpbw5sFgzUhRnpH+U3a9+ZplkjiPElhF54Rxcsumer4ARbyJJC8Hmjx1VjaOlJPBZlsziPU
pQ77ga4EoA9eQ2zAtZVlG82+OB2WT3GTIuX1s/VLX3HH+46bxZVUwLX1xbSFkOmPImAoxE0LebpG
1qwKPvoehDKpmYOgksoWoZoRHqFmE452lOjA+KRqdd7uwkepKaShgM3GEL1ijSp0S37nQ/uzhXTw
42imMJzYcxLXa8g/shkNn/oqjxR8bVZQ82qgyG3XVEh8XBhDBTO5IvVBp0WC972qgUiILFh7aizm
1CVvmbTIqoJmPxTxnFm+wT5vSS4gHai0fMr6EvnOI9W0962KiYgdqABl6CbBzka9IQMlZ0mEkGtw
tQ6Sly74Q94w6tQmlHHm8JDsZJpjrDgQimT+AQ4gQVAGjfk29Ovy+vYmbEtxLcb5p6agHilnn+B9
Z0X6IMJQf00gVkLBd3PSBUJIGzfjOvYnv+xJTavx6YF3NWkkqsM2QqxwHRdq9xTquWuL6/n9qPoE
K5Jy/EIX6fUC8KHefpAq1NNGoAfzkcOtWbwglFEAIXxxwfU8IRoXxs6CJA5A9oAUfqm21xBayxK8
ihh3AO6NKVb4t3Cg5dH14C7bNfG8njUGPKDKcKbfpTNZELFVQWVdlhVPVQRlWeenzosBqH0Ka1+0
2QSw2WmK23NGq6SxPtrWDE6c0OqyuaY2OaHUHJrDjgnkMxeDcPN89M4cK/+lDfSqq5WbvNa6kwAb
SW+50Ns+HBzrk9hx9C5KsbHV/JOYqJGd8VCYohYKBgA6hp9ooWhbntuSaiB9eWw9LcBSlF0A9x8J
aq94f7X499O8DJ9aqz6txXcm2weNgUxlM5T5kih+rV6Iy1E8sQMt7DxEjwVnrIzF3SmIh+cgTgog
IvORrCcye8UYs8Bj37t+NGm+LuBNDA1HwuWjLZOvJXCxgEuRsy76HZaPlple6Rtq2hMChcdXIjsS
XZZF8o5BD1N/7C1LHPmlw8uo3ZvdTnHNXCL2Z7G6nd85i3sCA3IghbC7EQIAuCf7bk/I9ksSvYaW
2T8JMPDja8HdWj7KIQdSSVkB4Mi/fu4hGLcyBEpyqyScTA00PXjOedbjsE8S9UmXh3H3JZYsR13j
XnYvYAC6LFXJTp7qul2W1FqbKDWglTwOTQVrjdBHFYpUP+Mg8nQEgfVenXDfm1KMeD4ySqVbn0d+
95CGu32DqHezwkMeNSHQSn9eKbPIMfyIhktc386tuLGllBXeGBi1W0C5aJE4YUYphGSLIH/fCkuf
Uz9X/hPyuGeALHFxy2na2Tpp8fglRjocefyu5THSxJfpGUlFVJKVtcp200uLyhrRe1ufk56V+cEP
5uTrufFturNFRvHu426z1GZjb3hsz/lQz3mHk49JFashI276yKOQJ/KfuN1GY8F9NBHFCdLvV3Ns
GuFmz7hQdRDMCW5t/t1LkZU9v2nHKg4IhBVROEur+kguog/zK6ES0j1YhS3CxttA0UuENmT+/NeK
Sfd6qmW9fYyVRWWvnC4lf/dIFRSGV7iQJPRBnfyebJ1iKSdDfigTYVrwQktryL79Q0chHmqFuPGV
PWsWUVlW+/rye1kdXVhTLMS5hIAdRgQghjThPeummcIil68C0iwiVoZu27xFbdnTojNbYQwaqjF0
rW8/KK4/XhpNGlV6NxJMQS5LP6UiY6ageFpHOA/LVCoXX3zCqJFEXxNMFDGugudpkE8jQEuUR7r5
DvwTCvUhDv9rTzmdbJXMjTqRmH57YuIAUop+oJj8KQOuPYehq787RMCK1OQ7ch1DedoayZ0/bt0n
TQdRWsKIPbmUFzf4lbjuWBvbWtgwT7UTapVEWIa7ngWjRBHrRbjsKdqEXgk9qOGJEyJhDkl4KoMk
r94r9rJJ3rTz5Y0xt/rdoev6MLavKy4liJv9CzPPZxPBZdk403lSlargGOkLxmBSpli2VyhNPuUI
pqM3J+vL/nabzbGHtoWUsoaDqHDUh7Ik5ccC+k5juo7r6DMwC/ZmfT/yxpZbjYvkfqtvuP0cST7W
VRDA6yYRAR4CN28Vo6T8+WBTY/GCJYrNnTGbwAB0X2/tSLpWwCRHkpOxbQlZIHngwSkBuaY0j2og
AUNoGDupi9ShI1beO7EGROxFCvqEtPRy6RRDD4mdJ18k9RCT+w0N2IogcrQnUSKWcbwU7uJen65X
I3CswEkDAyWK5iBl5hohrB2cfWegs/LuIxqMMJ7PcFfTM3H3rKYa6N9Fsrsq1qb/ogdIwDcvUMKa
xZWez1BBWQBWv09oHBSyFGdzV4/yQRu60EpRQ5njr91/IWQIJW5jt5qWnuT1VROiind8Hcgvr4Mf
0qfydH0oyPA0ta1VAdoQk4gbP969Gkp+0uAWo9C5Txfk1hc40zE599xlwa2D/5VPz1Vkg+Vvk3FT
PpwFvMZ6ocATOaH9kGV9ZsZ9NPa4xWCvsE+cOBk6FhGdtJPHaaPmCQQjRYL9NBShg6wk8+xVz40x
bFpjwwmVgHqWcwtcvCcLADU72iM5A2MlkphmhygRvkNyeDzFWOINUiwS4LIFvblxSScgPZhVRCyz
7uOUzZja/4CNIvSYaGpeZalGoTt/ZcNbYK83KRuGqhfy42/AJbnwmC+lQ/vkLBeliSFukdITeWnf
cz+dyycke4Oet2QslXQkCG0CdrLpmcK0M9nPmOBSKuB7WiPF2PpRK35reRrWeP7bN4mZgrlOWQxE
P+sCL0KR8pqJWmiRrTaRFyPE5kDkcL38Y07ojFXrPo3/uIn3TTMw9r7XyDmPH3tIctjyNufAiCa0
jA0abeSyPnerlBy/BlqYByoaU/tq/z7Ne1o5Fbdy1AfhMr6AB+fDHcW5Mqj28KzSHFUC6JPfjipv
D79t2JXo4T6z3XaEXsTPBe/5IYxYEYg1E4/iAOqMI63V+AiI/JfyoPkcjuj1db6e1FPvnMV008NX
bcg3p9N3yFMPEJQfyXo8EREH8gAgEexuB701JUoN9729luqeTk8JhoS0v4bbYYlMFREJTI1HBkT4
TX4j1A2//GVkZvpkVtCi3brMKkOJ/MJwEi9zj2SvMpYoCf8UnQ3BnCh3aKxa+Pm9I0EiLLWbJ20k
1Y01D2MZ/EAaq2hr1t90Glkf8dnm/ePEAqzzRLr3q84jW1TIjmyacp+L8jVqhCwJitxw5SK9ZQHE
xnQRtcyHwqAeFxrbwIevM68Rpmy5bnukjVnJjhQsdLiC7BbFDI230Ha7ndV8/LwbhImdzENDdv0L
89lxIcsfMmHVOZeshPbKalJsY/T1Zt74KR0CymYfTrPitJ9s65fh292D3CAAeu8kugiLYsIFNJxn
h/El8mx9FfAnrE4wGnIPQyGmI1uAp+ROzamFp3/wriJpc7KLzaQUD4POvlrbt4EQxayO/eh5ENm/
qTB9z9bUAnhUBt37HpJcVB0ZpCydufNiNl5E7O/QmjNoR/oAfa1mWNlzGqz0y5bHrROlUj69EsGX
vfr3QH8Bn1obFQ98jqNfoBZYHFrlTlNtNVnx/GnLgXfJE/aPUIhOSObwct10wPr0uZW5UULe/R82
X4lPZrQ8HHm1STPKZQwcyXtezDqN6/1mT33xDaB/LLd/ugQcOfeVF9cGhO9ldUJEPsEnFv5PfZML
vK9XkkIB7O+iF0uhBAAW07YW7rX+tUB2JgC3vmoyjHEq2bUsgR92LMkx6ILUjnvn3HwA56NO1HMO
hi7CckE5TEO1CDv0LpEiPDf2SMcoi2h99yNd5rxZM7UM4cZ3IIphUhVs1Y8XQi9jSNGZxrm5SRAg
Nx6CqEukTOpAaDDHeTsJ9/M21w2Sq3kf/HHTUshQQNTzTFCt2zdsDonjHwozthTrW7gSM+wFNlvr
PAJzPFWCj1we7icQIZ7G5LpUmnYN/gkqtfcO2IJTXm/vKnRVENPGqUWCwaKKad6mZbQXFUSgbfaG
oIXb6ZIk7scc2BdDJYUaKfogoq1WKS+xM+5UucIRFAKOxdF33qZ4SVEsGE7OZVocqgMGJe5Utp1z
svszw6I+XMU7iQiFTCRLJN+2i6yEBizDM+coGQ3KLcZIc82DvPDbzJzC2H8aKodhlERgvD1yxayS
o3NhPEKK4igUdnd5/g2ZKBXb3l2FC4Ute6FQb+jazwXChOptwqLKm4HYLWzxI3VE/R87K3oMhvRo
pYzLVIUlRSfdI0zNvdPwMalk19BW4SbTvsgP3fhySiIH/lIN1+5mxKwhRLap3X89tHv09f5ynaU7
Wc3GNFwvIZbFMMtx++LYApTseyoAa+K7x2d6Jg7afcahQZ6bbl1zip+2sxBzUKQMJhzkc8UtS5eL
F2AVumxJKXK5DLChHgkidoYt7XpjiF4ir90KXvSaNQsVDPexW+5Hvy+t8SRkalD8pcbKavIgFi4p
jULRnu4U6frtumJ5K9lTWxzxPJ7E9DtqvSiTHxMj3DLwnM8Xp0dvOz0wBtTD7IeQYfrnUMizfZZX
Vnt+dwkkrja00YxyvRRN3s9CwmNLocAiVunYOdsjAgzI+UxcAh3097uanVLV/DUzAcUw4hP0qvMh
nxtOGWqaWeBPIWce2/+DNHjAVRT87okknPgWjezv8PBjIUzkE+Z5JqGzEcW1wY/DZZvrHPU4knE6
tY5zzUQ4j9XB6Yt+n1M/LVB8BphdaV6bZuVqmZZzsDUeXKB/KgFzCWxlsbn/F7CoVlDq159ZuDOQ
RCoEQq/mxZiDW9GVSIjF1EALCMFKvAQS2pN62954QJ8czioGxq/wWJX5LxON3+TUCDq6/e06JcYw
sCH25gP1oijppqH5mXNYcC9nEPMDhTjkQFNPnLEiEG85VL7lffFnw/ZcY029MCeXnz42t/FyNtBS
Bckfo4r4aD2nKLdxrsto0ODDgeBO5O0RBOtRc39d7nkR59FRNGyllfFrHSi23/ZxzA6LDKYoGONZ
443rQ5zTY07Aof2sFebm1jc0EPmr1mv8przBX+sdtPV8oTJz5BGvuee3n6Jf9yx0mOqW1gt1iH8E
6+f8+nItVa57pQcWX/4RSm5RR9C8nT7wGJEe7L8MMF7m4adZ4z0UsLzu239kyeg57lP+3TiNgeSL
SFBw+18q7qGJf6kIUgNnV8vjRG5a6jkS4jQ9FSzozjT0JOjPIOUczPqbotWBkPZx8ihy6AxwuCof
1wgzNrUmJZP74w9G6UQYiAyg8fwZHpXo5AeFUm+Gc2hBTqqEhPo905GfO+Nm2LULR4TX2nkoi2Sm
Rbs14jLxoYkVgjgvTFOIVnKGbxmViDifIw+VwquASeD9LjgKc3OtFydEmYeYBb99JgStYayKbSkx
iAsBOoA0LA8pMOAadf97CyEdQ4xUbq/n1ly0YqRxaAeO1brWhkThJlw04eJ6ocnUAq0ACkXxVTaY
dc/Nt8ZYAv8Pfn0SNlhwA2RPALIcWNrbXTmNyp+9JOd6mFisOuQ0516dzJk+6JQLgFwue1k7CHO5
hlQY7izi02bSwV9D/KVaiOWhHzKfnuxA3OfdjfjHyh4KSjdcve1n+dsvuORrOCN4B22tLrh1rR+U
buMcjxIsZAeuvC6D11Y87xgdWrvRPPqSMcr2w6EPnlbD/o+MBjoKAwniV++2wMMp3OMwZZQIPTdh
BvK/RkjiyTKKlmzzS6oDWeZTYzgQ8GfNjY1vc48skqGyDctpG4Xxwz1Mo6cKbWS2Rf1FjABZ9GmG
PgXX8sbFMW0DkOuyw6hjO+E5snpIR2zzSq1DosV0VET9MiGhix9tJ7L7tKZzzdTM6iCd5turQ90v
ljFHchKsDR+gNMX2EuxSu9t1OgwJq5tHB2LCFj0zLT9wtJ0JopY7CykU1MLAf4+iMBmRwvzvXs2+
XQVuuv2rmKT7Qn87ug2vaVVQNnlUZ8z9nltkyX8Rj6BsZgiklkFGOJrW7mh57UONF2auwK2ZkDVq
JfoaHSqALSUgq+7ZI7SCCqJTpPwxhvvT/YgxlTswiyO3Ki6RaWetGIT9J+GQslqMvYaPDpJPYYVH
N1QePAlRSDZgZvlT/Rtl2Y5Sms1/ZrR7DnT7f9Pa8oZhvZAgp2za3eK7/6OpnX1oxlYqCaXDF8Tj
tWPkpd1u0QZUwTTZ8EUjT1OjJ683pHWtjDbHNavbcsYXuOngHgQspz+5czXXJeXN9HphD21tbiKz
UfxmnP+SDYBy2NlYM6tznZlpjdk1iS5cPH1/SsvlmrFztY8hNLg2PHsJ6dR3M6aA6th214zZ66a4
OeP4Me8dEVxbr+tFu2Zn5T5D/OQbbvvYH6dZTLL4nSam72tGVOEw57aRkfYDItW7RRALOOtPam/t
0/ihxOK3/JXyDObRKXoIk2dNb/re1Wh0IxUwrp6iu80pX+xTU99gEOf4woB7sk1bhQCGcV5plUlG
NBXUp4QwbJ21t5pohQkyZCmqGYkcPiPtlR9b8NXD9TmhyZ36NJ5uUYmIn8h4xKvAZ3x/zWq3Zu6t
k7gZ5pBLURHYuz+ym6Urm5nIZ/p5T458rMkpo/OG7FjSkrL+dH4gcYRhbQnG0NTDIh9/75M+orGm
JmiQd7lTUrFkIfKObsBRvgXUTRJnwuiDFcPLzZOMZ91HYnEEoqrLjQ/N79O29Tx1VD3Oy1snhqae
tqWmKNGb/c4g77aC3xDE0/qBYB5vehr77QlGgaIyIhWaP2n9JmvcCoYfI1NvT5Ac8QkG+CYO8C1i
nS0Fhiaa+Lekcz1pU6TBqVh1/jIOGkCeKbH/3GHEw0n/ptBcQm3fINAEeu8qaQoZaRqd2PGFeV6J
Sj/cycTXO4A3eS4eToJh/6ztIxcp1dVTXiLfowg7KGTC4I7d0CFv7nnjyA6wX781kwfyV3TTu+GL
WyJj/v+lXlcmojWNkEEhhuKypFOH/hWTU8FrCZnShwipNXw8bqt3Pw0TePfzgmCNc8NFf+UJ8Gbs
n57B5dujpDXas8R+pXucmPv8zk+FS4UZ3y9I8egfEYY5omtwlia0P3dPvce/FVMEdjUuyAjir+tJ
wr9QDsXd9RRkrJQE+w81QCVuY21hyyup6nhcNqgNU+Vn3TW/WyfyXsgMPN7jJgp8q8Ue9U4Wlzwk
aY4VTfLEWvHaowcjEd4p+17aziw7IPzC3vu/yKw9btRahoKSufKMiKRTnBO0HDVLX+hv9Z96nF7u
aPjapZne6Yvo0pwr04rTFg1bIpjmRT+uTnhAouJENG+hZNDnbRYqoE8GkySP3h3m1IJApmrXjckS
uvTb0y5ORSoGEf0INhwlF4l3k/+NTL8Bpft/gcUDWa+tJkuN2OvplBXrK2pswtJNhImtdxFfvxog
Jv18j8NuFfFJkYARPo9NeceMqPZsUW6TF+R+Y4MgYa/iQGFtmIKfDiAIme9jrFiYJHL7+rGKO/yp
SlUhiO+B1ZTRifhZKT1hYHUftnoZy1eB8Q/c3iMDGL3LDDQ8nkrTGlRFHARf18XgJd3OiLLZW2tl
Kn+mSvDjW5VTbwDUTMFQ3nQicVFHpifyrbIhbOs6Dc5W80byHuaWnVXrUay/i5rVSR54of9xsm2V
7/OmGdKrW6WajWxup8SOWQTVVuavZSs6P4ndrl7/tm1TlGmt9ZgI0ioGCMFae9NeHz8DGg2MBTTB
2Op5uuUjRBbnvyBit67vKU1VwDwqxobCLRQDoJCuqf+kLcD865ivoO3Oz8xNOJB/KixK1jS6tSK/
uEaaG2FOHZuTlanTmx2i3+OQWAUZtFGS5KrPOymHCCzRSJ0T4HRwhylcGAJrrNsv55upHg8E/DM2
ROvEYpUAi4D5ZhSq0Th6Mij+OXX8wEUCo2FF7fi+q+3+J8Y3+kaRbR+6REF3I6VVNJ/0oA1B3w99
9Fztf0InzK2HZ66wURM+Ge1YsoRucBVKArc6NE0FF2SkPB4zcb2L49rmljTeleLJqIXyo1Nb0saj
tyoUnA4ThWV8N4bX+Do/myou7hQPJwE3rmbPbRGf5Ce9TzgfmoPFyF6LK/Es3BJTuiz4LzwkAAx1
b4fDzCyaoNnTGSl3Dd72hbZ3WoTpgJKBjwWprjR9O6uLr+MUo7OmVYvt7mOWHnOvTn4QBJ287Ydv
YSmR9CXno31+5THG1ly40jgMOMRicGF9S6h2tkJShXwR+jiGghWN2VpCSAviyE7MKWaJno7pECHZ
V8E+xM8AODX7OWVWpwRRxHZyuyFvzdv2+A5LSOSNEJnxBqGkPv126gAf7kWNmo4GT1na19BMpmHq
+fb6Snp8nZV8KImoxmzFril2DmOCsJXng24qCLmEosmbzoMU4EubwddjjKS9xYr+kPb6h+mJQERs
TFJA0WcuOfz+kRtm01IZi8zeSkwlOSCgBD82X2HAcvm/Etfb5HnY0jXrBsbuLNuAq1NcE9SUrr04
fYa23efOUpESXppnBiuU+/JdQ0WWF5NP5Fho0e6v2JRxnOgAk8h+pJ878KJltDdQ/cYlkzaaG+Kb
nC4ZNs56we/hn4O6Yd+7WUhiz67xcAOhhf3Oe2trJZIB3JYq9f5xUHT4FZx31E5lXfzKSdxej8wP
y48geDf0G8WfI1I5zcQm2UaIWMzj80R/gYcb8WgTOUDuUyUg2dUIkwEpqvD7ORZp9Xci1xIbo4L0
u05k33aVy5A/qxiRrXqEqRlr865Jtzyj7KuFBL+IT2rHG6R3v/9Q0YYq9fRPHaD1fLg0Lwijt2nJ
4KnUn0OWk5SyapMdreWj6cGatNnQioiol48WSIITAKhCo9SWBk4vFd6+J7qKPauDSQqp73chjA6f
NMNDagAVwkdxr+9vBcoEj72Ky1dFz1sC1gWJyq+Mo9jrWNjxqDjsekOFmRt3nQdlxaHBQX6KQCkD
lGBi3K/fd3E+CtCbmzO0QcvQLKbLllFavKWQLgZI7gMFELGAjgx6jqa6RJv52ycJGdHp6YGZuVWW
O/k2vWk1G8t0pn8YvTVcPve5XiloznYSzj4ny2e1095/dciLqzM/GIc3Htrf7RevyyChTuup0JdG
+7ldfcBT3TbtLetZWWylCPI9p+7HF8AdBaVW355ZoBSIESbUvduensYrm7vNcJOVDAAJzPr8ItGq
XRwhJGr0OefWXdw4lmpfJhTyxa5Qi+Bx+md27P/oFsHQJpmfexlm+CqIj1slvqSXT+/e8UBSz2Sm
IP8VxdNmOadhBOpvNOC/qjMo0obcSsFSTu9zYtyr0sN4Nkxun1Q4vBzn3/1xrhpxYiv67FYVUHCD
8awkrVavsoexqj6JcCxSc0TL9AIB5odw22LksWUi9LuGqPhtE0/XzXjg/germb132UkTlmBex6hA
nj7S3OkhYd10QWSKEdzyNF2UeNbG4SJHHRCoJETvFivsB91S3c227eLNooG0FiZMvwif28dNU/KA
Y1+qbmHbYRqgf8xI3KAB1NTdPNYGFk9Bhci7Rk+Bywwc0dRPCxrgBJ4zgNvMFIeKe509W1m4PFME
Ummz2Z5l9SWelS8GjZUwRZBYXMpFW5GDXh7q1rGTxCf6O0JpRrpvHRCbfKHNA21fGHGk+sjpDbhC
AceZcCuPuiujbS/HLFWuEvcaJ8YGbPwoKRfciIdvuo8garxK2ufYmGP2uB7ggrxpTkJT4NcDJDp4
TgZtOJoJAr+yW6+pb6Ix2z5Sk9EG2t5JPrOYfXXBMlI4HtBTW+uMjD084JDKw0qASHM48E5DSAD8
OlT+0fJ/XShF+PcpKExixxQ2TkaU9m8VTKax2VwqsVKou4UY3/kLkwzHZtKjj0yEhuAtaZvKPiEw
RWtv1xkkUNGBJsoc2oJ6zSW+LOOSntqWmMiCbUwDmNKjtOi5U/VovUXmoz4CkF3tdS1Q9vZ76zwl
nMvFwNqElSM/90iuqWN7ZzfOsJmVH44XHTuQykxDFMYoU0BqNyyqP+3gWCQCeN/Zg1piFMqF9lgT
giL7Dyk2hPX0tHnIJ1uMFLjTApbjo8Al1GCbqBHOu2wY13If3tY3SGGIsNkGOryHcqvhevNZSPgP
ajJJUUGnw3bpDtHllT4oRt7Kg+yI2fRYzjw1XEfWwdACbj37INuC7M5J5rPcAB75XCtZYGh1+rgb
QsMFChMxe2g03Il6LdLn4nsmY4GRSzY/wVbb/2QKjM0JB5OH7KrrqYdDywcjiA20j+p/0auvqV1k
iI4TVF5C5sXxyvY9Tsoc/p6f+kOiGazXqRg0LdKR7al3BPCCnm6pvNF5sxwD4jX52CtHotGUmeEG
sT6CWLYzrF2siQ3Iq7qi545end2OV3jRY4pikdfwZhYIlpOydLC5s0a+eTAdaKIgFb2qAqPzaUTD
MMfH5sPFxWx//DhsAzTqyv/saxwofDWKod4YIDW0x2QHRomsM9K3Cq/iTjpPb1wB0N6k7Oz0b5Dz
6l/w7z8mZBRI0J9+gsm2izkN+eK8jkoDA59a6gEnfI1uBDDL+YDnd27xGvbvN9CjKesecrPwRF/F
ZrRZTr33WuCw1kFDdfKdmmpqU5CPAVriIdSsrurw6/h7Kr5XY3dERBLaMTeZG8DN+BDn3wgHEfxp
diNbFUDvb6zwml6Lq7Ur0pKMXPJVm9y9eMl0lrK668gaHpjCx/qRM2g0kSiJFiwRM7JvLjI+17AO
Ji0nKZMJbvUeXceMCnGflFJWX719EjcL4rKL3wF1K/HdnrU48Ixeh5UX9TDI77ECaJWivRWhvlzz
kWkcGvwQNYSovB0qrWWkm9Mr+7pKnV8yaZp/UDThqtcUeh6wTYTfFN2fBc5XKHU+dIHUy9sD8a+h
qmw7G3V1SJKZuHf7RfbXF48LTppWShnOl40wik1bntnCPByet6Zk5wCDQoopr69EZPpKrlAD2WhB
S92ZYRYlZXN7fgaNvfWY90nkCBlwmBldtPejLg1hQdMibDv4opeUpHBPZfFePyvLJPh6nd8lARrJ
09INLdWQAawdbA9EfLh/Jed0X7OKo85KGpS7t9aake+lcB46iUYOVBZ2swstadbXTFBEmAHkqBRF
5e8UpRWNLlplgsGJsBPGukmS3ilzDsyOphzIo24MwyZtvclm+hbSm+2oO9m7N9/b88jIHIbdL7yT
ezfXLNRH2qZsePlbYQG894NzugXcE98XzXPpvlmWf0HyIBKKHNse2/lDPYEYNGxJhLK9Vv6Q7L8w
cGHe+k7uurf42Hvcy24pwGXSOZqbiiUeROVcm5aRlovuHCubiZxpmCtHuECu3A/x4KhgRygJGvQ5
T0y9w1JWHQkLHgk7JOu2L9HV5BKDhj7eomRjqZqHxSGkuBKMrEPveC44ohbTW1MXBcf9aEa5pLpb
DRedZuHHvrS6kGTBBmO6v5695E9y4zBpWMQCsUSgp9FUQECEzfuu1bfXILlo9AWgB2xrQ+3Owa6d
q81ktVcu8gnvr70CYJrU7KHIOAWTGVoMmMjEbuypI27Jn2HJnj0G+g3YYgxrxLiwhr9AZBJ5oZuT
DJBpbXuGwt/6l0aFA3DE8X0drI9a9HXOER5NReVq4Z9eIVLmdt7V2eiq/cGzdhQIiHgBDGyJAvYB
4DUtp90oNk5FxT2qkmbhT4hwq4uxHL7SiXNg1KicNKJMpQnYIw6JBdze6AbkETL00tsKipTIC2Ob
lscwhyz2+l8EP11eFo2LIBzF0qLHQwUa0HuUd/L+f5TWmsUQT1wIFLfpPpUlezgUuLxp5GUaE7np
hniCRIj0ep/6qZHLS/m9a/D13hvtxJt1HiKy9my/3pIsFcw+MPhLGsFakNzEcssKi0Lcp/X72dkl
bpLHVINFbpgvpNdIAjn3prbuUpTIyMkrkKdCMXmS+pBshsDGFSuMLZaeY5SIXfPs3Ovic8C70vkF
5/LBjz+2TYoH89yz4liGfxVZXDBLmBihaj6Uko5xJURuGCMvMnKW/Z9qHeopX3My0xwT79vvTahd
oDXNEE+Ugy+4z31j1Rou9kvvH/oZRIcX+0EcFgRrU9euOAamvJfEi4LSL92VRWUkfy1ii3658K1Y
aGuzfLsgPHyKetHqJeVeP6dw9P1VtTL8DzgC4fQrFH5PrzNTkAZ1qUmGtoOEvszLiJ1WOvNy/0YI
BF3278XBt840HrU3TalwcT6RqBb9Jn2pwGxxDyUcyD68P2X5agCUlPr10dnIGdRH1DP7LPp9G0fa
/tt5RoDpABc+6uawbTyeqHqX7G1BjFhWZW3Ohgr28IyE1pFlnFFZKC6wdCJ87Jk7OCsd3ob/k5wn
LxyR3U9EIp+Zn3EPw11vwumBabRCDqgGcOyFKt5GhqYYlSm5mAIL/w+zsBbe9+91v9IHNHlhnIP/
XubAsgwEoqGbpWUJSVtVO6keu4r3Buf/kzgX1jMf+SGOeTgYXSZ3DnnfI1ia+SHXRavlT5vr7n8k
SZgkFrMdPqaI8kh9YV2m3fbAWElajm+DS8Zlv5sWu4esvupGX+/b94Cm4lB7x97lCuUc5RuIPF3u
frK8jZbqDw8sHtxC1m4NIFem+orx0IdBQj10mNgynu/xOU6keHCijE3mmeBnTJ88CN6joEqKAvS5
vOQTLSUzW7A2cRIkTp0QyXC1dhUrxoHI6+zAoCDuozOBBX3Fkac9JjKpCWRLdVrScWdazZYYJNkC
hSrVwtXTCGXIW5UwNcTMFMAxblz6YRYrWOccHGQ3Jftr70gtqeh0NDza50/oJm0GqeTygKJDpDha
SXTnpltdke16G1pSHGu0qXsTFaN+xPiWNetHJCRAN9mq/nRYg+ouVF7wIDcFGoX2QXhO8V8TT5Af
as2UUk6Zt3ym4hAO6NwCkp55s2+MNLdu3/kr2+RvmN4vOwrZKrRzV05lfihnQSe3alhUnFDq8Bk5
RSVvp1+Mew9aonVQ1pNSQK/oVPAjC05frW0eJSSqWMIzSSKCBu+66k2bsgeNJR08rhiE42kjk7YV
2b6AXxEGeLM3B+O79X0IfzyWAbwLUsbypYjLTHOms0zzN0Sy3PhT7DP/Od/sUF2KXzEevpSjtb2m
BIlzWvk70+7LvOwevqos6YmENhKQuGr7nhqoNjmM6wvZcFL/lMo2h8wR0BmCE/2KnfoCa/ZvbdQK
1A4csepZH+RckR22z1Yas9tXfVVhjuwHGngA7SmCN3VaftH38hTjBLS8z0cB6UHci12/e/1d1oHg
a/jfUJhZ4FmWLNMqCh7D8GWjqTP5tdvP+Wuo4EouFCF3l04bTYwCC6LVbjkxKvLY+ktYAbDIUsBY
Ajk/4SFE1gyEB9XAWwTSV0M5lRUzU+O3UGy3KK6w3fUabX21u3qjlqQP1syUrZW9xa+Opd6csKxW
TPymE35PCV/1L6e65OWByLxj8QcP6YihBo906+DtRWp6se35IOtgEeSBiF3X6fKR8zwEmd2RjAvI
qQvc5MX+5iFx9gjlUr8Jc4y+mOesX/jBS08tj9D26DV2SelNmR8se/GzuJRtgz15KhKM4HHzb2fc
TdHTAPkNkVgeifrlndjA6NOjMzyv6xFAVjgN/Bo1WJIlHCUSvYVj0WvYbnuy10l4C0qbZzlVgWNk
kTYQELGhUZGUN+lFjGrSzDLTaYTUK4IgZI7UfrxfQVLrIYvEuzE+6kc6Q2y3l4FRCGBGlguZS1eS
fym1PDH51rmJ7EomYfum/gCYsc0rylFtxh6r0/Su2qEqfX+C0CcAeHJQ50AnU20tS8wsi0DVqJ+6
e/033BeDH+tnvhDzJiFfa3NqkuqZosK3faC7FEVz3PK2TnB7hca6olcEHmYNTMf9BVVCR9Gvezfe
oxslLi8aDK/RtKy92xSssKTRj8vTRjs6KP7BJ7k6tcFWjo/y50So6+j3XHctf4N7Lih8pDH44ViJ
UUZuUG8fyL4Jos4nGhTDtj1mnf7foOVtyUml8gyjImLpYpeeFVm0nMuWmmIAmpvz2RL0oojiQv5t
0id81dE9SD1zcLzI7B69a+wY7qpmTS3wQOD5OvYuFPr4DZnMneT0T3UCZRs7uG2LzcRNdgz5Z5Vu
fJfYHIPDHVaBoB/4x6EF8/AEVDdsxvHw6iGIA0l1stbw5eFQg5K0UWIUVr4LC8Luw7R1b0FIweyV
sZg/N71dEjdpElP/p6S0Djs1zCvEtRtSABvufE3/BIG2OlTvEsvBMJCn/O3haLRjC21JyH33rCMP
L9JuK+PAEg/Hx/ho2rrldV/8URDANL5k61uMZQpkt4ZaKzcVUYhw/3ZuLytZKgDzGk9vON4BzOAA
fKtgFIFo+sYGevJ1IHgp9PWLAK5pyzCXrC+REmAHXDGvphrGnXjrqUOjlc1RZQEUZRKhR7xk9LWJ
7lW8fODhIVBCd8EM7WHFmbxqxdeWKh/ad4vBUUs0izYXSF4uL9ki+yqjQaZ1VwOnIPTsAhygqdNb
p3xWAwdMvQJKzaYrAeSPLs6+5lvOy0jgU/5ySspvqGKyj58Tsrn+osZplJGVUCN0aUg7NLZsuFAP
F1XZYIVP4+5Uai5xBCJQamC4GWY+vvp+KDUR0iJ5NPhpLyz9GgJ5MdbJ6JjVF/86s4r4HC/AtIRG
h86hPk5bTTmvtyek5SBuU09fqNFjmRdfhoLvICpgW6DsAPUDDUbxIaI7DJQ2NHhaoj82f/mKeyKm
9PLDYBGotdzJj6s0VjrOdqZlp2BGAkcWRN3dbbR0GTjV9fqSzEQ46canw7xMPYUGhqnAJanlRDa0
aUnWj7Eh+l5YelakD7o4t+wXvjKj1FnY2WICkzqPP94G85SyGDJk/HudbY2JhYtkPsxqNb6g2nBg
FiQwjcfAGZNLEO8DxCxehEuS74lpadtWnSU2fM6SGqv90MUXkx1oO8abbFq06V/sFKaaoivlcMmn
0wChQmD2zEWwezdAMxzLqBpCG6ca3voV3K2DwmxMa7vJQgJNmsrufxgdsrIdRZl51yWV5U6eUIpn
6gX146gkWDh0+6bHQnsAPnGnYORYWk1mn3BK9xxQGAQ3Ly0DxH9h58QWg00xY15mKc9q9QX4Cq0s
EhcrdkV19ibMRIW4DMOTCL39DJgQvqgu3+KbbP5vwOx/pWakKce9PtInx3AF+gEacZtnTw1ueHlP
6ediGIP64Yk0lxtUh+72Dfbc0zCoUMY4HfRyAYpjcBT9v07GRTgmP7d1kDL5ReRsWcih+zX/pjoa
kIko+t8A8HEjGCO4ilzg3cdPSMVVEikmldBu4YKM+/Yc5cmlb58XyFvyldaY6xUj+NQleCbtRz3m
WTXZP2DmCnMpyOk0R+Eu2WqTs7rgNO3Aqn5mAZecEsPzlqmG44tRqD9ZkCQsdcWbNlMkELeOFBFf
5RwBKPvJ9ZLItkvBiVbfMKI9biNvURuBDbC8pdJaOy2dc3VyWKVJrRrSXNJbRQwpaWXTzYZ4RA/X
FlQ0PmUgAUOPCxUsfk7qdjXtwt9c3BHHR/QXUxeg297AeLt+mFNeqa/TzDBeSwETbwd7WTKMC1RW
1bTFqBjrfNkPQfzgWyO6MJf7boBN/nYFidKJldOmcgpXkVTKKRPvwDlFCBFv64cOEWnRnJi35GgM
LbKBCw80KNRyaRvOtTL0gyqUrwFwc9hxVSS4HFqlAgC6ljot15t6TOMBGgoffs3Z1hNSDb3ndBLb
sFPGpK3bVJ22NrhsF7I17foDr6vcG0CVid9lfIoCfppzF1pzPAA+DSdogqxZ9IHjN44uzDzs7HrE
bnvwEC7+5g7R5uBrZRnRcJhcOgUf/IQeP4lB9IqV7iXpY1vH2Q1DxJx4NprW0hTGkjXZ0M/82mPK
tm7/w4dVmUe7sg2eEJ4Q50X2Sc9M/aYGunnfTCt4JVQNiFSg+cG2uz8RfSB72D9k5wX36lCUOByn
TrRYgwabUyl0Dojw/wavW5Rlj2QfFetD8vKBVAD9KdVTn5cIfmBPQ9RDoSBuwzjXCbB+Ctg2pbef
th1FItRRPkDEihvatr+ZcDT61i0xU2cPcyL2ob7VapLZPYCaSwglu677ed6vlJPNI97Viu0uUuxn
FVZi3mKlN7pf716CLShoa4pFzHm+eRERIUre72mWst7u03UD95573O32ADqB8blh0O2eLgHtvIIm
WFXaXJR40FPSnckmrpH5WYjfarwL6hBiue7zIGFUWdyWLJmVahocPsCCs2UxbQES6cNC2dbc1Smt
g+xoH6eHg7vJkhUaN4/p21yZbBXLJu18UCTfI5rbiNUZKc0954BIojUdFOvOeFZ1VsZMHMa+pZPn
ArTR41ghh1RD/YwEkNQc23Ag/ZBeVJ4E5sNRe/oTpoayxJMvBJ3Y4xTM8v268wif7CCrtfzC+STs
yfrOA+64JBaVUTBKXhhSPM3jyc+X7YMX9HHo55gCpmNgXL4ddS+kQ1ORzDsBXUk6AOjzRTZkw9UK
g4QTbSMS5sen1pp71sTrbw6ctLrBvbHTuT3M6Y3BgNRVdbK19ToMD1f8lQmsOJGX/WUWgxtaVZxs
UwobvWUDXg2NfYiITqeFJawx1M3vatkWJRpVwjIfX+KE4wC10tDT8AcVTYi3qBtqL7ZIU+qy7sv5
sC/BnacZ7HE9l6ngxpw1WXYvx7NxMJbPS/Br8NtyEVwuR1HGT6/NPdN5ccKBhXfnPPvQ0zfHgOnR
OXh9qkkqos34n5UGR3TMw/ADkA2P94LLZ2of65qkJp/x1e/pFIo9fq1c2trsQ2yBLXH4Pp01mIF5
9EMbarAO9rho424FhXiCYlU6BaxX4tRVV8rsgP1kkQpkO5YD630N/ItbwP68Lvis+Fukdzn7t8sD
4da1BFQ23idK+1+8lWvWpgJESSV+gxHbRMee8CUV9o22xROlPxtOtxcGZHqCTFWzZLoP6T7QtIwX
qngjt3kKw9osxhrmqi4himE0yEUJo1E2jpE0gh2bWFSmeqUz57P42jdkGmuwN3v0O+6Kv93QJPBT
wwHCNnb8tsFJRRPScBCjzxJJL8jvp74TXtqiBQjh0inCF8eg0pO2UgYgkkmBQ51fBSSj6BKzlH6j
GV+LORHf0E9FGppOICcFY0beU3i3/nLBhHLuJOASAmyud3FjZ2C088KGTRVuzvJQ2ro1Ss0Nqbuh
eAAVPzkgCAK63GbYmF6FwzV+E6o0++7qY0yAnqvtcVUa+xdxnE3xEzOdCl17zEIDKMqJHTA70PUV
4omZ2mcPv9HXqD0fitQJKJNKOhkASBP3wqb9GcKjBT776Gdydgu5XbwNcC1ViMpYXbON7bOII1PU
Z5YCGpQl9ftifAUTnCi2V7lF3A11f3U+lh1Xp1lFDgmG8m4+dx2QlBKRMlqFogHHuaEkwSxMvy+/
yaJoo3e0HC7Pqu1yBUsvSytO+d1NrPeG1O0nf0DfqGihAF2kHvYfHQSF+FfzVVE4fy5ZFk+LiIyf
Zaa1+McKnOF8MaiE9QmsqJWFprdT0gqI9AoWuPgSxSXM5Tl7iYUq2T0VRfoT1Ds3IWDM7HAkyy9q
vc/HoS31m9qZat/JzUMdIi+gYwHdeccAxsNkeF8/yWVOjzxLdzzpeJkfL9TNasrK5rTwINWhjxZp
qZEmE3Z2vn4r36vAIr8otftM5k+5QLe7EU1IvA46QpKGjtbaADz8ykx8XWgrHF1J64fnkRPT2WuB
YieXe9Aph/UOgv508/XTKvofA18gGN5+5zVHmnhXaQwFjm/1EXufKDniwDa4RZEUKl8w/1NvwxYE
17ZN2QemB8e3Xmr6LA6Ur4WXnhfq5YsRPZdD1MNpH+7Zw0M1wxjVhDEjNe1MalTjNAF7pwGxiI6M
2PZS+NIve6CKUM1jyAqGWs5OSbv1+yCiygD94XxvyWu6XpH6N8CNKz0Wq50i33hWYfpfTQ07weSq
819VJeSDHV1q9UoYfbcecI06QCwnOdxukxB/s2PtyEPFBiuq12sXzQY1jwLxNg8GOglVgUfGfMQZ
thWXfv2KmvRhXntoM5TkBQRIp5vV8tKDcrqEBTnkW05EphiFEho+rkIKBVLIwlYwhzd+xfl/xk4b
8gvhMeWbOGK9MSz690PIgjXMfENReZO3BndqGbQmvJVsTuvHc1Rtz71NA+I4Mjl+BtQQtNCtcA2D
OaNWZmojFoJUzk7ExX2cD/2EQ+g56J9ATUnDwzy9a6gQccVuco4gPDRKyCwu6g7B06hagtP0moOg
weaBHK8vvyK1y0nYJ6l06DRHlIy7mFcU4twTTDv/CiL/ubFSYn2MpjtkRShpk6Mr7CJq3eu0OYiS
psmqJtIhrmOpIV25LaiFLpClo64uLQipzva1+UZHMcv1Kyi6OLxa3N5a2jZxb9+2q3p4BdDJ++76
OhYMM+9Z9OMg8apYi4rL6H32/EbpZfTWWhtYJ+LN+sMZkv9Kv/cLGNSG0bpqd3kwnnP6VvabayD2
pnhGowBwsgwz3N0az85iQe47FXihh5J+KfBj3n++Ua7rICc3u36Bo60DshCHk2CcwiU95V+LY009
LA0UxkXRC8smgH7rcbhfpU6JO41SqWpuHZuzoZxthUD4x5Y5oD/cgI3X9lzn+U44aiNVzrfPGCzB
a6UMf1KJfstnwPCA+YX/OUVGE8z7MqErONNQjHq+bzeHhTRi6H0vnn99ie6OdvTb0Qr7+PraCQ0h
ZtXyjIwKajP6zZHP7OH2Qy/98mTk3GMydHTjNbOGEjNUg9QjBpFc7G1Qz6nOGSkcqUuEz0AWzy3G
Vd9lCKghmdjwj1UjLJ4MkkUnZSogh6zKkGHVWMUhzE2pF8QjY6TyJD6USFt6w4YRfii4DwKMNtfS
Lo+GL8Bsy1xenguEhIOiCJG0xCHkDW/MRsKV+q0iKyd0fgTuUPknZdNhyI2JXcnb78JiYmVkhu/0
NQJYQpPGlQQS31D9wR88FXY16vMMLA0kP07OwXi6P+WZjZ43z+/LhQQJLWrJ0/fDvye/ULK3uYf4
Yyl604CgZ41AcgPFka/6Q+t7cDAxBez/TdG+X47+k7H3MV39N0KlEHGan/LV0g9nS9jMvQZEEYE9
YV0TuMYqdVNyTlF/ypPaUxzdNNC/05n4hsuyFidZA8/AvKdwEqyKNAxOAvriB52ShxASnvK4YiDJ
89sH2XGKhIP471/nvbJiKEiX8NUrxBIXXnYjPJl1ZeADLLII5nDnsGjvMS0ETgZ15lk4ChnoTNrI
l3nKsYnwWPJWMTwpEwQBJoHXVjUl9FW3cCUaJ+OUQGKFurXHa8NHmgMys7jLg+Vnb9cTF+E8Si4J
MxwoDCDBQlD0s2ouuslEd8R7C/hAKfUUwSc565s2Q3SmUjDCr5/LNGletpkFwEtRhFkOlgRqfkwa
mDP3MT7KldSLW6WwmCp2PAorzAxis+OEtmGsvjoMpsX7OwPMJiO9aHQFswMiP7G/4FGNNgNMpj0N
immFgeWPSt6xJ7d7F+zZLW+HZanyMXz0Vi5Nq8Z93An3iKUjiyrYPSYeHYrJZfTJgEOzNAfsZqOf
ijRLbkMcEuC66mEkO4kXUX7QfrXcNljfvid7FQYz4nAti9kSH3shOiNJ/Lk2ptKBTXhDcYKX2u7k
s2zb3moh1MtxMOJil5M4P6u4XYcn9iVb7Go0lqbF9fGaY+WQBjbHtlovCevJyTVb/9ejA9AZGHk8
l6NgYXSq2Zr56D2+xF5n8YLgoT9nny119nK6P/YlqaKLOi2vOMJfrFqge/NpI8q+Tj7/n4doILE8
7S4JV+gQ3WlDitzBsrwuByoTimkPYF3InBLeXkpkq73Ni0E2Vv9+Yry09jDO4yNAixnz/4oSs5G0
XSDF2a5ziCGkhW88ccp2s8XnrXZ7RfvRFw/ZvZoFb4TML9Hn1ZmqVWsRZcTBVBbkbRkFttbS1tXi
CW3WbU3fqjaDQIT3weTwo404NhpBnlkCOjr/DuZQVlcQUTpqcViNboNvkN3iac1qZNluIaD4Og+i
6JtHZ8021Gmx1vKo3G2Tp9jk/IX0c4VpEFVCNDPROxa3mZvdHBJXpstOX4my5x0QXLHXd5riUWU6
oySuOIR3qA6OolrEXvf1j/l020gniI3/mEpeWL8Z4kGUepE2QwBwCeqfGs4bTFaxwnR4+P1Zr7Gp
NYN5ePhKShLQVdheMKySXb77fRDWdYdVNO2Cpdq5FImiPUGdmxBn7krzBd5/sLS3H2AT1uLwlaJV
YthifHXNsgS3Y4SH3+9nYA/93ZUPXAjS9qk23LqFD+5Clyohf2tXlyZSZRrsEuzgzTQGt03UBm+P
PFemcCvgr2nZedUVPrt0ANdMz6trgJKmNVaks/Qtdn64kVebteuaEBZfOJD3UvFQPp6JcGCQpnZ6
i4SixMSl2xgGv+luPXE8RGtk4gfgI6WTpTGDRA4ti+1MocUFt+ov5yxaebkHUvb6RVV1Kxo+76nu
kUn5HCkJOmkPMKxftekXcK4P5SZ87q3UhlbRbBHz38jLUFpFy1Lc4PYWzSYqGrVNd84g6zs2gOt3
/mMYPTD+5+PkH+Px1DAoSymbZMbX6NB6EidQwsrCEUCoAwKtJRRE7RKzFDDgQTDyy1GG+Q9vxeKL
wPxkXeacWIoiFH5PSMu+kydtmF9IOgP3dyb1ngIoYX5fDIcxZl6KuNrSdHlMm8g/DmIXpYetaJ1C
/gfc4dYq3Jib076WwyugmV9UYPNKJVpYvWlw5sjZPRBq2Dx1CWLuaqu5BlwXAYBSWezFpe51t8zf
y8/WtuLsIigPTmB++H6xXuQcHV8+QC4SbjwOmnTKRCiCyvadoouyIbfqRx8riNybWsJhPnBjUkkl
7hGbuBfPBV/fi1EFGmg1KRWg0m9RSZm1shG1da3Ptq9EOK6EAGetGfkxVsXdHacQaSklyJ7+OIsT
+2IIbdf05ZR4rDQiRCJiSwYLWIsV6+ZnHxdyI38lVocGn4Fxj+KZZ/OCT9gbeaAjeaCAnICLZvim
Y7uEDx7daiWN+B/U1xVCAvClJi8YZuBUhgXEcQhonTm/LJZo/5gGcg08Wqrp4woPJoBRqjEfasXB
pZEl2gtPJO8m4oqrQkVRxHuwVBc9uDCEHCDm1qUjr40uSNpNC8MsP9XVb7GNfNQdrXVofQGwD3s6
S1UXc8N3CmhpHbwRnLNlkssJvogmHrAQHwYG+HYiCr0E3f+SgCQAEKz3EmTHNbHfwZf0jUq+2OkY
SKWPZTk1mkTSehTGa82qWjs+gD7heKFbq4ihGhfvoqrsxF3Rju1IfAYgJfcDRmblfhY0jnQHBwba
15C/q/TYcCV7OCOkRKQWY4i3HiQPqGSp3O5sJlgRpMGy6wAa4Iz8Dg89Qg4J+Fewq7V5kEbByHBt
9wIXx2EGXkHVA41Edc/YitGggxv51JLN/OhbnYjh0VIFypS5geLAFSa3C8wHPCn0MLN9oKE0USHw
3KLH9HbLN4xB2FvWajb5X27DqL8JaeT09daR5Gudxockv646D2NYMa6/NogYFfxQscR77GhdN6YX
bCUcwzkwtrN3rfFDFUo6IqwFEUeWmScfuzoQ6n706xcb502iRYzfP5SdD2hZG7S35TStR4o0B2LE
hWiEyISOWMAlF5uNJ1a66ZSPRT6qSujy3wRQsmF3NTGkXdhsOeSLY60bjWpLp1iUd1s04evWRVSY
E7DlyNcjgNHSr+17pvmgF2YI4zNpwdeWOg1cSLNSDIhWye5GQ9j4+EKZW8mWTnsVvzMvgdiXiBor
/4nBtJ1SCXDKlIX0Wonxk4cOzvgf8XHRQvZAQ0sq4EFPrDpGQk05SZ++H/wUp2VYuu4+SLPCjU0F
EeBldgIyl1xmET3HZXt8DEoXX4YF6Vt/i8DO/fDM7qnmFR8Qi9xJ320PqM+zWlx03uT0CS8tGnPg
PLGaXSpx/rWi21+uY/AIpYvKwPlqHEJC9FVFbfD2+6zcm3JmEyRP0+mJdwDHG1U86+JBLH3CQzTQ
M/T4z5UcYl4UlgL7ujAcKy0QJE2ptyrUtMUUMWt7Fr8wPOvjaTugAmwqakKTH2Ov7AvtP41b6OqV
cOvh4/9hr8xT67AgOJYRPNYzWuIvH84yCrD7UVteYd5juzArtSIoKsv+DCRC1vlQicDS2PhwU998
U9BfuAwI+0jyWQO8HAu5CamU27H86g7l+0s0FkZUdndg3mYE9OZ0fumb0yt69nURnEBNjcjQ7OJC
m7IsrZ+xig2OwnASlrRQ3cP+KYnileoQa+Qni9qA8tF+4/TaNum1+JCdNaZjjl8D0TzXeCfVneg+
0sPyit27dnL3cnHS8/2xgMWP0Y2PeOfNtFiHM1S4TB8nWvmPc8cPX2O/COk8g/ZKuOjVqJOpUCNa
KxAQa8zhnvbKyA9Dq3dwGJHzpYm50CBs70QuRN0CaveitD39ueiFgeufemUJT/fuReTVCXdITBLZ
t1vP5GpN54D4JN+PUbZdK7J8NgCZLIzgiRJhXYl0kntzq0j0y4/suk6XFYHTtkxql7UzKpdd01z8
t+LjumOMDsmVBoG8uU4n+Nx1rP5vnfphjkcJBRjxcm0IiuftkUHoEDY7Au+LkOcVgi4/YN1eg7VP
secLlR4nuJejh8JFMGJypXsetExLvwq7N6eqd62A6tUKNgL8EuaBrerZOFktoC/HZ/XPw40pRQay
TSZgMEruG6a3brlusWajobf5CTx1yizhKZOczDN/Y6bXdjuRajY1ZdCk0C82hEUw5EzKqqEU1Nu6
Ohfe+ILDYE4WFdPLR/WP4564fLU4HPY892jYk1EOBUZW10ql1XBfPEPKwlKvmREQB3III7MB/dy3
eI50gNthgFuIBi8z6GTm5AGAYE9jy6xwfWmRexMdgMZELPxiJcpKeDCJgJ3fe33xkqhJozQCqVMp
5/ape7fiuBRff9NSlzAeoBlLKx6/41Xclug4Ps5g7s5ClG/Ef8AtIBhhjCX/d4+2MOwYdx1Vro2B
SYZe7iLIMtu5rFOPZo5pNm38I6cN2Nv1cGvQoVcniS8zuvTQl2bMn94KBEV9Oa4eq+1eqr1nsPk3
blHzZyjnAqg/8pVBQJpk5iu1CRipFkm3SEM3QEDU+EI8LpbzBIs88RQm4ZoIJfAuEdHgTnqImia0
kHrxFj1JbpYNc7PfXPRMvV/lowffXYYoR77WaThbrYqRItKmt9m7MrPd2m6YTGBGk1PQlJoT7knt
jurTtogHxlHvTlpI52ykWYKBfAlOSvCdvE1z0wlj7E4Q4aqm6EvrZ8U28BMpu619W0Y25FjV+XVD
egT11+IW1B9szoRtAvmHQ1F/cgUr18sA7YFBdIl8gLtZwVYnvU2KhB0lN5F0uCRcoDB32qC9oB3V
2Iou180R06sd7cYAe2PpcLx/uxiMIK9tI2mLT/kSk480YQzsvZq0yHbo3N6z9WNWtBrLHyWutjs3
UkeWyWVfjaTFWRNJSqRlzKBc6C8EBZnxsUfE+xIn6BQod8VCRApeSrnQmQ83uBttVrGBVOcazWmX
TR5x17ZQvc45zI7NyL/HheC//JKE0bpD5eNz3/JahefVjq72+IgvqY/hBkp7zINm28UkyZqotgP4
yMEcF+56QlQu2Gba/emOrmuRZdkYPkbu249C22Mi0/WreIzvyVm+W57OCfIj9GiWMliEnsOEe/iq
euUMMjPBgmuKDkDLvNfLddEhPX9ing4rHfBMNBtpIep6vF++Zjyl6paJ9syFw2rMQnh1lNcg+sMH
D5DyrF+XJkCWi8y6g0cqCjEGaKD8KWABoJxMHVwr3t9RdXjF75M7JxtaQIMiio5vue3GcZXy45hg
hZef5u935ff+1j8Qo4eiSLHKgRk3tlxjgwFROqLi3TA3hMF0sf79pk6Ix+Fh23ql1yrp/ZsSe5gK
UdPUcPQbv4YSTe2ncNTtZeKR1gp5dfxHi7nBf5GwaW/2gyuO7wO4aQTK6zTH9IzDtUc1ZueLV95U
3VvJGNansfZGIWSUhM3/9J0/06QBBcVnXewet0o5BZyvI+aWGkNX9riCJ6H8xeDM8havt5MCcHnz
zt9wckENGDtc6yOf/j8WjQLoW41tI1mz93mgAYmVw2/+bKhQwXqysvbPnfTjNlLjWXTXDT2JMqqp
pPcWx3NNGYbKQsjmHPCUNw2WXEMFLutFElVWHI0SXj1HfURIiQfyJHaR4+eAdBJCMwsZQ2jLtEoJ
ETY4XYPFpLl3fQ+qTxzKjNVysrxgW58vrbqPItSktVjBd87qncucVMuy3ufb0WrMp0y0DR45Um/u
0EpdKeH9bkQ6Bn19vtaK9BdQhDaezdbF4whaiNAn9WZ1hp7mNgBoKdHemEgD2Cm4P4TwKZwcei5h
yulm07nWXOlSoLOtWuA+XgqxD2rEBqqIXqbFkAZorwT3iEYwAI2I+y4whble3wSDhQ3B60zHwQMF
KkYmVAFiBpGQ/IuYVS83R6r73HEWyttZTMRvKi2rPz/14NE0alXeX530osDVsuj4F7r4gupyGYjQ
GrEWSdYfMnXx0dixepdSzkGnZBUHhPyQiU1iEsZkjX0YM0MEkZc0s3Fj+vfHjjJfINrEIXdACKDB
R24fgR0YUOkQ376NjuRTPxVMp6lfDh5mDzWtqVjRVtBr6KOTwkCgfOoQXf1DYzZjRllm9LNZ0qpU
/b9kucMF3nidMfSl1jmjNAGc5PIBwrOdO8K2jwp5/LbbjwqmiGc9dslrP/zwHcRzzMZis/3uLuQ0
3ScP27Je0+She9PPaEwWZLET/slPviwQSge4YpoMA9WaAEEqgDVFoPIBWdJWpq3lQRJDAjTZGm1V
5pO+Vot2yADix0kjdS95gbRkbM21lTdDAYiz3L/5+zKMF4+CdvwI+Nujmum+ywZ0hagMQhxxxSNW
8rEzR35uisBf3Ta+CQ6ER9rrq3uacor4vjCMGV62Oqv6HGBiylJFMimX5phV7iGStPM4qOVd19wo
+tDOkck2g7DEzIOaMQHcnRqIR90+5+2K9ZaZk5uxZ6Qj+PevSy7532/fgxwwJJwpNO0ijAJ5Ujmv
gDGrvYaSuN4PODq6gSnyZggsI8guzo+pFvTQwULGc6CJZ/FCQMBDdM+EwKTBziJntv4C5FeC6+6J
D6s8B/NslVD2LK2/fVjes3BCzAqujBHUACVsu7bp3EJLFRVOaIGbRfi+sioVZrgAV9jMCYJlTv14
5ZbKEOt43HOV1MddnLpHXD6fK+Ux/Q3r5kZjUlQnRU2PIlHOzZOrfbzDqR+Uem7ISst9YtVLNl+a
FZvZQO8AJ16v1Ieknc4S0vZ0brfsAI84o3RU0o55A5KnYzD7Cto316C/pctYfdUlEJfkHkwjadni
Ar1i2Ko4+MnuJLeIapE9+zVdg3VTsPvLFEzowbNrLyD7lPdgnedSQ6zRg1QpeSVUFKdRbCKiBK4z
jz2wRSIKLsc5rSG4M5kK1iKz9jMx+gpzBHXF8GYCHnS8ACQCJu2ljzmPG+ODzIXrVzhrKCqqTTJy
XfGaWqHRKSFDvYX0rCKf0XKdu6LF+XRd/B8N1VbQviSq4QdmlZIkb//n0fSw9LIHD2L1fx+snVQb
3vWNXzVg5fpVu/YfBNp1J0m/xd4HKylqYj7gA9Rf/wlAJQfhSgiSFz/7eZdihptEQeDfcbY8GBuv
cLsDRGwtJKrQBwMxSkUCwTbce1sc7dwDqAhoLQmiEg/hbw6qDhLbuE7CEstPLZaUZRFP8Ehs4Zr7
QbMCk++yHiwa7Yj3voNwiTNbitVo36DNVwSpArjCNIZ5EHdxF8WA2V00MUmJQ7s3J5B0KE+QcNKw
Ci8lRVoi1MPT8I9SBaDnC53C9RbJGZ6Xs+46Pnsc9cNo4UXKIM626O19OKHxIOt5BGB6dVmQhRTX
qRqpeMItDSL5/AdMeYe7WsSt78rdBykHvLTW7kqvz2OTscxeEy3F31V71IsKFA7mj0QOYghiIxBO
QwdtmKSUE04YV0cjqUH1cvfwGn9QChkYRqtax8Dp9wspFtDrxYnCuhMNthO5/L9YLixZjIVTKOZ0
oGb0n67UCyYRy5Bkp3lXKtzIPcH1UqIZaa42egn/FsrlrDf3v7hnKL7qu4C+bM8Wy6vg4J1a0KH+
Sc7wstdvh6K526kTVqCN1phWhEqVHGwsjrb4kAqe96G+NrGGLMUhprC4xMKbWOPImoyB1ccR9wem
jnBNk+HRc7NWZxvSMjd1eh83F+QVINygEYH/mUfLhLbmk4Rsr8fiOrDAmvE1IAQhCzU2nkA8nL1v
55Te45ULacVwdeEp3DjPKJ+J3PfwugCBKtIqmJlEz8LLczCN9jKH8bCvX4xvymEajTASXQZ0JnV4
9b8YdAr/v4VhHiqRemT7cDyEiVu4/Zl7a1r3EDDjMVKStFH7xJzeESRQluy0bUrI53EdzZwRqjcb
/Z10eI6uT0VST6o/1HDZRdjudKFTuB7DpPktokJHK8YXHfa611y6Z2XAHsfX13C8ZltOqU+TXYgP
eUba5xs5wFahSLJ1MIrHdDrLbhmU+1kJApG8zdpTButCFx9jCQyXosxpw6b7JgxHyZAqf2M19McP
LsY9mf5LEkDelOYG6VXfpAihAhnNlgsZ0jYPH2Iq8uFaj/mTCkJWXnl/dfVVvvirCsZq1Wqzp4GI
L5K/SUFOAqqhmMtGH9+DzBIdxLiPDdYv0qf6o8sKnybkLcO6pBEsYytDjFfAJZnu5uT36G9KgPFw
gwiz17CZZpqQN8fBQP7jCitXWumoCMttdR0RwgllwZ5wqmCmqPZS65LkTSlFqerOKON0PLv+HUCU
YQSe/pKesVHC6l0Zs+77ZPIk7b+eHgO3JWNij1QewThSTIS4x4nKEi2+3u+Eu1L/EmzL1X24TjB5
lkDeZLTa85OtPb0jMc8lJOOqWlJ0g4S7gTLp2I406Hf8AOqs+z6sHEkF59xR0wsFgss29Qg3zHP+
op2NRLQeaLn6RnNogaXXERZ5A1kDtThuZgvPo/Iv3s3nrKD0ALfeVVUrr2xwbTpqE7AKIFq782kV
eIFWgxZKWXPo6lhfYreLqCYudbfkLJHk9K7p9mAeMORmYSYsEmxBOlpxs8I01qWICXWTGzJU97jc
he1N8JkCEKzDb1R1f57WTO0YUu0+4xeo1EBWdjJDsOz7F/3gQraK3hzbSxJddP6cfMkS1/smIByK
KNOwac5Mtignq016iFrZ7hPKbCPpk0xkYc3oE/u02dcxWC3VOdsqG1lxfsbnomEeFXWAUVEVmDso
LAETaeDbhVxMsHyk0RiRyIw8xTItbZ2S+u+7/COPtV3rnbOMcfnfl8mOC8w95MNtTfl2r6IaGY6v
p9Rkpb02+bX0VM9pHXPxbCCyu9LO2eU+SkvvPlWctQ5pMlIQvi0Hk8+POKLzujNDwR72U8RHJs9C
j7JO+nSKpxdp0gBYIdlpp56JmlqDh26dvDrPdxHJi3Bc/v9PFW6SGwHa65Ac8FLFGdBK+gRaYVtX
2SYXJi5zBxyPBWTls1WQ6w6wdOhSwlKApSZAoCInq2YvtpumRYh2gvnoODrplwHh4TvVZ0T4jyA8
XblOsv8yI6bD+uZkgnDRku2+ZDQIZQEQqzjKSzdzyMVMsTcF7DkV1HBZWZrcjcHMvUkIvy9Hx/zJ
cs/BHYbmV9BW7hno7eLhD7rn4r6zjP1dsQjCizHsT+zXwkEY5+XuHBgXA6z/BM7lwz53MfzoMIJY
OiOCak2kIHCnhmflbErPqLLbPNUYj+d7aaKmFU9x0u/v7MqpSBGTHKK7pjcLJcQwol+f30Y6IkS5
0winjK9xikNuOivd8R3lMGMkMsA8wzquO4QVQ9yGPJBW6h0LdMnxLie3RWZk/apjc/cxdC8Cd/yz
HpHmxRkBT2OuP9x35yCzcQYR+Lk0tLSCG9cft6YBfIW7o4+XkocWc6Cg+VU++xEDhluFcNZoMs5Z
GiHhqANNCPFus36tLaV+7NWcGkuJ1KSZ4RQh3fLAfdhVpvgt8g3elvYJdWsjrYL+PE0ljiNXICed
ijjMG2Jf+3xw7DrIHbtvC5W0/XHBsjAQIAGmzDOUWW1+M6pX+mNu0/fHmNdjSUBiPnKnQL6m6BrQ
I8ZltW3ZanRvPiHy8zygu2xaHHFPGWFtE76o5cJDMLswjjJKJAqO9G87ixA3TqDOu6wEndjktHUN
7FRpMJIsp4WMUzT9U7O9uJwmEYI0+aC4lWQF/shq7SxLgPo9HkzasZoVji28UgTIn5zmjCs0KpIq
FSgkmr/eqitaR3BUKTuBL9ebFOPIsQGvMJTRXDOIFUCIN5mIt7QKA6JF7KoNxeOhXdceRjWhU9D1
NUCOLoe7xLfThsYtO/lwoC38nft2p4Cz6wsgI97VhpgPVzOV0QR8TW3aQjwSu1PxJ8y6r4ju3wbe
BZo4CRwo33bsg8N+uw2BQDCTZjTFJDDGstlkHz8qIspYoOOm0+xqiYI4d+nOVHKFgDKsjxRD+kZk
di2kZHakFvPIbSYftrxDox/d9a9q89eYE11vcz2M5e7MjWb7wDsC70Dk4vaTHRdHtQzrjNYcgLhA
pDOszGsxX7mXCvCiaTOu48NJzJqfg5eIcGGqrHxw7axH63V5aG5IVg1aWIy13OwLxVh3BJJzIizV
OBzWYo90G0TNAh5Iua6GpalWBsIlUBwc5oK+aE+ycieseo2tJbjzGQ6bJQdrOoKxNLES1FoNAM5P
3cl8bkYRh7YQ5iZmQTxNhiQDupfHpcmwP9501xWmigArg7WVtDL9Mdq/j/FUXJlNr2+wRXQt8cQV
KLiHSCnFfZn5RYCPwPXxbyw4oRC1jGuD+UmW8zv7eM0sCF7gyK88+HP6i0rfbk98bS0njtqZB/eu
LrfqwmUZrg8DICaO25R91/pvNs7lI2TsHm1pAG/v+r/mysR7CKFEmu53E57BL472vqrXJsokngyY
q5UVOAsxLWjjx+ReNZ283oH6LuPhlIzuRlC5k8k4KboSQ95dvmNjSkno1VybRH3RJgxtnCpWtVRO
Ze5lFI6BqqzQOOjKyoZNOkWAZJ1DIPJdn05rNnjwPoqk+xVCq8pGgpAHjM62qcBwIVY/nDpg9/LG
sAGFcOF20mgiVzLU+cRa4Ym18dY86fpdYBrnZSgRdwhuHdzBCXLqk9k2VoKO5paFGqEozZWhYd6r
Niv2ymvU0TCt27yfZnUlT3s0o7mCgk8eG5Zb9xuyLfBNT3GIQHjkbehU1J0cYW+KOoiKqqusEYwN
nPLtwVgwLRXQzL/TW9CZfXy02dxPRxbZOzi5tIqnDkm/rYPtz65i8u3vzshF/bfj0At1pBxcqQzr
Pg9KxmVG6jf4hqKhgx3GyTrO7upqaMEpGem7Mdv09wAPFlcns3YXZbuxwLdsnHIiKuduxhSbhPzr
SCzVwLbju0YEz96BbWZTKbFQJ9I3mwqBHX1k+pi8wgEK97T8Av1zA6nUNpi0br7cksdhQkkgQuk/
Xrd3vLS5sWyZV4pv176TNrRBBT90wg58XEKhveP98IE0w5FiXEjUPaMlzl1pxNng2Aw6u17KQk2f
SrmWpzOZgEvv0dY0QnNgPbAFUOsO80Tn5a2k+bLXb2D3envcZcyX1A60JWAlN5msqF0XIE0t5hc9
JwjmRodQpcjAdFB2RokYnhrW9ZBEv19M2LL1vaaVNzALdZYIZUezQlNmPKgN85Ri82J1OzqCowGR
dVCpiM8oq2iqcM70CbHdrmRgyjzHV4CGgvtC3aC98706l3NDlhXqsyI60icUtddh5PuQfU4EXE53
yL62mxEAAGuvkb3HYvHdYIq4SGuYd6ETdUVAcpEXPm5PD/a7Amaf1+4gZ7nMPr3fkSp9SdIElb9F
tdgMeBwKNcATEWIabXuJheoTTBWAGcjDEjsyAK4tohAWr6PFKA4JWLf/97EuB5OTI50tdOQUqo1Q
b0EPct3z30uvzgLgRmwTL+uABNBvYXOXf9cHTEGijBUvH4aBWKi/zlSNUgFOyMCz3qvWrclZ4Elq
/2MShC1PZVxpqfhbOF1i6P8WPmgKwS1IfwMHiBKJWaadi4ljjzfVYb+6XCDapL68BOBwo32HI7wd
si/tTjAk0AlTiklO9dnN3PAkHEW1VK9I//r8OSLRxH1WolpMmuYIcYFGtEn6xITuilDJFKOuHaGk
s4r03/bKX9of5Dvzu5h8nFZM3TbsqSIhUbFas3cg4Mpw+A80Xxr3Z4Ihho5dGyJRjUzAjd/5iMvl
88r1/wN/R7WrnT/jgzUul0i2BeDj7ulpr2OGokAqlM3q9cvdzmpn8XFuGI872VdK+n2TCL5xmnGp
5anw9cbVS8X4UWucP7sO9v8NLNBzpTPycohjbqos5iwqXAYgA4hnIP9P20TmjCFnnqKlixZzfx/7
/0qTl8GT7Do/xDDtIIawc/P5+JLIuUPXacPgzgtlVEZacg1U+zIB0TvoaMWyR/ggUX9GmyhTXd/x
N2XBx39giQqCRX81jP6qHht7u+Img9K62ToS5UioBOELwd8EHO2CqtHfAb+Lm9w/os0GO0CJhmR/
KgAea81Ycf74h4LxG5uR+43MCRCYeKky2GKuo+ZAwkzYQ/CdnRkHYdB9pQ4InUfY0pVVSNLMgnyt
SGKvKgJty8MIa/UZSn8r0102/GuMjSyYbUn8CtwL2wexvvnH8zbOyVv8fxAKPw9da9eTtLicGoIk
yzl7pR+lebDBUUEUgepWNlbJfGZ2ohK4EQHfE7s+ubywXrM2TRcpiZYcYqlPXFC9VydOadO5hshm
xRfQYiHo0xFH7e0EPJYpEXDe+V9Vv95epMPnBuHzANl0VcQaqpq9kxP+4fuBbZ1W7Jbwux603FQe
b3IaWTCM46u3hbj6Ek/g/TURcPTS+x7CZNkWFJZ0mXqE+/f4Sp2wM633RkZrudm/6v22cX6t731w
xsjwjtaRU5/ovHo24kM4HEAeEktNSeMYLLjzSvZJuM/jfI84PkTamNYnxMOd5R+O/0fovy007aU4
gR0pIQhx+Amvl2cUQqz8WerW6+MOj8EWx8NcX7jSTdhkKBWW0C/VfB8iKjeactkRdI00SD5DV2NR
ENLZHALZuOFOiB7uXxzs8H+dc8iVdKekJ4irDscxIfCm2NL3PxyuAs40C2FoEtumrEzIiOa/6Ygu
DQAv3JmTXS1CdbmSeGw7Jx2XTIIprZ7zjpo981QE71+9OmyXJ5OoDQQs3aiGJ2pJH2GGaGQT5iQ1
VVey7J0cRKHffrg5Ikbotmx0TGvPJTWkf7hHtFVMOOmn6bWlD24eUXwIwwGsNGoqj+D3XT8LkslA
E+/h6HLW0HRoRg77GoV3umC1MTk0X+lQHFmhImzqX+LCCRku8tVc3P3IFOtwU3qfzoWnhmEX94rD
qU9Px4AQ7RuquMz8q5dp8ePlrfzQPs/QTEsaaaVmiwVbVFg4zN3geA2d5N/Ff5tnYegALZypnpKb
knsDdUFdNTvfQP4T/Sx1wq72+G0gZOe7OQb8vyTwIeOG9nWv+TsIubyCl7o/yWKGwxC6R5Xp0u5V
kGQ3JwOL8tvKxQGbHElupgBhFBjgDyHnNVF0j1wbv3DaBZpLof+6Bk6PrJhaWg4XskKy4tGFNvnT
D4udEMK2b+i3xvxdLAOl2v6o0uaIUNJDmUZAybvVX4XmbZIxbtMETR2fAXwiWNCccbkEKg1XaUiW
agO/iUjiJdvbJ+ocslnZ4N/ak/f0qVohLn+OnIB9JnhvWaNi+ghRY7FkEW0hCdPvcYyXJ4+l+EJE
zr61DAXrceVBEzNH+ehM3/5CiPTOoeZBtvxQn8BDGBvZyqMEgqZruraORPAErJqNLrdvCjmkhAsA
KkUNhqgDMpBEWI+hXeh/xsawssX+i6moq2N5/KSuOpmLjysc4AtNE7mDmYPCiMogud1Cl9A09lgY
Pja9deSG5sDB/ALLLv0wumHQTayiRCuM4EDc/degGdNhvS8s4ysTtcaWbr1bvs3dPgRph4Y8heqf
skin9x1WccWF+OQ7lKMGZc8eM6I6WZOWE4+UX1Kls78vTYYF3e/gF0CR7fAM+z8CZm8OrP+KVeHD
PKAnyUlHTtFTsXn8YCOpQGQ4nqqG8sMCvTN3rHzWIMtSrWOWG6SDGywwYkt2gI2SAqIeuLBEF3FX
UuvuAzP5yYJAuuqeO/+CP5IkK11XnprWquda+FChrIEW2v+vqJhCc3UlXzQyQYKhdNUD06IVVkq/
VRe3lX4xEMdoArMMX6e5mK7F5cSTtYV2LMVbTrgAtNPJ8dv0knB3zt0e5BJSWlux266ndalZ1pRi
rcyeNlZZHl2aPPJWczFq73eMqzuimBbSht/MS0yO0ixlR6fxl+F5oSYV/39uOgMStq2POfgdR4w0
2E+aWHU624xBFbiCChqDsFh9NOznvzx8TgUmPMlk+zLmFfggLIF1UviDbafA5zEznyte6P5mSna0
98HOQZXfLej3sPvGC63pnEsgBq7exlw70ZWGwBdw8fZIBPw5q83bY9tWZ3BYie5vPY+uRsCwRIwG
70m6ISVIX3mcnQKPgd6yP3MmiYOoK5R78GtsoCkBwvEoOeAv9JNH9zMzSvEXoXTB6fPKgpxJ0fwC
jSBcKw6cC/ZnW+KBf5llq4Ge4Gg6FUNqp32C8dqM/iGRAYDqr1AgNilUVo2zgq8NBqooXdTZuT4Z
RA3Uu5xzE6LAJ6lM8Gv/ed91rqqEg/rli1cHimwCZ442uC7LxNvFihqOcftQycAiyQNsWlPOP3rr
d2PtR1ev4jUV0YAPbiVTxo00VpTilhcYB+YnljvglN/xxKlXQp4+PXX8CVPrOxnXsWTTQULd/x1r
ZMSP3kI4i7+QVUFPAI34Iel/JcB1O46oj3Cnrcgp0YiRSwOUecuMw3yL3Ww7XDqoyatP+bl4xEOD
zOLbh5PAOowrk17pGqoYVCxNbv6qfCXBTa96iMFOa8vNCoFD/howU05H6X1hBfd7iqXV+lPOBpyh
rykaN6dXJnwIB1xM5+RBg122QBSpaJZnkmkdIXwVzwnJeXjUri/e4eZST+HoUcXPzU2kxFQSmK65
UIBadQUQvlhWVxGmo6Kf0Rgx3ko7qV5S+7RRnQuSK78mkzo+ZBZGWDPagKjsdvczDqkXR6jvp7Lf
nGCj+IKnN6o3RFiTvPzT0dFzP8u6RkPkdGHUQO408Xao8l55Zq8NkOANVsahaa4Pgx51t0gVo9MG
FiSp5AISlposohFMWAEPSX0IjEDcSuZgA5UejS1GYFPmx7guhYHdfw7MgyeLtBm1W68h9Qlc8wnM
feUVkZ6Fo6OHwPZOLDI/+UAJozm5i38dMgCtWFVH/9xE3c1HOVbrFTzb+75n3ZMzdakX9hJZ/Gn/
FQ6S37R9U0G5OkhftLdnOgw1ulXyHlcyga8XE6f9eD6Ov+kccR9O/mejjspPWIJ5WSi5tNoMDBwu
x+d273vW1XD5kutnQCOrQh1eZybPYEyjqEkBXl4Z1iAxqW3hGpR3i3CIJ+x4fLZk9RE0MD/GbNc6
lPztOE2XZQBvNxfMCgF9iZNaEjnSvA48Y3Q53h64jG+YM5lGP2CPAGACZrI0GGIdL0k02qS4MOlt
eoo2jjOX4GpRAO09KLa2bdxiQwKwc9SUysUANSTCA8tNX354PHbyjQkkUfWKabOVPkiTVhPffoGs
iGO9+YTHODXXQa4z9AvUF8NpSNHW95dqdtPeZZUemL9Dgi9Qa6qvwcZHfXX+P8r4ixGrWO6C0nnc
RVYzJ/GpW/Vi0kHfT/S8cXmAXayb8Drz21ubwy5pGcYcl+MGw4HfUqtPq1WdLo7CgP/xiN7NpThM
hd5zEDYq/RRZ0RAytH5WOpB+gqF+jN41R4PIdDQRNx6huBUgy8fMRGKNhHURPGPS+M/lF7IPFkkV
iWcvNkUDzB0j3m4N7Emrqw1LS6+kkhdVFQMSmJqIP1h+Bgnn00Zctd4Uolbw3ubvQaYs/pbv8R+n
gq1jEmhtDHd53YHJJ9w3hXHvc1u7c04s8HuVAtarqmPFH6sG3hNIo3oJ2MLNPRtW/HoTR8USvywq
r6GKG2S7AXGqvAo22YaHp1vta1CA6fdqn/hc+zbMDpYgXH5Y4ElBGX0cUzCMhmw5QyYhikM5JKiN
au3jNxk++ajmKnSinac43SpQatrq9lz55Gj8EhUoxLRon4yikj+9wipA+F9A8r6/GFftRWrEbZqB
8mZtafF/7Jz7F+7ER/v9k2FacCaYhZQwsfkCKEJTEviiSbBmddXxMckMWXXdWbVIysdZLoiqoK0D
qWOQ7SEVeNoSjJCPa9dEsel16hAcnbF0feaclHtIeZMKRw5lISgnpuxXRgLIK+RcZw7ew01aqe7Y
6YlKAKOxmXFLdLNTtW6NpcvuqM2uw0DlWke1tuBMPTbyYRE0W85zKn8nAAROreyygJP/aYy3PVEU
op4wcAqLVwoNp+TBygRGnrlGO8MUNcdlGNIVql+8gje6dkMxsGR2wp0g31PKXaXZwqYg1tx2mNB4
kVV7icPVs29rVrmJEvMF+EsasDkLnuTMAwclRpR2PJpL6xqBjc2X37g+B6hCyU55+lGZH+n7rVqj
NgUOOhuhXuSYGIG+zJG8ymkotuytdrfakGZ1yLdNc9P0tJd7QVseB+OtTQEuqQzaRoLtFF7tGQa5
+SKj+IlhBEm6KPGl2CjE5nzKZwm8goV7Cyx6R2zwHGZb6rAD7BQQ+HxCHoM2YMFj1/L7Cg62J9eR
c2zMhJt/bRMNdpMMY5ulZD3+l0INg4IUUIlBVGQ5D9l8t6HcSje2EfXMiUst7IhFUYgroAQVlvJq
3/B1I0dbVK9Pj97pn9bABTm3L20cOxOddBy01TaNW5/8r5P7iUp0lTC9iqOBRSHKomEkJd02kXNs
VnMlO+cbFIGArWhiyE05xEr8upLslSFk95AKEDEQLLKS94euPvei05phz+Yn3mM8JH4dYlLBXgfs
KLWdAO92AAOPDhSzJRhgz4WSg3XJYJ3LEuA6SsW+PsfGWqnmMtzwa/0pxpGb0PMevbj7WQbX/YB+
Z/DVC9u4jfCo8f4XdJ0ZFh2u0Gabrx+vLvT4bBpvVdn+7iXXJ7djn43SKgxDuH3cIMCxp377/Erm
6QAnUROQ9ESe1LbpBLIrKIhT0JHB+ddCi/5+3OZa08NxSRq+CjYCGFIEHmRGsYDHvT5n5s0xjb9z
ZxI+JR10mgIBpuRfyBd9vydFaMUrXT8LaCOCyQwGMB9jzsJliYJbIx9RTK2pzP6Mu0IAR8ow4qTD
jpVFQF/uI77xaCp2m8TyopxXAlBhnABoGZvCo0HN3i3SpX8+qZFA8GIe0kBD/lL9v14COq/vy+M1
s4QFJdsl3W8GqS/rC8SBmpX03l/FM95TSF9S3EqYCT8sisvFiAKA6bTF1KAvCKX1DtmomSEbWdR8
Jr6WZcwXZCqvOc2juM0iDbbaEncvNTyo10eRWfHyDCMHSgUVV98F9nOgX2Zyk2tBdZX/rYL8Sif2
eQvE8c2vmZmZWiV4tMQq1d/gmHsuyJj7wMnFXCqml4VrRx7j43Ua5nMQzyrWRFtu6QX4taHsHeri
8rG//qJ8iMLFjzlorccKODxTE4F18wH4TZZqGZge1dEcu/DufJHqdhxaaiZmZQ0UlhZZhAcU7sTr
5G+yMJjbW12CoaLdl3CMrbKLk3xtSVx2S3yt5m32yyoJ3VG2/ehedfuZr7HDmEsRSf/5cNHE6+TB
cow/FzdYaVGPY3NL3E+9AWE2PuRpWaag/wjAj55HkJ/znVgPAonz5xyET1KCGc87GQqK1DzxyDUt
5MwlIcLeze8Vq3W/09NiKFETyAf/dwV39YdrVkOoWDYej6k/TES9NVlVmLn/RJqhQjKcmfcl6eE1
GzIqT4kJOjEMf3The80rOUi5chC9dTNCGK4s/vxD8zOJPY7okuYVzElTVlOysVpYdGglN454nDXz
nQrpkVaZA1ntClbgICAtmYM6J15biPU8oS6JnUbnZRSqwpe61eEWaYPVZCKJHJuwDixwTZhnXAko
W5RR28CSXJCpJoCENOcenM+GI4GOsEcBMNFnSdpFwZT+GWrWnR43sBKbi1XNiPRVuYYTUfwbuy+1
8ZxZjFvacGYmdkupyZSXLZjw8wdyqecbi950mcI5NJQ3qvHKYffw7VEbx2vPKEJheM55rCpLG0hf
T0GausZVBEV6X4miWa8MnoQA+/k5q60SqTerdoJbyaIPpR7kIvnmJew2P9s0HQhCDTxKVDxJBS30
Lh+F51PvB8VVdtevoZ0mM/TetwOLFQbxp/Z8sWjF+q6jrZmSnVjPWYG+QADI067+OnJ1ZPp0eSKj
0uFjNZP4XmQAo+rvxbyJpGeV5f6WhwWw+3QLaqr0LzlcDYXDXAnU7HifS0Vi+iC3XXVeyuwcCnsZ
HAtC1nKmEvV20/g+qy2HbeAONY1gD7+TX7zjU9hoglvtFeNMJ5S4UdIRKXWlCKFF9wCYWG/eZ6mi
9iMHvwKQSywscRskb0p98oCROMQifdcLhxkFjzOS0uGNipreL8TSFpi0dDhYIiYQdHAOfohL9mnQ
D3vB34KGwUgN4Fd0LfIRF7yPLAmMNgaE8PiycCmfKJWf1bSVjTDeff5Uve7S90Q1rB0BlsNqjOyt
qJ+5oKC/zjvXzw6w5jx7PfMfeIItacTeAIsHyXhX6RYvPPTcmhpGhXGFvQgGR1m+4X5c07nteF0T
GvE3WGXvDaSqciSDMMhVXfVGwXICy+2lXQ4GXV2DhVXl7e06PAZJhYRtRnWrdmbqESYjLCnziiWA
K4Im8v4qgNpR9UBaStd02FykQ6A5WuG26+ZgETnvK0Rf5/MyAByd+nDosrS78kpo8c/mAPifz+Ep
lr2E/WUull0DQZOd9F2rvExXAxP90j5UmVGWKUO/5ALkvfYXO1IBL2Ys4X47iQmA0vJ34gfFSvo0
z5gf2obJQNYB5J2zQnPeFA1ct8VvhOu5onNN20MEVpVZcbU09Q9ozpc3stRT2fa+fHReWlKGF+Z7
a7y9Q7Gy8HA4KdDSeikhC9uVgtKE73jnqV3C6ndnqn0L0EvKRKr8t4DzgYIpCNxZR/UzVX/kXPt3
ElIpXTcYmNfg1c+6RAKmp3MGOu9/zROqEg9qclwbsCOWWveU13iylxMAMtVSayUaMoUCJn8i/zwo
4M2ThbL2ykvkYFUxQ6qulZy9UDoWx/wByQAU0XlyEuL+Dtbd6AiwMsj5aKRRGicngN/bIEQxBGS5
fAHEj6AZ9nhdgHthtAmVH6qTz4vwWPQzgtLztwnkZj9UZEBX4+eQAtTtDRCRGzqMQOlt3SX5nsut
YAbd8SbXthDlO4JsG0WhZsMA93CSNMEjXFst4FHmJGM9EclmQPSZZwcM51ATXcnYUWLrlK0NmH0A
L1iDmEgj+MMwMIb2lR7Iu8mnfHJ2V9hPwXRneAAJT1DhlpbpRF8HeUBkItk2Ae4IGofvazY9sLd+
uauMBbxmOIh0yAEwEUJ9QRkw8RN+JEetzA7hSaVcGXJ/47JFyR1zMmyoWtXjxc+QjyHXJS7lwuS2
WMrrbsokYNB9X2DCreqZcONglRnQEqfu22qDiGn50j/KchAWks9mSc2f3vRTRhfHjJrRaw4gdD2Q
kl/qYGyICwlxP8vrmQNyvYKbXL9BUmqg+nVelhE1ueTvBJ0iqAGyBMpQl0k6enLGuHtLiL1gVmvd
s9BdNn18VKR2yhN31MOWx3cH3vc8pgZ+cUyw3dWLASdI8bH7HTcLBbVJy/o6IZMClbqYhqeRoePc
5jIzL4A66+Cz5iBCzCY1IicNJJsv4vp6GN6VpqmcoNk5D2Cz3sn06DWwynNktSrImpCgdQ1GciX2
wsFtU4MmBKeBBv2dCnz+8bFZAXxpdQl4V/HQpsLFcxXIIHhL7ZEecJaHEWGEZXSTCyZkKEa1Aznn
mCIEp492afzhVZidols2wO8qSnyNuBtMAgRGVqpklS2o5aleBJCG0NCamAX57DHbzTfZxJrG7GiC
GPsqoZzmIYHAE8r/G7/MDzDGfg1lpx8wjbSvDhjUs/TTiHMDxWRTh9S5eXXP1loR4ymA+8ZlNimH
u/3/5wC6bdffN+mDKvfEXjnTvhGb7tTVNujeuUKbyQ+iYeZW9ihEPdBy5f/C53Mkp9vYzf1QaiRo
/USyEHYkbHTFYuLrNFeIv1MF8FAnUo+mp6BnKpoiUt8C8Gb+yjDtz6qXvDqKi0IRwfTrorhVuXQZ
3O17L7QarLigCohz8XoqqCDl41PAVNlDuQjVsctwg2a2NVc9RRaMKp+oFN0HTUN333VVJfGNvJtt
Zbxl1ySvqH+SQpHFikQg5sWsrKz1/TlTdVznX7mJX65caXKwlvoa+VzFMQPaqKHMaUHuxSTlDUN9
3XS4nLCDde2S+z8olnHV0W+fx+t/8Fke8CcgqR+3APeDIzjpU1o2Awz4NYrUAbqkQRQ5Llx1qOTM
9IU8a6DA5T7csnsoXtuhl2y77t7Kj3bBT/TOfClLLWE0+oGA4BbIXlpbsEvj4S580Hy9YhH0VeAM
36KOIZ1jyGYFgTWDJS/PFgqxSIc/P149LZIzsKRopoT3UeDp31MsvlrWFsdh/vr3Rlp3LpbQXwbV
y+wKIBLJOn8J7Uqu7y0+HOng3RNtcctHfX7ozF7WVlNCMFdS/BqdA+rhxNCcxPf2ibgJKB0Pxg09
CQbuxUxQ6s8JbA55xuxJI/ojf5l1q5EOBoPDB8E/M4r+tb+Qrqzc8RFtIwDg78e0enZJbfdzT16y
2DfVHVbkR+8Q09QUei7iHHJpdi1130DgNJtfPoclM6sK/XOAIvvBe52LQk0yMQlHWn0otlwB0PrX
x0+AuIyG4/dmb/WePUtya/mSJd16SA/qr7VIyeRzvqJKrKJS8brtDKEoJboEACzMS9Tf0iJajrQi
EIpzv7hZObtK9HDayektCIo335VFMcow0PxP/JWXJsKUjMGM+DC5yze+q5lR6M6UarR/C+bQw0l+
/Abo7UiTeby7XWVqFFUWLHOj0620Cz0mBAszmvscLDj3OJog0SqJ0jl4+jDFefY3Oy8WBhsRyx0I
48omhbuLOm20p0hhFBBXMXScmPGDszAB+2WwVTrtYejl5axfAxKMDSidyUQ4Ayx8sXzcz4S0zper
TZLHcYOoD/zoSKx3vR2QjJMOR+EqnaB6zgRBMs+dyCAmUgKxETn+TqMHgBtJEM3Km7vDpCaPzMK8
mYUi8OrqvmDFyygNe+ToLlljOJmkdOMJ3QYA32SzJ2dugrJJLWGl6wLI7hIy+bxy8ezpWMM4AfI3
OXx1eTUm9YjStQcWUDdZwQ4btRciSBi9iVVOoVSsFyb8pha6ystaDPcycbIZCH0/Vcpe1l/4L5ym
g88bqXYod+qMyF8RAhkiLYcTsPuqK/+KAoxwbnZf4R8PDN53kJhMV0VtN4cOE5WsvHvZug/8uZDU
xpdb+ArLeLxnsSDpDLlE3nvdxYG0JBhV1zb4P1obeDZXu03lET5EW38qgrem+HZR8ETOTtL2CY7u
qlcpfQ2yNYE6FW39MKDPwOOOpVT5UaXMCaPlBT745CumGu31uKRJzpNVRrWexvBE9rSBmlxg9Sj8
/Jy3OfFAx3Axdf7SlZiZwIaK4q9W/qdn2vytQJYxQQXZGsgPOpRmla3r3dK2BoIrI67SQn0DzmGJ
shVSJUht4V23KHQJvVRZkUOfzIEVur8xifDW9khAi4t22WQbHMGLsWOg6xI4fcpbWTONbcLlf/MH
ofDMAZyIUg/VLrCU4F9DabOR5kOcEmOKllApX1FRS5Z0cgTXWpzvRFhZsHWUXEHDmPK8NSEFPlJi
je62fAOdh9j+QSz17thBYnMDnREr52/xeYRLiTWO4vcFzwaHDGGlMNTSsfiliyh0m4AWK9eDJN+C
WZNU7uz11I4Xemy4rpEPTyFCUoho9cr0xbzINVKA32q7y1tXiC/HHJXchqrFz1v4fJsbC8bOJElz
mpMKQiVPtE+KjXOve+W52CRPxlPhlVBsNjDj7OF9B434A3HMDHj4AP/jjzvEEDR2nu75osBh9YMs
QaHr7Mb7aZTHtd1BxO7mbXv8N4FSbXa+FrL8eFyupyt78uFoFWOnkWyHzzu1FiOPNAoVYmG4JIdJ
fbAV4zQ+RBKFr9uOOEuy9942YineYUuelXqRwfQzSpY0L2slkswIQewbRYiUMjpAPseZz/K0rosQ
0m0wLi2c/KOXaxtmBsqPfss/nCr2LA2HCNkh8O9mbEMi/kBWr85A8vtxUbdlS+41snf83QMpPhV5
uJagGvi2IZ83aMO4m/9rwjRRz4VFUVy3P5Cp17v8ceqILgVD+WiN164GK74mnA/aYKac+TroZROu
Ea/L5R6me7+thKcPa0qMUfs8oU+faT/EsH5zkCVOI5g2if+Giuh2WI0lzsjZu76QKtO5aMqOxUrV
GSI9hwmA3qUlyQtiedzeupDn+pcYFjPHjnvME5YJCBQdmZuzyEByA7TXmMA3SAXp5POUndCTYrFP
Rk2A2R/fPefvmTon/+1D3x5s6+dznp3iwCtSr6YuhEy90by4T/lX+V3s8Gaa47Q+4k7MwIN0PdBT
gslGc9ZrSsdIYO1Ngh8zES67f17LxLH0MlTktMUr/rXRIOHYOX028pUEiSAhfrNJccCOR3QKNPuT
l1Xsk269PLmm2Oz0T58z4KZS289Y6JrMyrVjDHbgcj6KS6r15EFYAwbK7mP0vZUeFL+4RYhHP6aW
qkW03UJh7izKl7/qhndd+ZK6ffxsUnrlWw1v4fsQR1IyRbM2TB8GXCy4RXtS+/oW2I6Yli+Z3gnI
XtkGXTGOu+G2paSsCekokcrXesYi3i/qVfs3hRtsADVlauj9JhCtG8MvdvcDmYoe8fGP2OdC8tpm
yKt6YRdx8R64B+kroQ9wqIJY0n+bwdwuKTXjPf6eyAh1Fgn3s4sNCp0imWGlGXlQep/OaCfWb6PN
7takVwStvyhtAFSthxZ9lqNn5RMLxM80jo+/EEOPpyHSal736e3mPNdeaPTVI6cNo223r1N0iHwt
Rd99Qcu3AZVp+MNE3hbPwwHEdXPoHMt3+L+G27Rd9tQ2uH26lZYd+wKeYGceUHSE92WGn1eN51vi
MRKApOt4Lo6+LduOknu8VUhMDq1ogh+RNGHZ/Mqsblj9Gi/lgW0ylWPRMoXxqJTa/t0Hd12xkM8m
FBkFqvbgbddBnW/S6ZVTLVGcOwuwarIS6+CZ513cjAa4ewXWUnAWYNeDnhv3f+e7kWOCEnl7E2fA
wOXM5KCxwUeHpP5uoSII3DOclWE2744unYIpgDhnCtAX6xXSrUIZJziGndxQipPuft78uCn2tphf
PIr1bT3rZoCJ+SvANKQSHlQ9muRN6j5wWNin3ac4tITYQXieAqdYJ9MMR9XLael1f8fMzEVwP1FL
F4CySUg0Zv4lvKqvUBc3IeiEZUtmE6E9xyfB2NBAxW43kdjkFryVDeov8rzhd2zMKDpxfBzfo3WP
+eBTV99XeIR7ojR7obecrYWTzxXqsKsr7heriykUwzbrlaZ8ZGzgalQQ3B5DohRR2XqyRhjWf+FU
TSiWS5RVgfbqjBUzJSE2pvefVM2Kz+qzGyxMixH32mJkrHPjI/fHbtUftK4FFrzEALjNoKnxzrhW
rb9CRN9oGeY91Nufk5oZsfN6d2ssU8WQhVGdJkWZCukWGiG8fTclv5cM2nDT+2eZxZVJOJw7CXT4
NZoMu1+sT71RlxUnTR1izA5oEwLGLlpA43BhaQYePuGNlMujHZ3c6d9t2Ns2vYb3oi/fXXEMbzHW
2HHB79obuvNNYuoglmu8vD2mlkqLQSHRqBbSuoN4QgXPtJMtowkESD26xjlUxMEWcB244ah2001b
eQX4p03gXaYQ5bBIDWwQ7jO8o7M5EyncBFTuEueFpE1mE3UgOtQk8FQPn7QCks3JlNNqyJ5V5/f5
bOzqutStUc0hzgX1cvE2vwLvexRkEHX7qIFIap5POWutRr4RGYZ9b4Ka8AA1mS3lKOL5x/SGBgkL
ayV32milBTKAj0+ybseqdELCNxmNCDMS5gozbkZvsHvrECqTCHsiMZS2A7JPYd7qPpqiUU1DrRwn
PMY9WC17OT7FRiY+ZvJS4ypSdwS69ld7HvELfavGPA+gsTNzUPAVJlHhTLHrhetb2a+ClQI7gth6
okOLAdO3mCnpMLY15Bry6u7Vu/oXO0M5WsVCbPSkb+16nes7dXxcZ76DtAsjIDeunXgNdUEKIr9E
Yf6zTJ5VBO8tsEcOwRNpcn/z8/AwMoMYXvqzUtL5aB8V0N/Da8lDrzxIcivJq4h/u3RDHNEk2o/4
Xb+EdE31E472fHP5L8s+jfH0GiL3C6bZ4Ga1dez2jhBHR8ge4HdiJPBXz+0YTecxxYudaVshd5Jx
wFXtbCRjWzZi3gHbcvvI4cYCaBi+zh7PXPCMAPoJKdqlJOELc2WoXb4VTZtYk6dPMCdv9CYciAgN
LMdWU9kUEdiuOGpXLe5R/z/xOFyMB4gYBXJGQBxOycfcngdoajKA2HvGWwdE30XgfVK+wwMQcjB0
h+CaQZpcOTyOLHb/ERj7zpPkOE7IlienH6iFggk9usBO5ZgaK3egInrzy1PUM8uQRshQZY7AhWg/
StBbqpWPKD3ZwlKnqjZa52AA4ZmQyYztdEx5unGujX+avQn2U6xj9vqZgxMfU4s8SzEeKgKY6UyL
XeP4E9ULly0ABxBQr04EAEhVlvc525NZnHUP87XcJn114/KSdrd8BxEmiUdEJrIk0ynY1CfnC+8c
Xsifcx0YhElT5IfEVT/EV3UJ+R3xaF0XNIEN+Chx7+nBu5WJtxhcAeS6J5/TEL40dnxmVgxt+3lC
faO6DH2PKlggHwPxNXqTIq2vyxglG+khA7UYbO3Hh0MuuILa2WuKw1kttI2ZYx8FwDYyX667PXt2
M995zCVekMc8HU9TYzo4zwTdCHZSOUGN4+bcHeYCwMdsO2VDzpuQRbEKZUV2JnUax5Uk8bH0yJpC
H1BrMEFKieGO9hUZMJoHR308Ytx25by9/IK/3ii70q+/cSaolNLYOHjQTXGmwYdjhzrrKvlA3HWc
f9n2JOU6ct121JFtroBQya5BvnnAHxsYct2zekAXENIxrYxl8pibC6LkE8JFdmlkWOAIZvGZrmJy
vqDPcwOV4gEBxsIUd1n2aOaW32NWDqWdgKew9lH/7x1fQ6GEdeBgFRPs9AqpFRAETPybL45S6L7f
jiDqP9tF5tFqV1jps3+9VWbUt364mx4fgumnBxVwaTiw1n9iQ0ftMO5+YrhG+3F6wIOVTtrtZDX2
EAnb4RS1OWX8Yk7Tpue9wOpLezPKybjOHn4+5s6/2Cvo78XtyHCpbVer6A3hrzviwkW2tVDp3tAi
rbAljVJFo/TXeqbZluNhzrWNYcUtQq6GMmxozumBjSlag9IiWTMH80XIohs5pPFEaYi9mWD6T2TY
0zgmw7N6k7zDyHT2GkUYLW9fwsPNKrG5yQLcyf7j2uYBU2FKJYqv5djI6PBg6gLujlsRyGPWWVbX
Cc7xeHXx76c1DFsPzDcBPeohVafAnReWFOUPgFu47zJve17dJm1wwRedBxr8Aclii3/9urVbLzAs
RAxatXYEVqCPlJjifkPHO+MRZiWFIlBc87fboE7q4jDAiSFkwnMyi/cTw/rJBkt17RQy7hcN3sGU
1ZoWFv4gV5Rt9EryS6ORWXzCp19XyMw915uEGVYFuxAenCSG/ihvcZ9iwrNgoD5KYwpjdnIFjSQ6
rUZQ10p+eLglfjRKItfrcMkv5xnnm2sjAzCL4SFIyOkxIq+jMx8cnwU2iXAUqSdkDe3VxnT0ARHi
/wx1FNU3KjfjrLxwtvAca+oAeRl4IEUY+1XuxW/d0GmreF7gIL7Y/rnoOD5/1Y1tJxqw+nzwsxov
AD+xh1RuGlh5EjvravZ1A1gqr/Bes2WC36ndSQYmezOB90wOs11hpa24vuak34kI9jaf3nUxqRDq
1+6yzPazRRtDfzcesa84p+f5ezvXnUpq/i/5QjtvTaFx2STJeic7t/CQtXEZPZIGcUwvRrfajin4
xq72odiZ59MP6IgRaCNu+FAfaYXQWyzNWqkU0yAaXsPjesiVwwKtwI7GNstYvIiS8Gv0xO2yyZN1
mwft7GD6VMAbpaGXxlb+ih9Txe1r3GdcIXnbc8cbS+dS+RYWx9V9TKvv8QEqqV9wNf6bSNdDIXju
7DRAJlR5tPqbOEszcsHwkCzFfqE61LlblGWv9Dm3jLSrur1ulazZbwK4FCCsnGTnWugDOUV9TvS9
DlXUfJRL1NIHzFdof2dxi6uLlkLpUjzR0z36TMfu+PF+bvNMKlm07ZH6jkvqIRDKexv8UucekSMy
wSqwEV2vWtQYlGpbco5+jxQ8oXdo8BXLklSPx57ZyXN+m/5CiM9fAuR8rdUR4Y7LQQdV8ClfXNqW
d+rZtLt7iOSF3VLEHjmTTB4HFqKL8XeIgu+UriI7P3ImjCKVvl0Rzajg4N0i0uM8N2e7HvSlNxoJ
6vZqngekWj8giEFkGms6ylvhILAceHUpCW4s7009Vue0U6zodcDHSJI688l9aOGOWQY+feezb+Yy
1zjWxCcBzCUus7aLUfhUL1irgjSd+74Z++K5y3kS4vraWd1RXFiGH41MWkmnlda+KUMuKTvxR1GP
2VGtIAUnh07x1vU4Tsk6djrsvTokWt6mdXh32RFxlMvCIHzs7Lbmzomer3h4PRY3CZrwSufMd09H
Fyk+BH3s/9RLzNNW/AWYe8YqnLxNTjPU3Rwlk8C/2XgE43bt7YSOy4gKM+OLgiiExLOnZTwv67Gh
obFMSNVVvH9dJCTSCHK4crhiTmRss39S6HtanGaygCmCeRE7m3DHcBCv0hHOE4+E+FT7aQNSrlQj
4kIW4fFnQ3eWg7RBZkvFAKybwTNAXXYJ4Sbey99Qb+bHg/Btl6Yj9PaAPdaBxN7Lfl7wBplcWycI
lhGZjJc3cfwc5eVuQjG45N0b+rkKVEyHXlfeZuIkJVdyja6X6tjlgIgY+E4hpgAv5TB+hCKqIziQ
M5yHz91nwHur3cWYOBkdezDGEaDwLA+fiFwJhyLMY5gen5MPcLvHwgsrHYNuvYB0mKfjvs7odkVj
xhOf1i7AJhLGqCRSh4VUY5xJAIC5MxIhWRy+Le+nXIl2snHj89Hu3TJsiEhYTvLcinroGhY8GuVf
4uc+SlldL3QuDa5sgSWwtSOQucYgp/XCYdTE4fvXysM5FTXSgeHt/Jj1akqmxsJtQpBGDU4/Ke3N
nfWTXARoI/czAYVxKy8gI/4ph+zKO8aIag9AJaOBjlw5H0CL/Z6PLUT2OCNZQPUowCMzdrgS0Ms7
9WzpIV0jh0XpMyn9vl6O5r5d4T15+XqxR2eW7V2YR49Xv4oaNH+v71QfNCHTkWPaQhtsDlh9DgEE
IZXM4dEx2AsRNmmQUEzQf79+64BlWSVZF6x8tyjjq4VHSjTGToE269TUzwdhR1Sv3TygWiMU9Nce
eAh6/7PXTS7Tjyor+5lHo/rnYpfvb7mg8PoMlWOrXJ2Wn315iG+h0LtEeSImyqSPbof1tLGnY6NO
V23zxwidCTvOY2v8Pf8xmT/v0gBSI1v1iO1jjgXDWx7n9C3QJmf2m6zXfaNVATg1rJ3Dz0t8x5LY
8Jwx6KJmMWFl7s9EI2kc7PJ0jObeyDG2cg2U1anvyoCU4NB/qKylyFY4U7CCwe2SpCW/R0iCBLXZ
tlDNEswhYFWvsKRFpw+N6031Gf/Thb54ss0ZRkUn/yhkEffWpT+h2Y0aQcP8t3TY2/ALA/icTbos
g7uR4IEiqAtzWG0qA7Xtx+nryBRtXVj4bRlXhoY0sUZJBXHSF4IzeoIbDee2DxKIfDvFTUrxwaY4
vTnF4hLUrmbXDoKz/6MpK1QtTz06vWO/QiAIEUtE+P+5mciba5fOpnbuHf7/yxvItY4DB64Bz+oE
EzZAwLGiUbn6O4c69ySQcyUbsFPnnD34ieb9SHil9uxjXKf9jYNb11B+8SwOPhiesBEGqCfrAOtu
BuK/tL9N/uepZQ07kmwdyhxwc0HmzJlDPxqNhjGabClrVvMyA5v97ohlVQNobpFNwgLtBQ5pUdql
IW4P0Y5JqsBedffPrZBlT8+RJQs34UhYjOeoNaF6csCq4naUp7Ylmo9h0vS/CBV7rKc446OOTun6
1Wk/imYFcoIkQWw8ysvbNo9y5eba9qNmqGTxt8nt3p/COFQ2ccgrDaXAq6iIkZTwWOhGloR18nd+
YJyRFHJR6WBGS1GlL44x/Mu+DQCcd4RXbmIU98VQYj/qd9xlBPHUsAKPb/ZvAqgpviSwOJXeMBHi
3KOKwFkGOBnLL08y8duA3S/Z1a7eTyTdhz98ce5cSS8FdV6s9fTDatKQ//1BrBdI3iV2JpDkcB2t
lo6Lq9kBz9NPiqG8BIAnX1YRihNeLNuaKv+fkSZRYjs8CQycZm+iMQ4BxsEEOeFueWmroFDeOMXQ
+GqWqik0efdgBTl3er7QJaiUp/gH1G8yHhXUnR+9LHqPoSfP+jITzY6ALs7VRroukLkMktbOfSqB
hsBxakGM67VlK9tsHItykHdzqD4kww59FuNdUj7X3VnpzKVdSLqFE6gy8Fj0pVCoZ3f+DI55kWfS
HQDHN92ITn15kueekhJraJFRlISpe0sNuQuKeMbWk0BOd3SOH92AG2QjZTAmAqNs9EvHUavQfr73
FQpBj9iDYwonaoF+1WEbe3Lu+fAO+3f+A6A/lRkk1kK+N/GVRv7IvlABSW72T54pQCKV4abg3y1c
Re+hMpVQYM7h5Smmd9QtRz/4/0Np3L/2XZ0s6iS4gvIgpro+G7VKbEmcW+v9QwQA+oCYO4ufvEmB
kcOEt+74gTk0qvuIGyAyyZIPHBD417dx/tA1YQ5thbv4gIe7QryGeIr37/B1ppsFCnHk0bqc2JMR
EP1v3TMYO0WgzLSi3q5YcZHOq95chgLZU5TkqNKTBOZLDanrGd1Deo4ZuCA65KFbdbsf3Y0ZMnjY
EO5aeZZAt5Bko+gqwxGWhCi17hXeRJSaEBPT7dZ5q+B3J+pHfCPXpGoqg1sthu1JYbrkXV1qrAVq
cldReYWLAxnTOJ63jZXj6/e2g2LF0b1uNRTyZlSp9Ddq4yceQK7ao2nwcG8HQYmCVx41YYhH8EJT
IJiGVIVxyZv5lMAEHZAfJGHyVKfaLQ2Omyw6D7koiuZYTgBDtrKFczUJyZNJ7zSTepTYSYvSikYY
x1SKBndd98mx3msjCmNfK7vFDc2i6+yixQVE3Ezc/7pPXCY4c8hS6g7ywe32yDMUVJXnyZ+1MgD1
abnYxOCsmKh+mBdQtJ6f7IadjE6soKh23plGLwR42JqB2UDW6uGaGTTAvTW78V08/kMDKnaOhyFv
lKA0q7Xn85J25fs4Dgs614H9v40P04vLBymXnGSmeDmNqRpgma9rF89Ec4ZiE6SyljewX/5FbUBz
S3ZqqOILgImIDkwsj9f/m0cZkYPXOzXIn0IHXDhrJ5Iwi8XM0QfvQuXibC553qDA/+9kr7Tz7pGS
7UsGWeji/W3za0haTsrSnsSLh9zMwXLRlM/DHQmuZlWtiCW/8nlDGLxSGk7ggtSBmwDLKmCnLI/T
DKzXlAWUH4+gZYOPOpguQ5GYkm0STXiL5PSHzclx8BorWc8JFmhK/xliMz+Am5jVS8SB7c16YPuf
uOuQodHKc/WVG2HxRPZcwgk/douGdPm1fpKUjphfY9ps5mvkmJeQOiSFeg36D4rygKlfZo37hpdv
4zcwp9Pp3PE65yXB9oGSf7zOtcEBuzVuvIayIwMVj3y0clBNKWs1VDWDbaSBuMvEyuqN3UTMs1m+
ZXTLFu0+jBeTet3dRzAFW720B2hCiyNxC9pYDO+Ur/YJckFH6+tDPBNKs20OotLW+U5sQKPBl7BC
Mqk/Ok3TN6dxHSGVL47RuU5TwalYQ28Ond9bAPwoPA0dcLVDBp4uTruvcdziXHvsPjeYAtYSrLdc
5eH1dveRoETCfn1Kt8Ko7Me7KKcuLNlTFwcBoZ9xVJQ3HpjF+l8Yo9haPTIDp07hWyvu8NFuVtgB
k51MafU0nGpyvgHCIUHvq0k8hG0lKH6xlZqBB+xXSw7Cl+zAXSBd8AFWqpQ6KoTHloqwvvR+k+/c
cvScEmvlupHVeopuQ8eV5AHzHuupEa4uH9ZzlSNcCaiBEqPrnNfrtyY+B1vCYl2FMemlqivNUfcx
WLx6MLJDcio6T/TJwWqW0sWrCFNe9J9Q1TXbokWm7Laf+nkFHZ3Bnl78zqm8stq9gCOol8SMxMyN
6psBLRSgWoQBpBymp24tF7uK7kY+0epFCt2KnDL68C8s44KXe4tWGqduVz49OXprp3t6mPsTpDV9
KPgRVHQlWBN/Pc1W9UXs5bdCOoEBlCgxSdoaedGASObvGhrtvQZqK4x7+FQ4A/ibwxhBPdtIVs45
QM7ltYQ4YTDcSiH5EX2r/vgEzrqBxmmUzdEx8ejb/6diUHsPoJnyJBlKVO7qH40Y1wIYi1mIk2sB
I1yqkEcztjaH0GRFossxAW9wDKq5GUNAWkgwK+FQhic534aKlgLgll9tTiwm/z+CTmvXIE/mO68T
v1uC5ylnVzo0YaksyQoM0xgMi8PV+iwCUeruyFAuxntOBm/jiPKbm3Zz1XtLCmSbyKGjv5rO5NUk
IiWmmp5c3Ka1GqDaonenTgxuDHxb4l9QYzqhpBHaE65gUMUlT9vpJzLvpWZNadV96zzQLEQ7x1s+
KPQR3Q974CfDfKX8FGERoz8PBZ9d9OKAWAyXPow6EeJeg13LG37L6I6yayUhAgwb13AMF3SPt5w/
eSplAGMuhI6kweErp1czv68Z+1kfMLoKbS8v2dedPaE+aV1DZxb56D2ZxQj8mu/ByFJ5rzEWMxgV
KxHO7XFScUe+YhBcAyL6jJpQdzAEsvOYNd3crflLEgXqbii5hiMgxEsxhF3AmiNTLLpIx+K8tHDP
Vw9kOSfSQcc45KJn/oK3zB+oX/Mkm/Pvau6ezCo6nnJtQSNWupepYLudYCFmU8Q317ak3o+n63KU
ATVcsid1rqublme3SZWS+RbJCc5kMBfjXWAC1cxALGgx33GVmHOrZpEsmI9XmF9gGyxfAKlvmK5Z
GSRla0GrHFuZ4D3U1dTczLl9z5QktPI5ikeGhXfOC5roxjq4ZTu6VoZjLHw3dA0QZ83CJd5ij+/q
ska5E4vYPz18ivdWyE3npvIUImk/oaDNM/h/GniNVjdy1kg8YXdCCB/pKDHDS5vuYKXLKJLE9AN/
eYpHWt0+1Y/XFOe29HJK00bAiH03agiu9vuxrh/4gRIiUs16DGYg+pRkpVD+eyyKQchzjVinsX76
fLjnaqw8Lvn2++jkIDhtz2q5ec2Ef8py5aQzFU1IG8K9u4xXdCjyhH+OLjSzIiToS27N8vGwSMHY
3HQw5KmYigiiGPQbp2mlGFa2M3sAwF6NrYNVNRKG3EqogRCxrpgbqjuAu1/sHdjbm5lewvwMon+v
wyJtf1rZm1d8FHqaWo6vWzizvTbInwhOsDhv6RGr679kPX86IllrZzXvvCGB3XuIHFg5qXdlo5I2
tXJcWVfBOdBm6Z3VqPI3C5z3C/bTHm+bXPuwEywq7YvfNnLXLtjZA/ltJ2tD1wAIM+JnKw9vnygB
wzrhe7N2vhZjSuCvEVb9RItBWKtRNDzoayoFZlfelUxypp1VHToZZ17A6S/sBfFtOp0Q8jzs9BWN
nPmbxcouXvd5RyfFRLHFFr9E/ya7DTU0+U2nMNyI80WPVNU3SCsAdQ6rQ5hOZS9jDsp8lpXPXCO6
lrksCxkl7WF93tY7uGuVuWy8Hq7IEyLg6MP/3tQWbOyCeK4PzEUvtl2P2mOSa6F+j0p1eaIlCGfL
Nj4b4UYty3C22P5M0jeZto1Hq0MdU2c1LaCia2s9OXbdNJErVMCeyge9DmqSOH70wfxmQxCfFeEe
DxefpUfV8jC6DgxH4RIVq4WN0a/9LEWKdT/BTVEVWQO+GmjNIx3Mq6BdeBiw1/a+3LL1873TSlpJ
rewuEJ1I3EerJ/EQzvanesmXXKlpaUErx3rOEoWdH9h0eyKcqDCgRjFBV2Mjo8IE+gpqxpLwvhvn
OLM8gIucK0Cww6rRL8Y2a0KBrYwoGBSRCpd/eEmHyMgIOzhQA82nP1xus1W5UTJM4RdEKc7gfQMK
hkz1duy25OwJPMQVLdeFzQ86puYsGk3finWOp+aYxMlRRQY186+OsSTMpflXQbUjA/12J+zgdMiD
hLgVThIwBX02ziSASfrcKlYtyY+9nBSEWd4mMZ9DpaxVTvEnYLT//mzRtkkxrKfG9OSQLgcFw5cl
4K20J3VaoEbR2r0lJFlvC4N12JdB8W4lvwjptv/ngUa6Nw/wTDCPXyUUP1HzZ3t3Yydo+Vl5Q02u
b5gZntCC2O/dElRqTXTtV5qEir9Kier8C6HowDXSCL9pIy7t0aSsZhwpI5qV48E1ruu5OxQGIF22
wuQOIzO+iLdekzYrpevrJ1yooFvOsdthJxfJQCQ8/J46hMloyOcOBkDsk9bKaJmdU2bqVTrqjzy+
B60w8++VWdCE6Gs3TPk8erqiORORV+sRDIs+w6xafNEwdf3vasAEYtYfEj8wgCZjakKvqOPUBk0i
XWCYgvmo0Zosi1NlirfHLuBmsKGlIoZaBl6JdhqmY8iB3HFn/Yb4dweTTei5qGmexBM/Hi9l8p6o
RSGizwl7qpYWZkvoN1q3gajgbbgpgJLc59VkoMlfv1v1ThbeIpuyxnHMzG0b/waBngx49l8Mtwwt
TI2nvcTEJ2UAnl7KfFK4sgrS5u17FhB7M4pT2r5Sksf7kMF77muzbEVkJSqkrTnCU47pU2lUgh7v
y8uHWtO7+uVYfwRPytJ8J2rDfPxxgP1JYAp9BkRiFBMzhSLbhZD2gYS+sxaSQb8VfN5UP3hHZS7S
GgISFli+QU+y9z44jks/fz+nApku/2YrLDk4sxQ7XZ2vGKyCcmFIuCVB0GK3laK/mUyDonLq6scR
0PMVkoS8aDtq5v1AX6uuKzBt/2AIwosXl62qn0b5hvbK+tJXhr1aXVTWaqsjN3lGyHdF6VDstLT/
yupQBZNTW8T3eI331DwljcImONiXyhV2zxJ1JVKPs1vbR2zqHAyJZQUWgHXL1E6HMOzhiOJCtSl7
buNjFQysVhHe1504bXhLXqOfS/Zs/jOwczOh1c4xKUkMFcpomAEqvFpk6s+3KePsbepKmSsCp6t4
ImjrlHiA4OEp8oqDFhIwfODUPHsFBcdH6hwFqb3LmUXhZyT2DoL0bCBArzG65HmDrNKlK6PWUQRQ
kETQY8X/skWs8ynzP9AFPb7+0iFvBx9lENJi2jVm6AABBg4Y9lT+k0SP92HseeqeTNBOny7ouRsj
O9Z/fBWcrsyRWu5pIritFdlI73pbvbnuo3WewnQNrrwENtNVOXGYgP0Au+EOluLO+XoZ5G8R8kw0
Zs73BB0kHrrh7az2woyxqWFcoFkv/3urj4XnayLyCdWRqICWYtsNSrmmb+Yfqoaz429hfk2KHxPw
X2Lw1Xsz7d778PvMdyIvnFPkp+LjykNdVb32zjdx2e25JNiYWZqa3UzMGwrkYaU+gSxv3v68f8v+
2GhMsPttzFu/oDNAJCFE6TggiPz1uVyOMFT3EGT77rLJXkE8FqKCUJ2bh7Hf38j/irx4NTiSB1/w
yTgnG4EUHrqpDUiQzmZZk/6c6ED080Pi2wqGwibod8AZI4jSbFkkz41W9a17GucWCvFT/m2wPzNg
nSzh2SWBN/iQ9iRtaE782mPGWrAmG9JhK+8AMZR+s0UfM4Th5rxLkV3T40wt0ijQ7VxG+jtRH2QX
DTTPu1UCMbxN2ANeGzpsOUbJkOYFqcva50JdHdRqDMOycNggE7ygDtwd/vcYJLX1M278Ax1+m6tB
NmsQ6/3a2Fokp5xfYa6LuEjiV8aCnQyoLmeouo95oUon1frDhL6RjDqRxyzIzFQun7FAzhttgloT
B8RqyyImw5D5Bp2VXOQNszgZ3bdR0pTM8BtM5KEd/uLQBk1RA0WInj0Eg/Y2Av1FGnZPHbE9asxt
I99LTynxefDq99SYqlEFjcXoVUP/RtKHmT3xxZ1Z6j0ZaepVtBzElbtDW5yJZ8g+tFmU8Bvcl7l1
lJ+Dn5hf56B4fSoPSOlYW6tmKwxn36C2QLyD3kTDjNzV6JWTvxiLbB8KL7X9jROhWSkNt6uTaSoE
c2pBYy12XT/P62OOZ34ygxPsEAjW9tfVlxOJUnNuNWPiiNj4nIN1utZBzX5IU0hUL601iVOkY2Lk
pWXGGzgMBwAMVuBjpqckMYfsZFdzC8wWeeBIPQQkxAburYiW8SrIoroHhwmCuiDxWKScbl0YH1Cf
axRLru9o/Nr8AvrgkDM9IvT3dEisnbonuggxtfjWYzT238hUVBz2txG/eA3m8Z38Ds2e7s4kOzh/
XnilAMwKeHGGdNvYA4uWGyhMWL1cBBCn9VXSlz2eCwV6gNPMRl8p19Hv33rNVhH4RD9I+bgMBxKx
4teHwLupgMr/q8B4YkIEg3ARTNCN8WBUW18i+s3fCnHdSVquKV36TAtkvxsjz8gjuDB/uTzjmLTw
yJrPOMOmyLe2+rZxEDOJcGgUBhoIvWrv/Bnqocg3IBSEvhJ2jA78+Qqiao75cXto785VEK2LPNfJ
uHMNGGxq1nhp2KGE2reRmFzmJzXmAz3mFiiKCVJTRvNOQCw8HD/DOasWmM2tcs+G0o5mORMQKPLz
ToN7hv++yXQkJ21j++GyzY/I5oRC7U4LtQyTop8vKen0Omnhx6jnjDsLaDzfO7FpuPJpjxFoRxl9
30xqmjKTUg85j70mWotp0inYnQqktDwV0GUx87zouRtIVILf2j4FIv/nlOh7am4QteqYaS4+EYjT
BlF+0MW6K17QklVyxhvqRltv5ga4tKx7F0tlrU+txKiVd8tzfw5r/B5r3vOQZOwTRgFlTZqBOTQ7
/CUKts7DrZ9xTKA5D0YgeZeDXw0rcM8IgikzNTHM90GFtcQRtj71NXl1h5wf2tARyWOw+cD+a/9n
YHYvOgHcestYTy8YKgr9aTzDv05vVeIZh6hsryBaSTcskDqDvaA30ICPQrk6ZExoKibcAa74uPt5
XCrY0/hm468bhdVdlkTjzSAPcqEBrxK0/R4lgqpqYfg56t0B+CojJnxNEKjQWgio/QRruaI/QwIO
wRSNDUReajhpVwJSWLq71rcj9+UBFrUoHvwbhgNiqvJv1CmR4ht/s1p5/OQrD0Ga1IIx5Jw18ll4
71l1veAXok3LkopEakZcV5RfcWHV68VayDhiclmZC3ZLMyC2FlMrGtR5VOjJyTCn2UzLBe/le6n/
wIRBR83x3L36U1g+j7500O309RoJ0WwO5nmpf5jbaB+un89DW10UBui5RUCoWc2W90za9RkMAIwg
HbfOjMW8toLpy4ByzoEGaFZVeIVDgjtDaeyEhgR4aNjvWG7jByXHcqhipj5wu86iuxcVVDmvPSvf
Ykde5IXfAdRu9cVNP/q6luSDMRyk9uUWC7iG+jlcxoa3KUckPEPSVuObD7tmCqSQNIQdMXtAxHRZ
McVltZwtjZ9gsacXUgqDT99GcrP3BA7SglA/j7t1K6Ph9wfbD288Xl4RNgq83JT10B0JKusrVRb+
Xf7fc0+eklRGIb1+1BswP45dlgn7mgeSG+gFl/5HEg4HvpUbDcnm+dkHP3oTwvobdTJxF8YpHAhp
ynhE7+zbwIZE4l/Pu6s8M4SAJscKNksDp5OyOlO3GfwwQEfC/MzHVzu0luThQ93Adg3TxFAFcgHL
Q1n1gDlJW9mw30Go89yDIXm81Pd07riMUnKhOdpg5nackaybj1WMLOSQYK6yqRSiOg+sLtdRbDcL
mNzdK4R6xRJfS3mjFL9u6b6x4TBV4llR/y3tUdWuOlRR+kFHlQxIj+T3djaSN3k6pzUaKrqt3V2r
+z5ygYjbv4S49kUGje0rkHVaHCRqVYsPifGZJxUS038e00jxO7leuDaqlxaL2MZYHV8mhHu/nXyy
qpnEOgeIjmH9yMK9tPjbYg4N84tdqm2FhjGy3MJnsZpQpcY6Egh99OdXYmhdlk1Itrz/FSkUTOka
iq4KNBR2b1DyMN/GYv64wgkfU7qLJgqqdhFwnAK3TF/l+2kvvPiBVR67SkyAZE43qSyscKt9urGx
DMdyBb3+umrXkg9TiXuQkGUb4JJScuvtfnLNkK5aPAVKPSHbXxSJTY6UusilQbPSTnofEDK+xV/2
6uuHIOleYPCk4r3MgenuTHCD+kOKCrwDCP5kMKIZZ+xnc61e7oydY+DwLxKgMaw79vAXnfLjW4GA
ZPSw0uYS4cpYxDXI0HqYVKVzkGJoZ2jpkhQnKfQ47KAtU0f2d9K/jwyEGoIx1ijY5xydWow4mfYM
QLIuTzP/zIz0RmIAP4L550V4EvPYhobBqtTZeu9hU4nFY/9vCiYoUJTGeyodMftJMSlaE//mIGNC
rHU16CDOiZKtaLVLEAL7POKO6pkaoEWFfcDi6rpTCi5Qyr9NVA0/MYuUbqwqtHQLzBZrU+oexIR/
VFRomGdpiiOstIDLQ0zdGzeg5UGwskTB6ZhOjvVK5pG7FLEiXwZb7MQm5eelDj2ZwIwzdyglOupW
/jXcPB+bKBnrgHU1u2/1VDEfHC+aK50tY1xIKQt/q7DTMtPCUIJ6xq2A+sSGhuKyoJ169d7pmung
Y6juzCMCv0r2QYUPXpGEpUPYbR6y37EIs4hIphNB1hr+SQmPJ1tCLXWRMsruql81y/doawne8KSX
+et5zszgJaDXMZsO/bimwcociG38lKWPxX5wok+TNu9mJCOPI2Ixvkrmm4k7TEDymSfg7iOhqaQL
gLPFxWgt2tQVWUvZ6OprIk5YY06Q6MEL5xS8pYFC03AAAXnj0mBA2EpYJPCc7OiiGSXN3t85Ga5W
J6SvZ2t/N6ppBlkMHpk9zgBG8dlcvUAsIo8FU/EGCIktuxhQNdV1clciHSjfy/sDB9U8eOk9pK7J
X3cVmtCeHP9Mp70MTWyTupyG+xxVRUdm98lTJjZx2j0oseaOAJE/O/H6ZUQ5CepGQlaZq9yM+7Xw
u3rxAqx3VRmLbeO+2mLkZybkoL2/LpP3J9QB7sVNYx8uCLYsXtV2rm/cLIKm6AjDX8yIVN0LeBUl
98oCwTlFRxrXIoLqz9SFbdwzNet7OKyCA95Wlpysqt2wXSH681fxVQ0b4+rbP02JxzaZsgZTtucO
0vxtUxnH/BIReEtJOl1TZfOqk7CWhgYZmn+ZjpEuEY/37Bp7mgsodgReuUaCACQeIxKNExO/yg20
H1dAz4DTNp4FkP1hUg5IEhViF2+yrG0vtQaPRJUbeo+ihiNOkEUQ4Mxf9lN+zMTldPhOw/YHVldN
eE5/4zCvUu04e9Joe7If/SgR8mkcSgsCdUyTbWQkiBjuyQ2Wjo5fXFR0vKJw6vnXth2aPNW9AskI
KQT6P1GiaVc6Q1JqqwfgvceLFT7Cr/fRE/X3Lluu0vPSO+M88raQkAUWOHniFP8kka38G4UvUJRM
oJL1eSiRRYnfHP96Ci+tiOBSO4yhoYE/9DodyNz5pWfHwiY8goC/MY4FbkkJOEw+6TYCbP+HbFyj
Z0iEmenpw+MnoHIsyvFJUK+7rOS2ceTGZNpvWaePhcHcbQLZxSjiEKcIoGVPRaG9ta+WoT8QHjhj
PklQbbRAojb5iKeja6/2wYDLYqk0vRMZh/b02P+MfdsIrdoM/qm8ZUSHrfwrPWNuFadZWeIqGqPn
7uiGfmj7rk3fMssCxmD4Kdu8Y1EWKWk+cOGeO2G+9PQipWpg2CaR8Z3igef430GYyGm/J0rYfye4
JNEg5jf7BuvhyREIeryH5g+aqmYWbXcH8ob9h2bIZlhr1FpQw6d/TGFKrNXe7OPl9vjPsKXD9kDK
yWJwPKtyuTELLqBgDC1eJnZwjSY88RMkzvPlUnbQeVuRtMUCagIo6SgTmnVMxWd0M2svQrleZQGR
mEGYPajDuU6xwUmVPml2uKduF5GkNjX6K8QNAhdlzZf6oKMlQ8Nj4xQexkhoJPjN4n7ElMO10DGd
8xkCx2rnIv0KgswfflmkULdMErFnr9z/gAoKTdWuSSljIHg5lbhGYnUGfJMVrRUV+OTPqD6/IqUt
bCoXxhiD6/JgOoHpvRzWoUoojDU7fEzGoA6f8BoiD/MhjbLJElwzPY3q35QVdjUBPLgNKta73R2l
RZBQbQd8G8SonGL0TwYYver45WWMzA+mlzaGahvxb0utCDXMU7Dk4DApb+Uaw3h2C+8hqiLYHV8F
HQCgXfaWJIIpjHPrZ34UjPpLDreF7I7d6gZgj1NqNadRWWlHBKKZ2jS3NQCeOAT6IVlT4zZVI3C0
nGzsOgK5khHr002enpG4rcvLMJVodAglckq37/kwBhcWTJfVljFo2l3qatV25R6R+QF+N3Jo3XKe
jNRyRiGB6BhC04IRbhwKodadewJLm4WVprfkg0BLQL5ArpIsMP9cIOZuqQXkqcQYup7RHxwrBjgC
7CS2HXvr56rOV1RQ0QStpaQrnfqygCy0hFeSmBCuLvxh6RAvnQoYFW2MRQ5LP/ZuHq+hhQxDAlIV
4Nx1UjM+NhVUCTMpo2NTE2IyPNCmr9ru24HrII6h8tvnU+q9WK3PovV6fW1zEHOZzLbqVJGrh6jB
syJJ8hTiiKW1EBb7yNdE2q20UYHzlCKNDZ/u1KsmJKpHyXJCqelT1ic3tRRsHrG0krmlPvRjYZxs
u58jA9Ib6xS+tIjMgKS1bATRe/JEHOesfsSCoPZ/Xi2U/GBeKqRQ/mrQ+e6k6N2OceWdq/c6SAO6
j5W2mX6m+6uISBZsZfWiqcbZDRgUj3MKTbhpkwqHXdjRynqvM3r/pOhDLORbr+Rqc1UP6gOq0W1V
VnDj+LBS3DE9e383EA2dWuGu/AcpOz6OXYKFSSD+op6Dpn48exGAtXtF56JP0OxHs/vGXJAsgydz
7XtPfylBEJ7xlSyUt2wyZeQtmYA4yIqLXOP4PtS1eeUfDNAQOlaxJVWCna5PongiKDJXVwv7T5Pt
YZgGF9WBpLEgxrEz+3w7yRxYEsZrQhgzo4mskiljrVXGsxZB/W3Che4mr+5nS/6h826D1OxryP/H
R+lpossnq8qPExxY0LNF6agxkpOXb7vT1ex5+HSkjik8BG74vQAMbLydgoMUZh/wGWktCcFjQD0A
JQaeRBgslmY9myI++vMnQXS+296nTTaHq+Tzmmt4J25A7nHfY9leAfcf0YVCpF/A8EVL6G1pfo0y
16+eZBhfJ9NCBuzwas0TAgbVBFtOGG/kcaeDPOuPveCjaFRNHR7Gc4rZLYWvqoBy40hNcJj8JiPS
tuAoTW/abA2+7V5V2+L/Hn67KwpqrZZOsJGWxvxwELdfF+SuUpsROzuWVQ01KNxtwupjSvvjYcdK
JLh4sQGeufMmpGrCFFmyRrfcQBEXFPWmotCVJksGRCZ82fSsbQ8M0t4naxwAohSwF/razi0b6OEF
SY5fDxyqJ3yq2zlBE3X4/mDmeW1WPAuyUbpokrjDu/nR/EncGHyAaRY0/ZEi2XF7QQ4bH1LvnXqy
sgqbs+gKy/kplOX/BYD8FXaQWYMTp6geYC5J+3sg6QFST29uF5ZQLLTqt/cmpcIKwrhXL9+j6SuO
jw7j6f/jsAKCy7+eYA9jqPsLrw5J6yIsSNzbWBfMGY+7C+5ZdTzdtfNquqaI7Q9VKgoZjivjnuP2
O44VoxGYKgixGziyoxcXrtI30tCk5ktZORSd490hK7ZL72S7Ce4RlyqdXqRqH5/zPaABYMtH3mpD
O82O5j3URrfptW1WW6aVUyVmosbv1gAn8CqQLdzx5U7UBvwVotEVDYQ1BZIU2yvwyVxjll7anrRL
YMkhJmX4MH/zyk9Lnn5ZMsp6SbDYro7dUujBAhLR5Qo7FY6WOLDJ5AoQfr983srN72NX2wtubzdU
RyxEUFFaNs1wJ4ipjM/2Jo+sWtkD7DTlRSut3CqCUH4zgGyFDqWbk4Mjo2RMztDvPJv2huA8fhaI
N1B8Chm7EZKiRoY41RlFof0BSZP241pC0u6O1/NYNuW0ph8IfhraaH5OGX/0R8Y5Hcnj9SSDtaH7
d9rjT5mZPEIr0N5FeeCmx7oHfcA8J1nvnfhcA9bwu1dfgP18dOyQqO0W4qTB6gs8H1Z4aydCE0Fi
CUycZml8tHXKQ0TTKZDy1ch+aAqY9RKrBR05RB0OKLFA9R+D6Ru+x684oXlhiw7UT0F8oZ37Opk8
BCJrcd9d4J11HNDuQSo2X23XN7iNGLpFFsXzru+hyxk+YsAzmsTma2QccqEfPEbsrZ1SM1uNLl/X
GtzjERWrmpH+Uk0+6yk9QTejxnF9PjIwFe6c/NGVQBNpQES1Xe7iNxqAj8lEHE2SHfAu+CQAHs5+
a2NKjFs1ajIE1Dm/9XTdC3gfiUDZVUi0KQ6CT6aSLEnq1hR15ts22um14AexPnaL+4mT7+osodv1
gw+uSiYEwvcBfuG5t97B8uoM5bWzaAkwZO7bBVVuL5G0/QRHqltfXYqup1gbxx5DGAKlHSwjRXFt
tUIYiS7p9Aeclk+hWh+hJKHxoxGx6byL1n+yg3CtACF/nSW1SvN9TKGyxzEL4ZUCSL0SJhJrSFIK
/c/ntUKq7nbqh19+WipS6RtoQJxUpNUbeYtTTCu2rLyZTyOT3fE/p7cF6m+J8iLgIU7s1mca7P9g
mq2ZbkuFOUvNfahpvVPKk2gL02phhrGmxSX861zHj0S2wErw4ml1vXH/W8SeiJM6mTig3NUvNemo
cMnVKW6rePHjZM2EaMehYFlp6AG3Sx8cdD4wJe/IFLgibLGiedQAc+LYo4SPuwcpWB7t2W1TXQB9
rqyKhHzaQCvFo3WtbaZLIgytQ7VI61DXH+06nH+T9ABFtUf7NMHG2puiq26Lg3w7zJWNnKDoPww9
WOUuhQtsxUOV/Rvlo0wgmUfKdmnBlwMR9UL9gtRP7DjlJ3nkKWIJYTrWyLeAlHz0/FMm9/5TgFEU
5UxDz6andh9s0bL/TeHmsSijVZ+Fm6Lb0iimPrk+JmMLDasxBolke3RbJEJRlUO36EIC3FGeN08l
PGIuSz0jHDuOHKNv/YYwcwcVONRrVcHXCK+BpxNlKSUEbCIk3hl4EJXoyzPzFP4zjC9epe6d5ElS
1GaM9XXkmjUmzBcfFO7yoWxXMWB61vrMafg5RfmdjcFq8Zf5zmwXtd/GdbrqkFIFgcsATozjNldt
wG8h8BRha6VExwjocWmP97ARgUOh6pyeFxmFn3C7cOHMJuIl+1LCHSdL4iwODeAp1s82/3ozlsYm
yS/ABR8Wq7RP4hgJpcMUjeNm+ZNxtPqBkJv12BCsyTmLRg65lQojHh2xWXyt/g1wSDs7F8VC7xQR
Vl8W1b29lvbhiq0h3IAJNvKJlkxpaIXkp48PbzMBbnup3pN4jUyXthCuUldP7OhwqIHuPq46YkHi
0gHfdVq1sjpLoi7IxWzNqIHEOJf50vdx+V4H4CFkEwpnAYVgis298qZPQvf0nQ5eghRNUuREyShM
CtplFo8M/x4a7PI+VZm41X5cVkWNfVPIPcbXvgmZajZkXCznolwV0SwQqtEC4Diewr3mtLTWcsMO
uFdxXknxCNnPe6vNYY/++fP1pG0me+ohw6GfpaMwvXTHwF54NxFGDXP3A0VUIN/GIKlqz3VtdSMz
Oh9QNSwS0ASSpGsw4osKumb57phYQTLpwyvo3rPHRdfuXZ1/VdhlPp4+5WNb8nredXX7CCrGI3a8
8ttGbs5ihddyQMdK7hsot//xk98RWH5QuROp01XnzTH9hvUvh8uH3tfaPNmiKCaMU7N5OYjodMnS
vxq2qx9vxLx5W3sVuIy11yYd8NAoJm+ig/YVU/13opitsXNOjyD7flE1Md3ImsRTyy9LsxpcXzLj
0p7ZUWAP1ReDht/Pfr0MHG2Hn/KLoPXFlPoZgDx4emrf+NikLsCXLWWkyQGtTrDA8cIRMWxyNrCA
dymhXjuwJhYdtqtCmDLwG2DhtBI5Boxgr0N7DP0pcRuyXjd2JWMrpMk6j+gFyxZ2xrCmL3oL0vBc
RkEqOj5Knl3+OKZGRr1BvNLwU//CSls4q4L8s3DD+RQxNNNS+bcSft18vaBId6PqSmjn0/9nkAGD
Gx65DNZn4wlRbvYgRbLCdWoU1O0iaW7iyTxgfZ9waaVXYASMlU4uDXmsErAtiGpUbh+5NjG48R+C
7eLKV0Godlq1qX8CX+5FJw2qJ/7hhJWoQUi2XuwAC5hL1T3JiEt+HO6nkpfEesnt+7o01RQP9yoZ
YFD5l++loZBkp88ouUXZ65ASKp13X9aFIzfFEi8JM63MucGwAUlQ11RGV4b8e7VJZ2jOfSO539v6
GEY05gJlPGptAbBmbNtZql1rvckpwF+VwOJUDubfW5E19cS8plzd5J6JuOlGXf9bFPnd0szhb2H5
QCGJQQeA0KhIO8L/H7c7fofCPS+bq9qQ/3gmSgp0Dg4WQWay8Zl7KAjSL6ZHynNnShGQ76stIIzN
rvKc/LiOoasAqjP3cZQuB9ixOCp2erEm9FU8i0wKkrJv1o7Mbi+2fY9GONmfni6xHpGHvBsTDKEr
2GjZwkPkEwz15aojmX9aGrLUalvlP0N7xOZkBtKcCeefg1DcMR4DOgtqhAU78E06MrYIgT6OJWrD
ghuMl9cE29evZP6/LVa9j3GFOu8iG4H9piFSdy3BvXNoQES5B+AGIB+PYaO4ZdfU64aVM6Cy+7Q5
pZXL5uSO0g3L6tIFBlTCevWrRngv5GtvUk9W3IwUWpftrIMg3wZMuU5GhrxvORh+jgQFXCXLoGbX
66u6qOXTm29Cu7Nn/zf8HGTkg864OkOYFg8OcuegyoeDeHD3xRyIN09UhUxCWGr38RBFt4ilaxUy
k3x6xkrCAx5RUiLW7Il6lAvsqeJnOskwRrFdHLhkbKLRdKjlmxTRSRD1ey1CMmAtqqIHCuLEOQo2
v7tvNBHdDHmVQlJs6FyLgYGyNOUq+nxM3mjIvKww9TXf+7rJTyQB1tq6LNDE52WZezC8OIJOJgyh
kM1JwhJPbNAE+msXPZeQCkOROy2zrUdrbu0IBIaWTg3SQDf5wkN+OMEaS3xWNatRs/5RsvM/HK/7
RZ1xZtAtj9RX8aVhKpFwMAoNG9BJG3WY5+UCW7mBAa6Iinz5RZu4bdx/LbcpPKjimNWY4IBeO3CL
YA0ld8P6YfrxTtG412KKOlhY5qnxLyDZnBtZyyTBlWy3TCTvZPzc8WTTD2n/CSPz2Pj0Ds0S0FYs
zQLC/u0Xi20NapD/W+612IQt07+QAcA+ZfEIKatlpge6JzuzJV4f1SG9zXdoLfemE5IhTAzaGwGu
nYmq/1bStqXklUMGa+7c2tGRjyxPdn/FBq7xQSzjKbBtr3IDZQfMeVc7JPzDMLClT380HImCnRVs
aUPnddbD0dPqvVw7T61W8WY7F1uaRYEN1Cf1FRP62+pw1xd5CuR3/MRCU1Q1AzMKtjDDpAPMJ1B8
0J6OXBMC6Wm7Wp/Gk9J6rwVQ/JsQRZTpfdQPC3+RimPQ4cRmws9uHT8BZ8CJriRigoSrQyKoM43F
/Tbq/B/5BJpncoV1P/jYd/FcvpvmHOmpSlIniAwmymJwSvJsYz+KwbYv7yHpdZa83QZ+E1cbn14y
F2S7hmZwIbJFeJxmTy5CD6cwzxRSZxSxklOP1VQ2jVSfTiKlxkDCzoB6LX0iT0zqfOkOXdjIcE7w
qFdm3RMvhcuaQvI6C3BxDg3dumluWZWKAkninWLFDCol9xLuRSic5IH7jLZ45Or90PHth3ycAhEC
fcPicH9yz8rbCu9kGQXguSWbAHNHML9J3b/x1bUio9/RH62xdD0z91A0ZmDVdAN6lKw+b92FvFna
rFk6LbwjKF0Udg5iey9F0KadwDBu4VjuL5qeBKLublwn8GKEMNtiP0WZOVWwFZbsuynpzAGkE9Ad
cN5ZeMQVvTUSrCoHw75c+eWZBXTp7xS7yTGA9B+tD8o2srHQez/+e+S8ZtEMHdskudsxEgCHe+Of
o4Rmsm2Pp2qm5wgf5QUA2DqzL+IdnI/YUk3pR32grqq0UIBrKfRvBIb3KuDMoeVZGdU+jV6cN3hc
36UVQaDP3q3ZmwD/Dj9HzYx6HFG9Wqx1QdSLoLxT5zVhNY8z+39Njr0iqur3cn29Tzsu1EqO0dq0
GUFArwAKOsO9Svq9HkmvlbF3Cz4+Ui3QAogF0ZZKlh3yRzsPkj1ezES4zo2Vu1QUgTzOkg9UeGmr
A+s1R+UpfYx1nB86F8C4JLVZtxEuQvOoq3VrN+zVXHrfVxK44dpeHlJtsxA9vnelfUQ1ZaLKG+qH
ahVwSy/iZZg4SqDcF3oULTM3VCSzwDe5mvFSHEJIMn28rQX47rbXT7ir7u7lGJegrD8W4c1PCXj7
/rJkhuyW7mWb2TSLe3o+/zUBpM/m7lGAbUeZ+DYKvjCnEb75/LoPGoTsTJYN19LEX4DayvNTz9m5
sZ5sWVTnQ3XZ8quaO7u0jdn/561DZy3mdgPedSm8/VOig5tl5s2KKlH9JvIi0ulQdZeCnxODAQCT
TUvCooSN5z6+1gyOzzTAJAuCUloZ10I1Gqw9drXfBBUn1c8RqgOeOCC5Tj53ZruAR9YCXmXuIhEY
lx6LHrRHDl4PJmRw1PtqemcQu8h0mWu6p+KZq2EfVn2FM6CKijEnTf9f4LmTcpPbb+s+Ph9klfkP
gg1BGYOT2QX6xGcAFMS32bxTlaF96YHn6bOEWOuvRRKc2MMyc4dcc5uQkU36rm2Yla1xm+xZk4gu
y6SraMEwROxp6ni0/w8MIkPyFiTAMFiloiTayljlBeQpZg/t/eZCrIz//DIdtaIz/5zShIWUjoeY
Ry5YUgkM8d6ipSRZKINZrLyNmYnZS26SNpiKvlVcSp/2E6gPlNIooJ0gsGl1cnnDnIWqFrJza2wp
seV9aaIBjRJ/G4jAh7Zijh4NK1EcWOqmY9YGBV2fES4IDGAo5MSqwEHJaHU0L1r9GqKxTqe/wYlc
oWIcSQEzImyiYs4MPrYzRe9+xkq8pvHLT+fznOvJ78g49vxZqz9wmouxvDZ4/12GgqL0O1PrH+Gq
fCzg8Ee9PIplo6VHPZ6LX5YFGpEdnMPzMB5HHqVwpY5OmIJZjtrF5unHoQ+vBVAtZ+aI0bWIz6B+
Cu/hRPnGByrGVLgeaaYgdfpLrc1cD6g0wbTmVSqyMqJsHCpXCcK39gjcKYXC50UxdlecK1cXMcI2
vwHrrmOxh707jmXUvYwHn8hC0YihvOw3qr1SyJxxSCGd6bStmCUdYKzE6ie4WD8Q95vwxO2SNrg+
0htfNWLGTuDkaCTdCz1BAaCLBZOh0NLyfJN+XSLQg/CVDXprjkbh15/6UXSb9mjz17nd+LRTbYBa
TIQlUM+YWmR0tq6L791eSNdaDuzeY+WEgnQTZCQfeT56fSCYpChqfCxPxjJl3YJ5dSeOM4l3wtTd
2eeinqPU3LUdvntSZ1DOI0hVBCJtyrbRgCwRLOPgvdbzLfSv66j/Ha+tZnPyRJRsFSrN+HNwIf5I
SGnVZrrZ3EAerECsG6TLXm9TLqf0iklFKCjeBpXffGbJceBNWWocsL2JDmJZNmlKZUUkSxd8wfy+
gYpSysqmjjaDl23SzNPVELOk7chXPRQa5eSE+b9jko9I1Hv0UovwEUGopLrVjzphlfmJjv+BBXCm
vjHhgFOCAykuXjLfCqRb4g89jey1FLa+umw308/2O1Unr63K+FK4FivJz3a+B9uvmfTYhIa9rqY7
NVnfmqdYMhz4edlwOiH60LxSHJu8wPo4a5YgAgmLXLrEQoDu1AjpOmim6BGlMt6bZkQ7/yYVPAuc
Cq97+k+qmbIYnmXl5AHFo49cqtyk3BVza7gUeL76hacwLQofQNnTOPnEvra/UN6lh9IlVFC7VJdN
b6X8gjBXnzwixaI/F4rCvvUW4/yIKCnwlGnEgMUVMcAj9Ya2LX1JhW5cRrPMdiTGWYzTj+ZkUn+2
OaWhEGYvil3s9Cw2jI3dQSHR2rLnf19wS/Ee6q+LyZbbsRs829BZeVcsW92AFBFy1Ln/zkbp6RD3
tNOncyRjB5gmfLHf+MeWWu7rGzqTRN7EFAYg3vE25PRUkn1LBrAFG0Ujquzt8dP25j4LmjvysOXJ
FhkyhlvfPA/8aMYYy12ELJ8Yy3tJsDK08hr61qCrSw9zAfV+cwODhQSGifISl8q3SMdVbd+O7L9+
jgRVYXzOaMQQFG7FNbH9JUt0a3rhvGRfdWULhl6wt40DDqgnlyYfei8EiemQzFwXNSF+B21tc6uw
8CVfmvvUTmpDh+BJpu/t8EzyhUHZkOxQ5VoMI9rMBsPJhIHIh/fn6PdF6z/OgWfS8tsLpCk9hgvM
ir56SUN+sOUsQC7jYkFgSQMvWJMZFrd2+LphDTD76QWEOewz4uGQxxrFWJkU457a9TP232blUXRk
kSYAas/Tk0VRbEgWI/HPWgFOVvph4NGIqGgej/s6c6c9BfG/9sdzj1FYXPshHexvpPoPsCyQsJEP
Jaky3pQgEB9jckkdkzTYBp93xmPNXJBMMHfIFR5qyOX53pAIbt9I5Hzw0KyoKzcFHfDu0GVCwfCQ
I7GqePd/dE6+9/s7ism8KxaOtEzVTranxRyd/zdnVlCy9To4dIL9HEzQnm1UDhpezA+pG+0gS3dO
aHpMqGimHu+VeTx4hPGeC7Vo20XamPswGSGRkzAHWnjphDo4aeSJbx4ZQ1/5cefRAGo4eK+AbFQ3
4VKMu1HwdAXH/LfwXYtx4vkxHqwwCKRCuf/2iXm0BxngM5b58ZYdOi67/b7q9ke8pfFs2ejF1BIu
lX3LbW87eNVshmPjmvd/5He/XX5i/MbijUL8Jw7TIOQsHXq4GptFxUH7SAqyJ2/LiveCxcf6X1AZ
ZGPP4J9UFg9+s8XRI5FZQchrofam0W6NUZ7DYArmjh8gAGW51qXk93oq7vlkd+YV6PHrUQCbKXcO
MISI16O8ohTAbqfaPrvsb3HOLyo0PsBGolB+LnU1HqBKn1JrM/oEmni0F+346lEeUuhryZIzrBP/
GLT0Wl+RAhMUnOlsfyt6qRSLXyR1oLv1zUcWlR8I2lafjzYQ9G7Me8aQ1vu/xE/3W/2sl7aRE75q
ZNmU0Pun+fanra9f9q2mL2KW0+LrGceD7WmrjDU9b5xub3AYXX+H1gW21so7OBIoS9k+8qI5+Xig
aphujfBpFDlJVR2RwjO3S+YlHSllFvh6tK/UmGkG2zJYhPMXF5nrfubIXRd4ZBvY+2edo6nJV6Rf
ksDIkHsfCF1D5a/dvB130/npwKuidb2rtlwlhITV9dEx6eZgG4ls05Cqnb9R4TzEPySs1LZs6Ir+
i1viljAG3bIsP00Ipc3BBUhL3K6ZbqpqbLzRqkbrpwWIxHGCfWgthj031aIeeQn9gT7SmOtEEoVa
kg5euAwwoMb0RRpQV//9be+AgxgHi6rLKUtQfU5GNHnbCKCXswOHaDqR2Rxuh94noSw6aj79cB+K
OEceQCXPTrdjPG5Ue6/0CtrV3sNXPMPcEqXTyTxuYvjEMw0LKRnNQI8bK6wxyyiBrlUdQzHt61l+
sPuXIQMdhaRYylMfEA4WXOuoiSLrMsSHhBxaPdRuX2AbRtayxrXE8xNqDM3a/qa+aehCoiTpnRLJ
rycorOx12vMreMLrGn6cXmSnHcjQVejeN1LzP89e6hixf6qn5XJmFP9TqVwr/FzA+0OcYNWhb6WK
Qqqc77QMhsLAkHhGIFwQHdaYr63JI35lkz+9kmSm+BUWq0Mn6raCyYC9Pz+pnC5nUa13TGYVDmzJ
3GVFKcJ3MQoNtU76JZEV0mbyORDedyWER0BAXq/9w3kvQh3MX8Y5lucZKxbuzfFAd0GHVzAvPI9n
JKlj9PN6+lQiysUkmIyh2H55IxnvjpO4A3ixAUvWHKcia5m3xwllCNI6tBa/lHteiEkQha8tgfYl
Lxh0Q5RanQ+92kSYLub3OmVp4bo4jayc2MzjMwsdV/5djpmAoSjW239B++yHz0ePh2VKWwxN9YVz
+myefSJT7HaeV3ieBAdPINWuQgkSGO0LWLMCJphy0ssyrp4uiHQryqUTELo4gRKrE3FLlclxrPXh
HSJ0q0KO0FnsCvDBIvTB+/b/XXuSaTnNM4NCxKwxYryaTcWcyt+P42HdC9acCU5YdPBwVeQmeoNR
66on/ISn5qxUtGS+AjP4LCDWI7VQh0UclYDSmEyyILy7Y/HwNjMRigZT1c4IqCyVzyPv5fkfOW8K
q8hVYsAmYATjjjOxrRTh5EQITIAaz/aecOX12ykZMxKv62mHbtMlfsONsrr4tLHHOhVmLW7APCb1
m9ZIBzX9x54hT3jDnilZoATniMf4PcJcBpUTVyYBxx5+Inx5lnEOXBkb7rbabY3bBoV9LBUW0xos
YPFpVzHWwbB34yLT2eHz23mBj92Yg1f/y/LXQWF2wk5uIs+KrwJRSM/WYvpYnLq2Zu19j6iI6bF4
2TZBQzuqhxMAoG5PB5amTdnaMHAYoA+TUiFXC5Gkzww+WNhIDEaQM/xKqKoJsVjbVfq5BdgztlPG
nDxhCApfSI44cmG0LSgD40hQyGIfQlWYDirwXVFXSeTDDh2KX9tki4KWOsF+aWONG/KCuErYwUtm
nQHNoJo5EABXer8FiUgAmiicww8KBvF0Eb0FE32DEadlleDukWucnaKy0PpVcSHoYWYljZXovypq
mpQOm2AIycsZI7Nrrlk+xbblm5rOGINeDVaI5cA69UvhXhm+LdtrsNdjyhjlYWCyXUmq1u6KFUP1
d8qe0RlwMp05cmBc30hBIyFe39u6aOkFYK5lupMafREBVRE3BNrFHz088N1Al7w/dQDTfMn8uiaF
pqpJEUbGEQ3fU0p2Yp+APuB/dNW0xew13pCGbUAFP6Tu7/jw4lHsMGsFf6tNXXZCX3oBEPHtyPP9
BSr+xKegoCtNHmyBKFW57T0MmDlCyvOBplAdBNjFhW4q1CMPzauOdkZJvcLuAGTNVxb1l7bkYbRd
AWrHlMnYce4H9j62xGXctMOEGZQI+WnjXEOdu19RXdxF3nfujE/KaQ5TpLf46txYdaetMFJ36FyO
KARMe1lgWXXNQDCJ2PvE4UYqIkZP2WKKJy5wUOKjCWVB4TRGoS6dXo19Q7WXcig2tUrQ2CxBqyBi
nK5tkhyHH+r/FYoIsqInFN/mxV8XRqjb4GXsOYhUyhmRjd30U2sJulvXyihQO4TbIpzUcL/1OCmB
XfkKG8a7Mg1og1IsfXs4bMif3ZgsJj1D4Eid7l0HUFJPrQyPbLybr8bs1S3L5LDPVWrtwpTABAH6
DUXTsx+0osqT76TXQSHbgl/eQ1DuUvtWCU294uJikJWvxqJ8F1MBSjXVt3qreWgVHJYaq7rxWLpx
3876/T+G/jUSt7GMoDT6WLTWU35QZnt6NuQgCi6nxpAgIwGwPV3aW7OPVyoy/1kLgA68BQkibKEx
qL7XzP5i5Mkfm9IDI7QOwUq1MsmIXzDNzGsnupTJBwSApKWbdAxt95jsUSwaBe2gZ+5iK14DHbKZ
m2xKkxaBOZRS740EyYEoHICsHTz59YDkV89n7+ygeOO4QASgUCEyzXm8yi+Y38HmcsJDXR9Z6Csc
KJlrxwzt9fVZ/Q+x3WwHM6hKN+JxqgxaPZb6rJKGAV5ESiZqtaTSXlkwrRIuOW7UHGyxvN0rXPCr
o/8B0s1SrQPOlgKse2+D6rRfHv2zqMY3E7+DMS5eDCPqnZFiqN7P+gdtC3hz1OYVbJqyTDBNn2KF
2YLesaRmjwYWG3K3kaJbox9ITkzB1qNNvSXQLVmi967SPRHnTKxDwGvFynz9M3LQjT6TAaSs+7+V
z3v2RtxpdPQ7JFpfvadTmPVw+3x+CDd3OnrJhpO+4fSlYEW9P4oL+3EgNoTMHWKox2gY2x5rTDro
kwwnk9CEcRAgSJYvcjoNfKmcmp10PooOOR4FZGIqOtBleXcBo9s4kM5w7c2lU65HnCvtwPhQoIwe
Suk89WiZlpzjhsb0KxBa91tYMxxlI8T5pZ7zB8l83hfB9hfs3sEkWyAm6aW/Ln6rhavyi6c4mdjp
/2T7vTTr5REAKLpmZF/uWu/f5bT2GXVk4gma9YrxGL39ypvRsAYyBxVHS5dnrDlV8MktCsttD4ZF
St3mRt9ttMnPR3oVEVo9CsHpgHqD1yB+QUpSBCENDs//qphPXVDjzWgAc5Q6R8Ij+JwF9x+rdFrj
6bqmCT77HrEL83pmc2Gx9fzPh6SG2rJh7fSjC0owtH/PJRwjgv7A7ZOFIr9TOEhoCtEsTF/JaSmF
mPmdEUkRvYMOKFtxFHKIjIPZYMDgIC9eaRrW1AA9QG1O+nCtpvsrTpktxIuvwRrQ9WwgPL4icAwn
rjKTxLtNDJObekrlwMjvXppUlPxphsb3WY2YEJVTNep6x7n6nV9oElHHOapwtKNN3LZcjLCG/TZy
06y17TdZJtJOAexWaQjtEu37usmuL74FSlfqH75RIteWPwmEw7ae/XqXK9Jypso8LKbhd44di5+w
L+6dzfyuv0ZJ38J2ggK9KDQMJVuFlsVUgcmNOJX0kMZbfC2Bs/y+t7dVLZ6yYN9HCXqrpwes5xRM
erEucW62VXp0+RwcjI0cQW6imdloLKwTluVeArK1VFDmvV6NUvWmFf8bHvQLTC/UmygdXhIa/IPv
TiPyFr26RxRgShEeYLnYsscGdSztFhfVxJCb/i1adYls+cN9vFPHgJem3EvS3hdJ/hmbBBqozpR8
55qfvt4gfJJeAnN/xDM4aDQ+nr6RCwHGBTukNN3a3sNKNtsZO83uBk/lwolRhNIpfgcrPJSmsQvr
THu12EibDWFp76AzPkIvz+rmBA1ejPEH0kA+jU8FMmHXaBBr9tgSFX/bC2lAX3kkDFdwhJEcfOFE
D9m+f6h6GuxzOO5v54G1Kscb63sdlpM0sGkWycsO1WbYupbmYd8gW46d9/nc2tptmN7AYrBT6M2X
kSSLHKdX2FeLNKSSBPvPS2KbYsnCjbYy2lB9mWPCiCSMcRbfwZmF7/2wbVZecFKaVnJ1hubHCZKK
/gTFqIJbqrHJftbglGj60ngrxhctgbwMxMpTaFsZfnXQ5YtlJremQeaQZqDsjEvFva08GQemlL/1
QKoGewqNWM7wliCS8h2tJZzrC3Djt1fkkM4Da+7FSKFbVkqjfBLL2mQiqBHSrKPAZjE9hM/jsicU
8z3UZb+onIRhBzWeH4b5C9ql4urmkk2axxxCRwlPTlRVqcFITtfHhd4GS+SXm6Uc3XaIoVdi7P7X
JeJCQTI1+vXdIGGrD2FP090ImkM9Ps1HzhdmRib5SHKtZWyuJMi1aUgSymt3NQ9PCdXl4WM+dTar
MN0bg7hF0HEuxoPHTNEoHCcIshL62ZpxTPt3A1IoO9iuohtJbHfIb9Jxjw73Ub1bu7SQPxuPz1x9
CIm3v0HbSsHyF9oEuY+v0wB5kF+HYxWRwkYyes/hJjXqZHXG25s94IUsMZq8+7iGff3Y77LQEjbW
P4lqIcKOLLPKSU0UIxOarwGm8BX+VfWjjp4HCfY/oU6bJq14uYJRNNBms8+w+SIV1wj9d73HnJSd
WT/9hEvmVv+RQRvfotjNqOu8noyuVW7hs5OSIimf3QcUyvalKaqLQOjwTUhRtJOJygmH5vTNY0aB
yJUwNawWU3I39m3MC/Y4MZ+lV7WN4mz0S+cWYGBOPTDunYRK0TNQrXF+XL+qwoLZ1m6Mi8Svnuvj
3hwxxCkVp35yrlZNgJzlcH1L55pSN9uNb6S0n46UETHqxcTghzEhpDogu35bPBVlsZCkTUNH5m9K
W/Fn23UD0cXeQWsDi5robpNFJR+0GZx6PnYIeN1O508R9MDWQLPthPV4+q9P4pogN62d5Crb1fZh
kXo00KKiUYPHUNmbUkQztrmwcaveNSceB/eN/n3UA5wCdImT2GnKVFtfxxDFrwfhJw7Nwvt71BT9
9J7WNSxL/pEUxTG5WJnlzxen/kVwedBmR/PmKqDcFFxfA5Xr6Yxp53g1gqqObdB7DrVkrDVY+EDl
ZWKmYfQ9pgVr8qwGAVw6KLK8wecZc47bF1j/dVmQKbNVeFh2ZUe9oAcE9lmafHayZhnmqHX+jQom
GAG81kTUHG5ZnRkWc2UaigYUxaAWKTivs3FnhbJsorIUwXpLCbUdHptg1Tq4qShBwRO59eeDk9dp
BWrRebYJ5eVBu9veRQDlqSit8/eS4cgq+uaCunkap/nJ+wTPtX7RKO0htjVdYRp2kEV36BYFxMsE
xwXER6/tbmslexPgqbBlfcpZgNdSFJpoyDACquWDSdOWScuiyB/0zzZbabqeRObZqv6OWZ8dE7yP
KOVlvzTGYn2xzY3pH/Wq/AvCS+/gt8iFFSHdY8tXLFYfXv9U0QIyLS6zA3yWCJIQ1KUVJP1YBCN7
olONR6LWXb8elIoGLEix+GcbfL6TowjBxJE/x3Gm15b1dYaEDrg3O4wOpeDK004NeHV1nOv5kxiu
L6/xtqxND9PUE92ewmSVWK3quC9YAP7yrTbZYRXBW0MXF5P8Fck7CTuSXJkhRaY1trjALf2vUpgC
4lsMXU2usGJeQ2xC5x5fU5/zbrgR7/1tLlS593Ixpr1khgRJEb1jhwI0VZ/mYG9a60JubLUE2rMn
SEFyGE6i6XyeZLDatLOQ7Tr3gBKRaszxTa80NDih4VMSUlZ5ENpQWxPAYBMUNVA7fwXPszMGI1S6
exbago/Z/dCs8QhYb38To76ktwlNd5kGa7MhQ2k1TNXAzVde3zhNfRScHKrFbwU9LjAGz0KFqI9V
O1nbpdaIjvMp5s6R7ZlCug8n0xZ+UoTuSUtJAMNwP1mVc9LbJ0ct2b+Oz65TLfJ67dekligedO/h
SdZr4A4++w21Y9T+KyoSHfYEWxUHHqgFCz7iuRJkd046faWZLSfLNyy7NwlBhpWHOQnuHMlQtVLO
283JgWK7C50h5QIHrspY7RVbBbEzql8tYUCpuzkuvOUgOc9X1rYFpYAJJR8OOLFMV3fTRHYIvkGl
6HuD1vixdRoiNZzetHroQsRn53JCcs0QuAC7gmR/c8m/sRa8K3hATx+83Mx7rkB6cRiKSFNfMJCC
YDBMoLZCsWgXS9AtRtxvO7qTmwHmfPNwdoVL0Rrii9x3MQHJ7TDSB7CsgQ7alb1GEm8EA9BDgv6A
johGMTz94ZCXZpH4fKISqKIo/9ELUZbZq8x4PsUOMhevEQOrNeHaPO9Lv3IYEIUyXZihzQ1/T57k
P+rRbO64kanlIsEE9BgisNGcehuB7I3flZ7Z1bmlN62s3h67BsC6mw9h0PdNLKfBAToTt8CFIC9v
bdsOoOG00x44twAwtkkQ4NCSeEn8ygZoLD8xwpk6PkBBXVH9OnG16dD7mULLAIqvxorjFS0SyePS
QCo8jltiBJ+yWzQ/jpWlibSw7Rj+VTcEBgkfJA7CrLkO+4/9HYvsXRVUJ/FebNT07QvIhBoOqTy5
SvjK+ODoSAB51ucd44zpajX6q0HaNxEk5iENzLS/chtUpVCV53rdgDyyX0GdGp2FiEFVmUMY4Zxe
b5oKle1l7wip+i1wzGkJS+cYVs5B9xNTnv+2XyRpMKiS9CS7xQq+33pSVwgaLG88oKBXxH4EYeXw
2flZwBbaZ8lE8l1/9380PIB/vsuFt9HVTSaGqK+LAecLuk+CSgDwKapXbXdYgMxEFZRFPCl6EdvG
iS62r7CPbmL5npQEoEBaEo10wPz4YTyCUDHWSqs1g7Mw3eoy5XYai6UA2BSwtarQ0ffXAVM7yCKg
j/IESydRsAvlKNiT6D/XwAPcLmyZlD6Bq94AOpDXx+G1vJmUU6VRATiEitBQBeyCZdkdfjXnqFwY
AI15B1zegRmvTEcvLpzdHDLyCFzqKLMw8eTk/DAqDzWj9cJOSCl9nCLs34+sHHDJ9JMQBPl9T7Tu
EQI1ZgAsYJlaQGaM37yW3k7APT7+bTpcjohHIaShLxGEEkjDX2m7X8fC6hitGn0O5iAAK39qR+HZ
PWhi3pDWdbGTnp0GUGsFRivaG1IbJ39CbnpDBIcXmkRhfmMWoXaeMgmY/ND6Jo2jRMPVFloe5YkM
xMWTNJy4adQ6qQl0l/vlYoNkXHvkK8R5m0naeQCmwFv6KgqdTDHBK4nqQt3b2OimcZCG4XbRohXd
2JrVmKccWDpZCv9mrJoAeLxjq7wFKXxHdP6D+242j/kEXygg7AVR0at/9rrXifSHnkCElBPbhKQR
YTrjz9sMu3FT6C/CnJXBO5WgSQNeXm/BNTQmYcHJLCKoa9Aohg1U55F/M2RhuXMrCriWsgI5IE6L
xrOBZ1/I1TRNlXQzsciM7rjD0y91DiB+hmsbnaPQZ54hhge1vh3syLdYeUmYKsqgnnn+CrcXc7dy
Q2FOVkCG/xpIp2YWIzBaBhPozXxW2RPQu0hAwoa5jJCAHCPdXfsEMzuol17b8IG3zf4xCjklpDOj
3O6kHrNb/X2S92nay/Rc60fzZAyk4C8IBPyJfzPBXSNq8iGScXfgSB1yCDTPpRDRsKZ7MY0hMTIa
jRCjxGKDDGTS/3cJhj4a3L2m8XA2EeebS1NhEhQzhI/9eotnwxVw/RVARuoxBTb58akVq/uPAF4k
LINOEgHestZ8t3VzLvPbleyEFS0dU8OcW9uQdz9B9Smf4uYKmE7bBvRgMCNeyKOX3X80yi+sqaMb
rDiWCUPCg2djNeFm4J7twlj0wTXcfg8jFX6tUaengArqD6EYJJ8+rFsB8DfNBg5ywkLc4q0WSJPv
alC1XCL/tJAQv/t5TKw5mLa8yS21LdiMfJi8aV0W2j2dP0IGOHuu7FIhjpBc6fzSflqE2XJ609I4
MT2OEeHorGI/VyOdvb3MoTFZqvum/jiMegm4Wsms3I01W2JYi29U3V5Lv4p1XMZfh3EMFQcspArC
Bnyd18TIyNdqESnnvBA7ON3kR++t0wtS/uMuOnv4EgcAyP53sWyDt7pNfrqEd61SskhlIwid9YwH
6Vd9jGW/BPYxL8Za1JVcoELyS3zoTfKRp9i9UkuGnotFjh+O2yKikhBL2hluySF2tdn3wJCAwXmL
uX8+mgVVizzvLXfEGfNj0W4o3AllDEKiW8Ts5eqa4N7alxg/JtDaj3z/94b9eN4L8Zs363Xqh4XE
/jwMP2ZUW1+RvDWWZgKprnSwtAo3kDrPZrIWJqPN1eFhuIColJsnY1RDud5FXelZ7s2B0RZPx79m
0MbQVs/gH7dvKg+y3UxOStA5Re2rSuwCj1UBROFJ4zcDhiCmQUJGf1ppV+OzI/vP5NtdBEMBmbii
OYAO9MjFwSf0ShBVi+d5lydjkLf433+fMFJyD7yxmX0NPYW6iwhgDzVm07Bvn9FdzstZShHgjgbt
vx42m/pLrBBKAcKqhaYNTNUjOKVRN1aX20s/iTekqoPH4NrrBJQ1HmQYWB4zi8YXcsGtzt+0U8VE
UVb2DNLSNwIksWv0z3czcYPVl23+mKK5ls4TdVSruNFrbOi1Y2ODtGXNl3INA0b4G/9CIMBnrHsK
Soud4syceoEh7vDTZr4B72qON1+s9U6yM0/YOJiWrAgfjf890Sd+9MPKQ2CIOjG85m40l1ejmlKk
NprjubMmTXPhVsIFSkCPKrHx1LpU2pn9+6bBvyHieBRilJrbdgCl5WwMOLhSm5KrhaxLvhL/3qIs
NZUNJK4tnlfSbqHMCKUB/VsD0eHoNp95Viv8/DFfrXTqJOXJ1Z+eLqWsKW49llcX1QgMuidLPU5d
EkOQjVD2/eLf7e6UJKEE1yJ0UaqV2KxIhFEipBsL+m5QDzjDX7O4DKcLkml2T1JFFwfhLuxByi4g
flDN34Ol95IdCE/oI76uWqfW5fqZVQpLMOFWf/TiFaN+cTARHetbgSP4NOV6WxOzBs+Eh5stDZUP
u435armaRRFSnWgVs5CBhZqb4Od3CFWdAd77DUuzSl2D/iri0Gr0Rv0eUEdK5SDyasIqwBc6eMBR
WqA33sqh6DoG20a0uAa0Xjo0mAfc1M18OBvggqn+JqbK1wb7L4MrCLQV/9Uro94BT3Vy8zzcOmQg
1+ENt7vA6Ksa9WAy1MwdDs1L8eX8ABZx/r6Nz7wrVQfzHPB3cmPnpJse8j6O+2vTjNb5VxNee6eS
WoaeHPffJUeD/ao62UVqBKYtF58xy8iWjieySS2usOpTjGMRS+HxdUfib1NxfRBKGuR0CFPzfahs
0HUBFu8axQNpyHQ8f4YUE4CxdBY9Oc/I1HZXwCkLIOEDVytrc2FsmUn2scoWvFdCs6/Y6Qbnr/fT
t2LHgs+N1F8vW4VVY2vjO+pyLT/1EvgEFr8eEDnkHn3oLoyfimwhwFSwXHfsIQ4FrBvJR6CCgh+n
WSERqHNLmm10/4CaJZKHZuZrrZG2keXbbHUs1/Ocbm67dQsAkhV03M1bxKYx5xnxX/HDg8FWN/hn
RkA3eGl11LuJHKyZUPZlOMr+G/HlSwFpvxapdqBrWN5OlEiuRo2r5g3PiYKX4B3l4fhNBvxDom1b
R6aXYSIQXyiHl3Ra307n9ICALpoo4oMwD/gl3ycD4Ntaygi6kFHOKvYfYoTShPDFjMgEk/22/Jnp
XVMtVnMfcbt6MNnu5yiYzjmT7cifrUVvnBQZIzHZNs9CrPzblj9m2458AycEBpTlbTnR0fG1flK5
MikwB8yGPXEqKmjpxDN6JPXkryT1ar605QvhRAE6VYK+CvsjoE9ddnCERPlC+3JgRpOP3L9LbrEM
s+839fQK1E+eRnMJuyGkYHCJMfcpJUDMfMmty3nNIIr+wS6n0Ko67ogOO9XqCiqinLPlPoR4u3NS
iCK+koOU7m5YD87pRXxSD+nidIlMpuMNuHDF8ABvcMQQ4DpqbtGNy9Qn3g/uNQ97gKRv+0v1JHD0
GCktazRe/q+ICjVMh1YZ9a+JJVpYkwY/skILQl0eSfxaaeqpB5Hg9epUDtp4VjhVQMF8J9LULgcz
aR2s5vQcYqD5g9YsDrEATbVUenGn2xy9JOxZXAwgrDSNgQhyymr1/NfYt/VqQn5FODg4zfm3bQ1z
C5iMx4ZAz/E3QctPKmj3PZoubqxhziyda4BTdCzNzZGWlFyPvopwbIbMdNl0jN8sS5pI6PB2JSNY
65EO0pSMO6lQFXFC2sHZD+NT36z7bNfHKbOqQ0rY+7YvG1d+8LWeT9YPjnzExrzEa0JPWcoJTC+v
PNwoO1iP0T4lKDstOlVVIowYPO+l8fiodW2+ZHqI5z6dYEGKfvP1qhssLbkQEDW5/4GbaPNkMmn0
PU1K7rE+ub2HDWq2RJr70WCKmrQl7gY3FtqrS1K+psOVqCnnpZbcRSLDHoco7Sxa5XRaZI1hMR7M
/bfonPdGItCf7xyf1WKFZgVarzr9urQUZbxb5GW8zYlxneKPTQApQg4NiOYBrEjnDupKXS+F6ryg
KNqpWiB0ORPTtUdB+GJrraru23TgF+zImrSoGMFjkrU7jqUkR2FwJB8rWj8MVbiGoqhj/IsWvdgP
Elp7n6LIfohBfdt7F6l+6uGvfvoi0WKQXbMMqfTWloWeIhJE/zPFBXm3DB6rC/mJVo1LpfM0arpW
MRz/+X2TZB8ToXXGI78IJHtEIJWTEKBt7pkgHzo4XO/zlU9qOpLs1Yw9wWLXjDoSbAPdbV6kdb6v
39tjiom+qhBB39rU+YLBMdSV598067NeTq62aLBezCCWgVOJC52HgFe8J5bPT5R0x7EZQxgfUWVz
Kt32nrnp1+dL2zCP6m4Gf5RZMZ1yTu/G8r3FeENNs3n1ZXKjGQ4Ja26LvDz4ct1v2Tg0pstebVdq
LcS5mNQNstXTFdwSiFY8cMF1EWwoNH0FZUTrLUmPykcY8ykkgXhNgJbV9ZX33sL+NaWMqBzWX1DP
5c6aJf9OtRpKSsPDfMjV6HPiVjY4M58DXvFjjGA9EfmBkoLCm+2K5XDoVIo1q9GInJIkV8V6wAwr
21RT0HSu2IuP3xpETEhszUsXsIRL409a8uEsvujoO30mkx9xpohogIr87UfQRtvgZOdq6rjK5R99
vEU6jvhE08hhIoOJRI6BXZlhB1QRo70dV5mI5vX3N4vWqRi46MprIzkCXNPklzdqlTHRYDqClkf1
kFkEMLKVoPCtusFW4RWXDjU/cYTq+714eEhtbSjguqVVxyOnVoep7DwBr3VtECSTBeThM1/awkT1
eyDdXvU8aE4fhBBs/tLsgRO7Epgvh+w+v5VfF3STjEQwwNl8TjJDCulXM+P7SYDBGVOVIwPXg6VG
PXiBRCQfEWUE57FlJ4Xzhr6jpQ0as172zzCsZG3W0ZiyugCpusZ2bQpzbKJFftDrDKmzW1WucFjW
9G4I4esnKwkQJNz4Ftv+fyGgbXb9EglXP2IsYC7DVsZo47Fn/BPxhxrL5uXaCN73+kSb1vKUmMgz
QeW8OEaeUgYon8SooJGfCjjmx6whfMIgkL4/N4N+4cgx43C0WrHcSIKvgNWpdDj7A2D9R118KS6Y
kkjPeuph0dqanLM6JEGR84N9xNTufoE1FCZDdAphUA6z2SvUfYUNLiVUfaPm7ygvSxkQyRd/kO0W
JRi35LCwncqPyOxlCWP1oM47xpPY8/Wem9vEvPc02JjWKQs7eRuRUlq4Wp18rViNtsGew63EYnYr
0nGONnkPMLor17nTrKe1QNVxcsYdY/LDsAghvPvdiYrqGWeQ6K/wNBgw7qczD8Z861OYDR1E2mVY
qtbo+VYr/YZZxSJzDmp6cw0Es2xrmrEYdg3Oj9rnEm2EhgmnBDXAUnVpJCKrE4arGY02lW7D5gW9
sPr8Ou/nkaSe4bzRw4P16eZDlilpKXEDsesfkcZ12pQ0+DWYnBEKggg2MEijzJ6Igvk8TI0dmpTZ
habfZRfuie9hdDOLc6YShciuMViWddAbrKVBc6XCU0PqWxfYs7sGjg4ogjNbHIwahh2SDngqR52K
p0AOEUc+RgAnPH5YN8iQL6q0efq2q1R3jfZnzGFczruvEN6hj09MvS0u3gnMg9yOlJtbpvjmL920
l+RAzMFDCo550ccaejKf+rvM7vk/BFjHcK9dd9/0x1ltOEh6oSp+RZb1o5UX2TiW9hhYfEob4AFv
GOXTO+jltL/diWNzd78zudU4pzLIjZGT7WNnY3djdun2uXrYRsZhUp4n0WieRZ0otK2iW6XmALoO
VaMMHf4Lr/J14JmzHa5FFqemtvNN8IsihDr4cnVc3/Pdux6hZjeoBARTlg3d3jQMqkZchJGbFUpO
rDVZ8BWEKS0Geh8GZtU+Ro4mQPDdPHT5AsUcKzpV0kSXo6F4oCC955GofVJwHe3SgxaB2fVCKnON
FlLKS2EC/5+FdOEWZdXmXjh0RUjLKMzjb/vKMnjCFjIG2ccdoMuameqMO4u4J7JHcaKjxZC4/WyI
ht6D08prXZbjX6q4ELXHLMhcB/ZrH+aIR5mH96yMWxV2nK/7MfHMOiH4gk3fxliygVwmqrAeJaS3
LtB5CLhtvpmzaThfaj3o4Jz5JSm78pI31u/ZHZ7ndCXAPDSiYiR69X+UdokKcam9H1ItlPZXi8SS
U9Gwk/4AErnE8AevRH3Pg+pLaJ3QRHckjQUka/2lSEDhMj4+RTS0KX31GRtyQtHP3GbVGwRit6F5
X7nLj7B0fgTohMqtAw5LSqijtW51sk9LvZEzmxS4RgZWQoOxQzfD4QEX8AfKfNP0pTayydWbKWLR
lnt+VJu4dJPX6qk3ZNlrrNLFwrrspSL8+mTe29dWpjDRVh9iYX8NsV028i+LQGy88Q9bpxmQHDv2
0y+LsFucXM7r3GPTWksyk4NpjdJ+HGGaQOYcq3yQlTa5fOv+76wFt0kH5IFryNdT31zu+PGNoTe7
9Ghds02BPiQlk3L6Mcc9duKMrYWF5jP8+kLJWb5zTZgn4Nl8j1ZFDcc8OqYh6gjXM286DpWqNj+3
aLf8GwuqL9EhNiL+kDEE0qq2N+7eZyLGSklDy+fcL+Z65oKVYh02Mw6cHK2tXawgDfvA1lwJr7l9
lWFfrVO5t+Y8OnHGuMV+LF68DMjptE9A+Ah9G+Shyxk8jmSDV3x6zyOJ97u0moKiJhKvauwAdlE/
+GR7vFJDzAL/V9b0OnqwD4cHExW04zKSPIQt9C2jTTWr+ZYkxk4ycNOANhUtgNcsoWB5edAao26w
BPc4JsQ3obO0aHW7d5TcfnRY+uc4y65XE67Qh7yObGmfwLGXtHaPBEyoWVNf19O2w8cpHdcdaqDp
LV2QM37PdhNMKMFwQS/k2+Rrd5SO99YVxCTwX/Lw2KIX073azYq9Lces+FwcsWjXujhS5Ah96csl
wwNENIjKJ+IFTLl8BnPNHqc/3dQ6qvK2B3Ej0goq2+4sqjrWuelGm9bGvqiPSLRXYawhvOi3/VYy
m1S8KjWp34SbLtFQ+ArO4JWNwwkV2teOOWADzXNPLVdjaVzrbjJwluhY+/JE9WefaqXpHfZSRSsS
4G/qjxKXaJcSBNewUWjroW4kQfaC3n0RDstrl77AAH8a9S/cy3SvqIo7kdvU8csgQ63r68nJu99q
tA6KoJ91hUCLWs5RqQafigUI7c49nebeX9IYzmE9MXf9Q9H5wELQRcXNseTclT75mi1A95SKpygi
wnOc2Y/NpDHl/cJ4VShpYO3VjFQoEsX5MI50H9RkE6mSIPbJKXyHdL6iB4+e/h0yHwdLudD2/vhj
FlZOusDh/TlsgPalZ+w00g2UHASZs5fSTa1Q60+viAi/sJeTtvBpS4/lxnJxuTQw3HAtIOf0tq3V
FgB9X6RODV9oOnh3RAYSlf3FQ2xMqrrrrjFt69Zr1XCD2V3lGLQKk9vWRqGsKfiDy6s7YgreK20U
pNnDYwqVaV6PkSG20OYIojV4d2RkCbfcPk+z4JUn5VWPjQuW284tR/OnjGmKpxWiDL0ZUt+0Fnfe
PULVYD0rNPR/dAt1zEhpKG+Sm6tfwcpqyoF1l8jGUsxkJLxVo3wGHTS/dZpvJuGbJvB7VzsJvQPR
2d6r9BQfTkxHUVIodR19Ra3b6wtxQXPVXWHVXHOJXRHBEvi+ncBwoIlGDJUJFyuHJcWGtxtbLmql
/UwmVABqmz+wAJAXmxPEPtmyo4pqbkjKeSehl3SKcwqoCrqoIu+p8DxpJ9aSAScPfdX56KoWxUEn
a+SzoGxLrGYDtHWVKfnRDbPolWu9EhEnypNqHV9R9ovlQ33Z6juYAeDpmSH+Mk1RhOVvGetrjEeh
KWkI3A24YhGvrvUyebzza7nws+Qi0CDRPdaC3tKoNCaTkSLy6XE8dPMfFgzpWcSKoFJ5df2D51Wk
AN8lBPB3z2StjZ1q0DaWpYbIvCKs9FA/0hhe9Ht9nzqKyJVmAMhR2C7ESkHIlSBSWNZgzNEa0uY0
LYYWKoLD6WxXUIg8r7GyCAaq06kSTvd3vNFFwYcp11UOs0aq7+gbZhX3h1gMHfzLcqrPjsAviXf1
sRWw4CtlIgxKn4IlnTVjZ9hC+MMfl6aeGMzQMr+jWSy0VuCbIVoaIonSiAWtfm5o1dKnfA97+Vbu
Wy7dF1DOsSo7HDJ6VeFPtQJQmoP+j8YWS/On68kC/gIIq4nwDSJFEY1HQFAdr+xYkP86C4KkGcL/
b/UFCnJbRKgS9OdQFivCdqxzkv+S4n/rF+wuSxC6XrocvICx7XK+y0zIZlpj+nw5sX/xGLBSZx6X
9NjIvcuLtxa1rTPtW6H3K9u7Sheap86OiRNQwgwo3T6u6hSkH2NdIQSg5TTa63z0lTadCt0lveSN
c2fUzquKxazPFkqptAYgyUJqAKEDe0toUlkhlk2HrZoubuUMQxmDSI1jAiLAtiVYN8DqyXwU4H3/
FD4I8w2ItERbK/39AakhH6GZFSa2CHw7CpS0rJxFsg5q9ud/ddc0T1EVH7ojDjSPlwmr1FoPZYMW
qKuhq3L1+hMBmEk6qcr7lBb6mpZKbWWI77FERi4ER2ODmgKSLKr4mdCNHpi5/w7uShflkb900yhV
XakVjsBsJqFJvY6PKs0W2AWFgDk3hzW1syv5ZxUaOGv28T03FTDqA/4IUYtcM8zDVzYymjas9ZTV
BJJgWGgr5RVV5djs2U/rJ7S/GhJF+WzHxG4ePMfy/2idBpGac2s+NApGuKLzsXysW7NRot5hybY6
K+Y5DXDLFBQ7YKGl7SceSUm03UOc0mufUr+cYERxl/C9QBK9uRb+GAUHddcF87IdLCqIpKUVRPTg
S8vVlDmupoDuOqWrO1VDW5IFl+R239AhffmGqCjwyjsiGGtTJ2kBy/9uXxrAJleRfkxQRilr8QrC
1wsbf7IyNomApMrisKxx5fO10s4RSJv+h2R2nT0UIT6Jp3fdF0hNB5RGcupWjchRGwneydAMGlta
BTL+t/4a3PWT/7kUPsBvrDocuTMGgD+HcXIyty/9MUvVBAh4WyzwohFPKL3GaOk4NfA+zXgWf1Pp
Tg6CLyp/GlFJCAjXalEluxDSVCPNz7C5+xgKdmZX42fg4vIjQv/DyHd9leV5ObQkORVgVxbjzpYV
jOMNf+UDi43yOv1MP7F6A254XEuGcNGTQZPY3+3+4kvZV6LJCdGgNw6Ohrtzk4tnoVZhGBd5V9Jp
m2SNXtBdAn6JwOoLepYEOnxKkpPzQ9e011c21T7flqcbNmlBy3hzYy3ubRhVAH7DUVBTa2i5jb4L
EhlbjUK+fPkUXqkmqsThstY4ASfpn2BVaFln43XFT/WwLjwmEtlGOOFg+OYGYD9N5Mq2/vl9l8DU
ced/CX+nx38zXexZygiXG/Tm66DwQ2Ry2kW3S3w4w2mu6fdR8Ofw0LeE6bCka54/7D51LoK1xRtY
C2rA5BmzhKkpK4sGE8xhajgQG6ioZlxjXIfPyxhebl1Eo1OJaa7YfBnpGuEYEeIekyjtVhQoruw/
TV2Ugm5jInHILAEZE/cge6guT9tvJ5cyg/QNRxwI2TqchCu9nE6P3vXRjryNOMycxwgfkSPabqY9
foEN3PymzIMbV1cCbZCA7sUVucbrYgzWfEzE2wNUz2xZ53PU5LJCfCq2XNCPmpGTTF2JcQqwjyBx
ohGVosu7JEYi1AohsY1nAFFamw9TZPWEAncORdM28Ax8iRr8sODFpO2kVbEsPBixElCWxHzT1L1p
vlWqAP/hcGDRARmT7bwIGxcD9Sxp8yTVz568BvuOlrf6xeZKXpmEHa5zY/h8L9P1bECF2vNt/PtH
HY0DYQBY813zl8IZuOzVO47tKiOMb8d5DC8zMaiGUiZp1x3YvWZRBLmGQ4YnY9bf7SmknBZdAwoA
bYI0Hkt3mIt0CFTQgFyXhKpAGtFcYqS62Pxe3xdLOoJuwvwDkraVBqGJ5u2HcRwRY1Ndk0pHZdbc
VYBa2QN9lNpsnsxR7B/upQz+UVCWR/2xDWlaULGcJ3rapgokZf9xusXPR1szHSi3z9mZI7Jolpi2
FZ60rAeLRiNenug0HZJknmNxDdqOq5cB/BZFRd52AXMUA5zJt4eBVGmviVVcWE/SjlOce85v430w
SD7L30BGXsXol4Rh5fM6Ev3MLCl8Rz7kkxUqeRbXJXU3hyayzv5UV5Y04gvPqeYupYVcfLLj4QIg
C3fW6qxnW1RlOdPwUSfFZd8taaqTYpU9sFGCXv/5jkmwdxPADmgyhSqitLG0CmxDTHnNWqOkv2Jy
AoxY0sqPQAdd5orMqlCHb4gEprouTRoqkXg2DKxfvh8mBKmHD6cCxjB4UN5EjTZnDSFNjlJRx8Wn
tq3hyh6vm95N2rEAo+5zE56MoRej+0PRfi6hu8N2ZpmXUNGChwMeTtDoaDI/maon9a2zNBclYERZ
RfdiF10vy17pWPZEO5jhSG7eljktIAurzI9SuLDNx6pOA/sCAH2pKYwu8GX8CSo8K/8eJlalG/VU
aO+KQqicPPij5dHrOU+8/57Bym2qj1uLbCWGmDJr9pt9ndkA3E5wRFGcfU8ELOYtgfEIdd3FK99C
qXUrCmhOtj47cOcMktYWE5z1KIpsVAMT1RqHZ8JK2xIxwbqLc5HaXh8RBEB5pevqHWOoJTydyTc8
+wmNkIY4k+yPd0vMH/pQ1+xxs8A7/pFzFrI1w3Cn4LDUZrh7fn/Dl2TnPFASOhcHvxN6lD2C+vPz
SHAGCEwArwkdDpY7DoH1IBHcODQdewXZaUnga7blSJGOhZXJ32Q/nMCCTk2DiSe1nW0uFfL6DTMP
WqQz5JQpocMB7FrCTiIj5Qn1mttAD2w6/fA4A++dPTpnseX75eTdpgs/cR/SWZhNFDwzAmAEpaTy
/GD+H6bQunR07f4qqKBbtgj87fNNVJDGFmNra6pnQk1M3dozExxaM4z1dKXyj+C/9eb2n11kEQqk
d9axaYVtBKucvZAfqyoNdTAUkCFohH1Uztus7ayqHJvvQNx8OL/vxzyAh4Fi4B312jmJHDaMVTBK
TxRp/VkEu3K5sn5amtHeL2U5gDPxICjDC09ZH0ANsgbXUWC/hfwq5j509sW4ZQlt6YBgN88/CJao
tXb96KbzRuqMOluDmMUW/1TzE5+ueAEYrHN2NlkyKdOrf3235/ohkrhLzy+KTOKAR08PoE5IlUlZ
0pZXNZ+Ya6ZE+4Y24nSqsDqtNv3+TJRNJCEHDi1QDKiD1nJl193VjLBj46RLmht16MWWIOgw/3tV
yRyGAmRAyA/YrHOImnPXnSYf7BALJ/XyGP/ERBB1ePlslFWbaZFGzdSbzO6rcQ3QZMTbMH3Ty88D
S4WhLQtJ0gG9MhvbqDNzYEcoW8HoLQj/Ptx4qQltkmTCNJMZ8y6S7jGHp1nvuZ93XCgYVRTsQmpB
VfmiJAb2gMpYWASyUxAVnZHCfpHXTEHwQD6E551lwGlfWJ53NYWft1XdmVY/hX0XZ+iQ2jAeGIZO
akFUJA6i9XkBbhSUlsvaFdIJi/2WWUrYl0CXDlS0h1YjYM7jFFY8Yk5e/rUnwETmUtKrM6goM0EI
ttE5BJoXfZ1w/J8yb5IwdaiJg+0HiUTw7765gkn4uKTTiIQEwZHGn16bSF+bFgpk1lc/BZUMiIwZ
khmtQ7q+r3uAbRK3r/qzRYa8NK87ONyRUrjDD/x0IPOqWH9NidaBfynvv5bEW6u37Cce1znpKp4m
0DkeXoZNfmJl6FQ09+9TWdZuVixT3s3lo+XJcZ9HLDe5uwjG984iIPmI4BJn+NjkF8sTFzibU3vb
WARUl58eeXRUMm2dIZ6/o/js0OvcJO964fusJkeRW+HURw8KZnlP0IbvJmpAH06VZ8JbIBDLwa8I
W2cu4pyRE8yPgFP2wxUK6T6O8Ht/wTrkxVffvHD4/BjrJtCMjJgrbMwdlT9oZmM0AqcBuqptYBow
AiN5kkHyXJrI8aXRngtnditdQDBT2OgQfpHrpNEDrFE41utz2wCxV6hoJJCu8J4LZyZhADkYTi7r
Iz3z6W65UL1xO2pZM3JBj2f6y8tsAmwvUAsMznSN5/tNeq7BvNDtNWU+oCfU4NmoPtWXBzm8zh16
MU0oJayyZhFe2oWxsAXQKnqINc6OR5/ZZY+5ORlbMNv/a0nrKoTeXDijglt+us5HcyWSpc/lAmAL
hKqUt1xjDsiYHKZ1fZJf1ecW9VJmjFXea9A56Asbks3av4Xy7E8OMN6+K79jgYzI5pv6Hz0SrQze
idVNRJbtmaWRRA38HwH/2seNMbLp8OFW2qQhcjtyOkbjZVWNAjUghLqBzJdisvUOI+v8+K+1E7hN
/ql7SxVdf2mUQD58HwQA29wNofPoTbH667+8VfUf+bmvTtR3Svg2E0qhNygVbD4IdfjxlLmn4x31
nwuWllj/5R01Im1Xq/Qas4Jh4xDN0Z2aobabX++EfXwqyALeX3tu8ODpbRUxzixmmhl1eTpzFOZQ
2IHpNj6Qw29SWzKwyfZikI4tQELjSjVKh2Bij/T3REcYmIgA+Yhi7hgsPeRzm8l5LPeD5haCeyjt
B0ppZC3Gf1/9R5WmUgaDe7IPRk6/IIxOZ9P+s0kZNEKi6CJRZ/YJJItCCC3Lc0i/YiQM4J9jZstK
1z8Bru72gEQidwb2U/PWP2dGnYc4zMpy6MUvJAR205p5s1iDQVUsJ3tRXYDasXiGW4IE8/CQXwVB
pejDj5uz8VIrvBKIKozikH6iE3QfbpNA+vJlTBRoMjbti12Y2ehoisBFTus3+iVNNvPB2kViTrGS
Vi6T4qvlvaOdRrS4nB92oR+uHyTnWnfOIxWCCDRagWWj+NMMjUisMTrOJLf9SXtU9H4YXSiTpl2H
4YsIssSy/RmyMHFV6EpNyE+vo7uHKUsqH4ZzGd8vyL843+NjSqyuUJrMDjadP9mNeH5M5fux2U/o
5TYDvbvoUOVovCjmH4gzz0Q/EG8OGhEPwVBNIMVceMCaWTvp2DEMo5pv8qivQjHkRF1UvuCBu7jF
+S4JVpQWMaObpiRDJcBQK/oThh3L86LZznP7n9UnKkRG2k7QnCBBVgRcryYy8rLYPafqyXHhkrhT
yqBc/FqIVRo4BWHRWnTH8IqQH5zGYzp//3ngZ/w/9Y033jw5r77Y2SkLgnHUyOliMjgitGJoOcMt
woeDZNFyoAIJGTOPaihL5WQsifIgSC3U/3av8zXSW0tQQwuz2NlzfpIvgT60iNF30ZK36PF1+uMq
yGNlcL3UrQqxTBUsG91WvuDBYRE082aBVznaDqpca0FrjcXYXJ3FFEX0YxckqxVvE0eV8MQQCqTM
Iy+uzEmNd4XHy98ZyPxaNKv8e5q+L6smtAq5o2WDU/rR4kOHJIijfBY1YBRKKWTgWRc2uZBwmzUJ
xHeyavMuoEVrZWOcB39NAIcJr8w9ilVYZ6bNnlWpOgL8uBOZJZmKXcK9pL4vnh/L6Bt1gqe/meUp
ymDAtJbShbhaZ22sV0T14spXV1WjFnYo/eW2MYen9qGJveYb437eu8bD4BoCI4DXQIpSQNZ+2n0D
xOnMFxvU1QLcwgKbtXZ/22pbyWZ6xT4HZlEwWuo/zMJFmP2f6/wpIaBQ4ZRN84JpejweTmDTWxnY
SRuVmAAA9xqBR21a2U3m+xEY1Ei+FQQ8yCRyWe8Y3ru0/mTicFTSUmrVKdZ3GCA8ONCOedmC05CG
LsDv9d9d1MHz+ZEvQHw2mFd7xs96laiVqbbyiqh7s11i+PQzJO6Tke4jxXxtxP9IfPTAr+EcpSQY
jdW98fp93MOscaG3sUswKWXJDuOjECEUkWmUQ+O2h5NBusAFFMlKzJCBcvg2yhx2s9zLURXrByuf
mPedsFHiVuex5aI5wQpi/ul40GrkcUYUj636YwN4W4bEW3vhRH5Im/CnUKEb74YFY4Tde3/+gJ6g
aNO/+sSKbrSDXiDu2a5Oo/ixPpq1vMzioyXsH9PqZmnG5w1Wnh3BedrBAGrnoyDn4o8EvZB9rU5f
dTMxas8uEa3Y1P39hTCZEaStgIZivknHy1+9UIjCQU/H1dJln+WOzZefP4vJLKvsLuEp6LCWfwnB
LZp+b18ol3QGWA+JDRoPwbzeufx2LTOGgazTRd+dWySjmCFlQCVwdFjGeXai2qnDVP2ZWc8fyfY8
2iwOTXkNQ7a4qGAuxeebwcavaen1QwzUQmPOsnIis976zJ4wSUS0d6OXaO9rPgiyoTCRZf4fA2Qx
BX9GNt+UfNUSHNQevrzkLPVEBgiq73XM4qIpr2wz70AW1WtFw51OBDHNjeJOlpu3y/nynYDkUoYl
e2xPT+mpKmlTtFh5Ba6KhPhzr/oSQvTCnfpaMl7iw7Av7UoKLVkRPsxsuWn8zpsleUt2yMMdRugV
snpueAcDHTzweab9r5i28Yy+oUy+e5iLCutJl/U1EWp8og3mI2u4dObhz2yrgJLcCbKXLLKuAG/e
Fmuj1jyL055sr0/cni2L004/BBkRLo61YVPrWlfOnITxj9epX1tTF/7bfEbvssvk1m7VCKcXhQaH
gMk4JTAdMTEw37kD9GHWfrgeBKlsln5ajIpY9qOF2OMk4LZvmrJzd/kkfgF9GLwPNKvP3NPuvz4z
wXA2EcpF70skw0CM6NyP0GsL/k9A2MsXXIGfN52Cnj9vx/tP5CxQr22n/APu2GuM+gVqgHEkOmLx
tu3HEKVe0CJDgJ6c/NmLI5rrxCDFwFRIvBmMGRtyGWNmQKxmxHHjw40k7q6VI/XUjVcBJqS77nWF
TbvHRJb4cDq8TBVxvzA2xrL3Z/JshGk4NaxdG80KNT74y2xaUipK8DuOyJW32G2ql6AsQ1oqqff9
AYIl/6KbsS8/lDd4effgH2NlP6DIxjtsFO5FIymVvJR/a+KhtUIlHr2OI14dVfkf3LBDL38Gw4B5
95iEiQCyyKEoU/l03d4uKmdKo/POkQOGd06f4lLVVWHbVkahlCV8gCmscTtXbwGg2GTYsmNeAR9p
KaHlLWtGY27A5NWhAVQ+wcCKMAwsKM2FeilFgirOX1fX3DfB+ROmyyixsvzxEGdjVDyCru2AI6zU
wMrEGE8l9dXzZZlLufcRlGoTj3q6iAVd0OJmVufbdN0w4TObBuk5ZW9wd8HzOw/R2fnc0rDk6dDn
BTsW4ldQhSGeNTTYZjk+Gq1+gmz2eLdznkPzIK0fHeh+iWYwqkhlwEKgndWibwkVdQBw1sv4yHe8
2/pa1YMoPscAI3WzZLDUijFQ4Woz2jnXLn7SqcecFTAUWAt3GHPPH7sGfPiUqX3Do7GlIPF1O17R
eELKBvEmAQZx47JSpUxXELg6JRKnQyBZTlsB5wn3Wv63kJ3yJ4G1779tZPpr94U9PupNspj7n9mF
BEAEv5s2mOtV4pWe3SE7ZcrMX0McdBPtiK4fDQ4TvysXHJ/dhKD9J2Wjo+c0hxlRGaHersvmSWZH
2W77zmAxqbnZV9cPf0AYbF3vOa2iaRAOoJZMFXpAvvIBnmSkBWf9EasR3S27/4Kn511GCeGFCtW/
eE+/5Qekn32VRzsVsoNj/iLJ8BSXY/jgHnsVg7eCyz+sXy9K3jLpsGJkjab/AaoGumpCn1uH8uoA
lJALKPYRe0sM9siWhOZCSGDKilX7Rg1A+ObNdt5eXm32IcLmGCEwrYkzSnyLM4fJLl1qXsREkeUR
Nz2KR+xBQzesrGyEBuxjbxXy+S4Xmk4JPk12e/PqI0o7BsXypguyCaCqlyORim93tIJUIvLaDRKS
nMjZ7p1z5I9hov2l0u6Cy7MX7DaquqeSXyBZIyhjwKScm4wi4+Pw3dVv+3WutnNrn9sn+AUy6eeC
OoFgUAUKhgBUAG06DLhUqRm6CHBocWV+C5Wdxw9Nh6mi6NYI8Og/dHM48y3806Y/RZSUuay5Ru8p
gpRzIcAOU8ZiJLNE2v7fRw43J7rWSYKmn4ygkjCC92qK2pBLaY3LLrELR4AYXi1q8WcKTkkqSPmm
uOiiaIZF+IIpytsXwdFcp/5mR3eFY4ISHQgF2MYK6HN5tvgxu6D1zQ3PVfauAnVtlCnDhZ80Q092
ox+NanOmZUJ0Gj+hlY+DfMZE2/DdKdLvLcPXwxa0aH+kEyA/CfpYej7UyBgd6Y2/9H8CqsFRitnC
EkYbRAahHhjUa2nS72htcPcS/kz4OksFk5EIWI07NHlmt0aCuHYl2isIuYidyTbTCJf/lfXoK20L
XEOuj4NAGMyrJ5elKMu14/bcuSaD8efH1E3n83xHJV5v6QokMC40VxsE2nqNr4PeuchwwfkQWtZd
GBBGhqU/WLASTHP0u+Syi2/AMLMMt/ZnwHgnsN1KNnHcigcpGRtyp/vDgVksHsmjXc6hH/4QHqWX
m/YHFG1AKucZ8BJD1irSOceH9USWpXXcgq3sjf+WoKC3Y5X14Rehfk7PwavvT2OCOmbhPncKle4s
ZnNvs80qqPypITOGNWjNentGP2X0/JZGjzqQyC+r8eWM0x0tx3eUmTjmjoVsj4Gomv3AmxJr4nGy
6Yu1UNKhVyz5g9XFSouvqFip9LpaPWuPd2P03OB9BTvUO0Mq8m7hiet3gfTONEgBDYz/vcBW8aF3
i5VCii3K8FVt79UqUJmnpV2V5hBEXvsvWnWLiD0DdujZV7wdg5sp1OAB7+gZ+mMbcj3m2jMJSjao
8z2fqFVy9y0l7nQ2xHoxFXaYU0CNLfmchL66zwXF7aK6xJ7INK9CTZ5iyvlvpsmXUEY0PF/BVgsR
R70RQ1MKcMDh91uXBsDFLcLdI92u4N8Og4+5A2m2g5RAMjuHWj9eoA6WtcK/69Dwk88Nt/OPxU3h
XSKYnb9BPf1uvko2nN/ytUoXg7inobDRacKkygC0YlSaF7MLrHCNmMVRfNkgPn3eNACVaveALOha
Ab3zQF/f8ijEva1aE9I9L9bKG92HSkxYBCTPpDBXmvmA2bzpQjr9GboUXvHzXGgRKRVwVANLW99h
cqV+FIkhwoccTo0f5cNc1RewVqJgzUWdUX0sOtgnxYVFkjlAPmKyHe4TK5QU6hCesSCk+CeGZZVp
RB41+BccOaGjqrdX6g+3Bycfyxzj1PH4BeY6GV0/23qsxjoHvjaAkJfgVCq+1WXq2SCkxcVy+l8O
tyvlY2eBgTc9BqR4sTIstxJEyzASMFj5SS3MeBoxW5g116sdY01MO6pG3JbBAar8CLyZSVkAbTZi
/RAzZcwgdn5sYNegL4aT2bTn1ck7ucCMU2CecjJALGmE4V5754IT7BOpps/0Z2Q+5jNw4h7bWxnQ
PdmU+yzsQ2XSywsmmEpl94tNgKo2EXNsNUCwxWTVA0LTDQe2gfHZcZMGpxN3DMh+42+cS8UsG6Zl
f9sRtC+b3L0cTgNGu6qeKiWv5GROO5tcGzkPU1G1HW+yZtdCby9pU4xQQL3BlDReMi/2X/SCYALz
3hcTiOKiFyFEvA1+9PSfMNbtDGbT55So0wY/hPlT/xP0hpu1umiv6I6QbwyDSduaBGVcdW1qhI8o
vNIj0Jf/Xx4aLHvMeXPMArUBxCeL5Rkl4GJmARc8P8FKo+nV/kZ2Ekj2MoJ6SwZQF31Tl9tkLbu1
LFdujONrdOHXqVZ/fE5FqZVlNshDnWT1VY66ngel3/tgi15bagcBeLF+IziN/KmHltYtQXiyPJrd
O0/6tRNcQ5BazSNejYubICeSZWH7FjROyBOb1BzXEgw2KlN+mHdMfHNGaPVgFdHtfY27kSK4UnQ9
o07FGVveDG4FJe9sptQbXSdRuN50NRemcovyj1KDZNlBwnN5++SEj5BVGD1p4L6eVhtvJtMa3KmC
mrP70pq61G6qGUk9oyGvGENc7HI1dJArnsQ0pl8z0MwhfwaiDIk86IEzXPbcUshnEqEFLAZcZJN8
btRlDftN+rJrxJuCPau3gnVQ8W29awbF8Kz0/BX4rORB6SZpNX9N/KuQrk1Um22thkjYtZkydOze
vVeMOveuITHaY8vu+227m/QcvapHM2gWWatl8VHpfb0W2OQ+85Lh35aQLap35VmI97C7vOBK4GLs
dD4QF9SQysV2ha8jWhHJjwxLppHhfzxXfUnFC8pTC5ipEptjNH+2c0fIz3bcLjdUCX2jZ8mXWrT8
9lV/f3HwtiMnQq92tr4nQ7PC86P80Wgpwo+uD/paBlORnNsqv8UIXVpFpr/MaJgiGP5U4SiKbzy2
ubEAH2uAwabQ62c6z+T1h28qgtz7dMoe0hOlx89Ix/O9uA24JTE/mZOZ84kVgDv4lA/apYx09Mib
ALIqkhEBNFomL4Sp/SGwbSkQCSfBGTcdFOu5L/m4OwfQzWQWqxjotUOufyLN4gnxN5TRW/1eyuHF
pVbq3sZckcaYRxNfVh8pbr4C8x1iL9o+s2aXD2OtprbKKF4FbDtwkT7n2iLrk/WWPQd1tCtBhQip
DPThgUNRYRn1GgXIad0z+YRnZ6p0g737+UyW+xJXUQBADPPpzkgJ7qVqOdiEgzBDYikLd7KkchLs
LSvIMNrvviYLFgn7QSLSnKeSxrHnnWD8k90JM03Tog3rhj5rQuWEUcRjErgmHhjZ50DBpBs2T1k0
hEqmPzpqeRGweWNcQM+DtkdaGTIo6ddcWrG00n45/0xbMPfAphgKHEINbxqE7jyDBzcMF2kUuKpo
126+pyLdxXjJm3oplk+G7SjmGgjuwGVKIle3ZuCWmZ6z/pXNOqte/pF4eoZIx65kAYZj9xyx8SM5
wvVWzEhP1GpvdN7T/63tzxSgHvxBuvZ0zNg0rveuNfhJtNHtcSItCbgWTJ6NhJ3vkH7MyYLxLPaH
X8gfW/3LSadfqb/oh8/mfwJfd+PSCgGcBb2tbQgjqlWxGeLy1oBUz69bcr4Ig4rhBKAljI/6dxnJ
z4p6upfHFePHw4MLkjMuo8hBQn07RmqQVUqnVsHcziff+jxiN+fhfLOUBb1guKl7puZoo0QHxaMy
uyhchMVHmmBhRlZT085rykLaC1MDQnoft3K2UHmqQLZckcT6xIZF9s3IUfaXR1VvbSGhPvZ3Yozr
/DL2QlZk25tjuNhEBtHe5aySZX5cKYeQ5g31OB9MVoUCwUT4FXqrLqEe6VQqDHOP7Cfy3tB8lTsH
0Spbmmd01DEfECCE9BfQcnAgA5JpxkYD5pr0troU6LcuC+G4tYOcB/si7txp5rOM5rL3Rqqe1+Iy
ZvKwkh3DCInfrHoFSVr3w/LT7/BdkPLh2UGNrJQ4QvuuCX78TtWBkzvZTFylZaq3yECou/Qnv950
WPvBaameCLDducSZsveWvHsOFYHF1JI0WlMJRBbVwAd01uIQ2QL73NUvsb0z3s0Q1sPMCpCZxeq0
IV0KZQ4ir+kzIqGmVPPhDzXV4xe1ffSspVLHzGhdb4RPzwQvfKURscWLk9t0wSw5GPU5MdtYL30t
Wca+SwGq8IlsoNp6+BxRrBzMvwMDoZf3HdRWVPz8mok4+AKif2+1BbLmrdKp2nJS3//2RWHRO1b5
kjCzy+JaCRoKcC9vUA2qnrF9Mf7yTM7a1LUDl4o3quzJSK9k19k9cS68iluc78i0oFKfUdMgAhEv
6HyJ+Tq1CVNxpuRyFW0Omf73Z6d+tYzElE9hWV83e4/6D+S8mm3A3fXf63KNGe1M3JXfBVbr99UM
Sbkx8PL6B1l5qVwbw6aDsJmxAUgihisLvYD9c4rN9JxJU9V6bsxTmGI7xtoqsP5DDPa0NNFatTL1
KJa6+QY5PA9hSUDteQJ7Pi2dCw+Ca4PZmUlwT7kAs8hSn8wmBXTsVqKzvip53HihqYFxjlaNJSkF
SQYIqoKN92FBGADu4MQUXyx3bEXj1MplME38I5ujwR04PkNy4a+61k1SKfd1g/VIIJxrdKw1jjOB
Wg1cSV4CZAqGPe0QjSbh5kfgBQKVCyZ0Hxn50BNq5ZigTs6gs+YjITrWiRGPY7M0tTQsbmJVZkU/
pVsKaXu0yADQdhwDbVRBWgzknnrJM2FGkSNhRjQU9trTThzxnjliVsLNXTH6WxunaGhYSJ5LNadP
BTC35a/g+bqSaSe0p9vJk80dePJFLyLOvN4ZUAaUURq1euWHWg8U2Pv6nJDC6zjxIyGYYbSB3viU
8MKQLqEbc9fsw2zvbUVp0ulvrs6j06p908Gw5TfBHMDG9FnecWglOaD7M9b01cnVrFzUOHLbrQaj
k1FTdepMwA7CTBCZvI4wZWIa7qO9f6soG2KWc0WX3HRbCyTx4KdOeWeCJ9Ix1RxpADIv6E56QhYu
cV3FyMbDXpWCF9Pyklj7hHywq/f+lkM0vDr9J817TO4lCavwZZT6aeA2IJvv90vf2HzQ0e4ARXBD
RVqWvvvsVGMSHnhvRNUNp2sMa8L8OC9QGa3OZuDYnwMwV+/iR7uJtKSD3vGVnvIvMaiQ25w0nfQJ
XtWob9c5VmG2ms2Z/n41NgnDP0BLIJb/NIicuC2d2+rkOAx9SqPVRHoCW7MpUvplXjaYNvXpccGQ
pJqHNlDcLaxpdywaBEp0AaWYHiAfLWLruxDZd5pvw5J/gDTxaoHg2Xim/iLSn+f/XMCIG8Z0BL+k
PFOSQeTWmtwt5b0u2bzgbXYqFCXQXRyrf3FdHc87URY+rpsRskRu3p2SxYgWk11uMjCOb+7dpn8e
CBTy7tlRnQjnXd4/ZriUyXMflWQMFXbX8AkobksZQuol0TULmszOKJmx0Lw66gwIwfdM/2ypFDNX
rGinOG8u1isMhsU0y90dS0V6NYp0e70K8KZxxwSGT9BtiOgCkf8Zbjadi9War3pHt8d4GiHs40bb
TcCqylVL5zCBY1/NzBwc0pgNoMfaKYWOe05ralK14PA+cg5voc/rzlZaKXjdYhRXDG6ggGn6FYgR
JCooC7TDQ9yq0RoRtxXj6mvbzuKTV3qJC5HFMSmN1NaDmHVOS6zYEpSlItlOSl7ZcFzpEjgw+ohw
VQkg5ZG8gBY6Tjbx/IeBX0PaWAJ2BMemBwUAh2nJxLxFiyTKhdTnbJOVk1t1nU8eetLqjJD0ONP/
b1z/3WF+XSHyco4jztf67Cop54PQ71GGxKg7MGpItv1+o0M/nHcixtVybKR723KnfVdMu3CQhvlG
i2DjQ0NblGNHij0OveCU81Yh1158fFhwXLn1CdqDXutKII92Dc3dYMMeuDWR8p6UU5E5zcs6Y0AG
lsuCa50kbFceRf9Trbjm2ivQ7v1b1xGThanVOHDbsHcLWOoivGm+5tskF+SvMFv/gjYrrreuSCKl
5hn0cAs0uDkXtnmnqL7+bzeUk9J532YDzy1DgMzdLIhrz5p1LJlqBQ/ICFTqcq3I8Wcy4+oJ6cjb
hqfIR8KAaTZ4FoYvSrjXn9JR/A12vLMZ+YYjtRYbGg5qGjq5IJVbyBuN8RymEEWKX5iS1dOJjNdS
CTAFcV1TX2axfKOAnFCwevZahR4Nzk1HoM8Mccbfe0fcA0TIFpsKZ20MO4jFHHb3MaumDdrizhJE
8PjAVh9MYPpiG1RYjc3DGxH7j2ljnFUMPWSqpHoA0xXr3pkehEUtzNC+533phsOu8xkOoy17a032
w/aHS5USppIRRfYV7IYZVlCCZxJp/On8ss4X/mPu81f0zdfgC4FyMWLs/zvVHjuhitPpdlCAcQfr
ioYUOfhH5Xjzyuc2qDhGzROBHbGKuqHzcpzN/JI0wxFAf2UZhiVcYVF7zMV8wSuy21e38ySmNB50
dzmWopWoZT1sCZTGf28VKnA/pnaPrg+O768kL3CY+bcxie+wxI2mOxF8aQOlhvOjve8RSsdSQa/5
Bi/gQnUO2PsYK4mS5D4+FxbraIdvc4JnBCDC3GrrZHLMhbop53rIR/poSoxTTMM39P49gIB3F9q6
2Rg5yH5JnecsU3Q56k3sJGG62rihim0A388u7NY8r40JxU0jxAz/cl67TDqxh+5k1k8HMOqJiLBp
XS550xRpbWz+9eluCPMAjakV2/P6OwwcGm7sb1Bu4i5jaZhoPHALmONQc0cBOy1RNGlFz7von0Br
H8holXeNYcDjFSjcl1c5YkEgCgaroWZ7O6CUp/PfTkErmIYk6RQtV5rc4rYA6iWZpbK64tVuEfGA
qWd9UDwmIf6Ll5y/reFj7NTROma+KIZh34x6nqkqJ4gRkzjA7vI7IHAiX65Nonw4Nbc5/8zUWZqR
bfpwVCsAs5KvyxZ4t+1QRYuF5My293usjoWf67wj5v4IcmrNVQIuAn4y6oOipwHkMWOveuoW3wSM
K59oPYHO7kuWQ+R6cWCcY2Nzfg7q+tKQVvMMiRcbSQxI/u979niMDOh4tfJIixlm5Mv3GFSxHL9j
xphLh11In3lJuGGj9cOhYt5iWWro+y0ZHj9EHpqjVm0L5eNzIVmVpm4C0eZ0LOmHLav4vzlB/7+R
kNbroOYJS4L0wfe5TzR1Z8EhK+eg0Fh0fQBhdTfkAwThBxZUhwv7vGRAf6Ixy30ySIiu+oKnXLJi
XmoNugLguVTxQDyDGn+V+/eeTR6WKIIWsD339u+PlH54DT3ThPWJ6hstagBDFdzp4GphE64EfZjs
tFzmboBrOvyqQT+9U59kz0DtpP9hg4grDR6WkK9T31vw6TQ6CjYrxctanhKaBpO2O+5qyShRxDUd
RAAujf45s6QdAw44E6sL9T7UhgxBBlBD7lYqN3lW99ulWc3wdfp177Xnv17hdKN5DIH7u/kBH4FF
Zap5NrBoCrk/1O2IixyBG85n50asWO9DuXSlZudUkHX8jSUwUHw0G40+g6r6Wc2P7j1KoZYISR08
U8u7LaSsHpWvNf5RFo0R/d+DUcyayZh1EveyYCGtqpj0Wn6n2T9OL8KJRlyrQOPghqdgaP+bGJOL
wb1tT5dhBgsa0e37la+7lL/MnmE02lWRwyosJhADxcCShFEntsJCUdNAzuEkI+kWKyhAfz39Ur2q
9wvDgDNl6u6XwVEFpxMVMt9yZuepTcd+1XGjFkSlukYl8lmlCqgLA9az433Vg2bZku7PIRl80mlG
lTbXlR+Bx+N2V2VJVhONyeaU01JHYaLxHpVACYr7uvG62oF07BwuGpx0tSbtk6IZ01Cub7/65WAY
nwpIRhvtxN74WlaXmsXublqxMNmu156i25OzZWNYb3CGytNoL6QZwqRXVNI5yQDkti7Q+Klu5pms
QIVC7Iv1Bv7Q8vFGI1wE3UkolTUTmf29TIBwYpZuaPngcGrP1jwthjGpB1mdL/1wqVvS31wiboaZ
3WtDfsTmKidT4AQqeFyMioaooseczbcx1kntmN1ZMX6lTkCQTzsu1mffBSbXfIP9OZcQA5R8HroP
lCvSLFBZv4iGRq40uwkGBYlYUXXB/XKUx2O6pJJpjgLPCWHr6feCsGwRskYK8jiLGGfG6P9QKXlC
gRh0H200E48KwWBA3/HhDTuE6rmudg/gW0n8uCwsFT8Z3TaImoiJGzUcZvAf2P6lCoiRL0U6x+ba
SSxnMTVqUrH5Ob13pi8fnid9CzhnlaN7O/ChmuFLY/SfFAhako7S47p9VeMzNm5GYzOM79kHq1cY
kwjTKwq0sMXhrtUwvX2LRMsTeI9Dhmn7wFY1R/h2eb7AkzgnR1B0Ma/5fYzyILLxtY31npoNiq+E
cldSAPR5gCh480mYYsdN0hN/2QZsEd+OXXkBpO6qYtGLonhcf7y99ZVbYICozFG7dDFUM6MM1eTJ
2o2Lzumm6Dn/4snBNcvUNKJdlQ3YkKlf71ZfhEGSBy6v6wLZwuzQjMTfNMz9xgBRHr5z7TRvPduG
zLDQYzdQQiaGzd5+XE5xnAgKVym1RMNkO7IMKXVkzoWSCAzxUDNR8UjsYvp2QEevDbryqd1F61sE
NXfyP90+VoxaoCWKhKZCuilitdKrwM54mE+LciSiKXN0t0qv975OEBrpI359m7jDczSzI8lF9FpX
LDzxE6+9EWUwgCu8Fpf8vhCnZIZKc0VuUO/eqiUTFR+AW0GCpGX+UurN6JMj7FCijFluXaV/PXcq
uyywc4T1jz9wQcljJfPiBsPRxfyufbrKBZ6JgQ5CrJ9ZxUgC4VLau3qW6DwMS1au3MKRw0y2+MDe
s8z8TI97XZgxXgnFu08NOKz6eNFWKKyvy/gsB3yXcrjkyNWEw5bg167QwjhrmcPdwf47HGuMaROE
qhGs6Uk0LiElVnICPXZqzxAWQ1bXGavrvDJZ3fNezoPYrxGT0s20cGfuk/4iwUQlVyxFFMty9O/1
gB2NWbiNYboqpp74aYVykh2ebZ5vbNVROEUd3XDEZEFPPB967PG1p3QrJ/wENL5LGwBUqxBed98/
cLRqZLF0g361T4zJYBGmM0f5NZel7IcI70hEfIKW0ymilEf4686KPNihEfbe2uFGB3nJNzNgR4Ba
QwhxWYLtty5AH0dRqFI+qJKyr6W+9jiGAJalG0LdDnyfQ/TDG42D0hwiO+Tot5JGlhc7G3GRj4tc
rMhuCAOK4jQ/KkgqwIn2p8ef8Olg+2L6cZX1ZUTFd3Msj63i3zWhgEKsdnJdnlbmx31rIir5wY3w
CzaEtAHwK1jvMf2+LjU8s8qkTRnVozRR6ItVIaBHBsEXnFVQmsbwiLLZ8eE+fwssuG2m5xWKXixc
JHFb51TJ0oFSfCiy/lVpVDivpFbPmudfWEHqKt/xQ5AFa1TItajffOUnHxpmN8arI1dNYE2eyso8
Qv4KkX9ZVKmj7bmUOPgzkegwHVngaUzoSbSx47oPYm8tNBhcsVqHf3f16AgI5iN8jJYpGJEPOfvk
tMfBqwUZss/2ZTkYXesT7x7z03An2WIj2rLUvr/NmlKXiXkKMxAZJRDBxDy+75MrEKFFafOy+IUz
kfIwKnWFfvcRAA2Ht5Bi2thtQytEo+mutcgjVgJPWxp/1Kkcq+c6IWNeyJr5f6SrpTvfTyaa6Vvk
67U7AWiF5TskxeQokiSf2ja/IQQbfRas7giYTxddbGYwJUG2POah/g+0QRxum+U1T6bIT+8V8QKN
gHO1xujGZ83FwPf6Xci9JPD3oOJN4SGydhfVkudIVUgPHlJO69jlu8x24sjD5+8ynYO4G7Efmw+9
y74dJ+aJLvLjvsDOqjveGMMFUkkItBRvgbIHYrb6IrWDGWEe+jcubJya2464NlYClTAUeVebFYh9
6s3aEYZEFYZjji+iFv9dBg47PO2abGhhs7ccMlq2AUW478lvAjZLoV7ZP6Y9V6CSk8Qr7B+S/VMQ
EvX08Tlq4uFAKMhJYm8rWOyKaNh7kKoxQSwksPCMD8mzgLittXZoh/yc/fzZAr/IvrwM4TN0SWnf
Rs983vPVVXZt0yZuBASwUR+YAZVbcpmt37TSxz1bMlCIjEGgGnqMOraYx//aJ1RYlkfOE8qeI6ds
KWaPlXnxwR/C7B0RmLIynHkTpzTQcdWtLpemrsyzZIMLQlx7y4DFs9Dmq/V05Sr8xw8Z0y+oBKlX
eofaP84I/VVNjFE0DuCORqV1svdI1oyuj7NJd151e0VTR4ujC7mpalTNl2XYEWP8CkeajAgpf16x
aQI1BOO75dxqnnh+Z3X1PV70QuPNtH+ylwPBnt20/UQgmuZWPYtUR3h3rV+uY/ls5U/d2qyvd1YZ
FOmiCxUUw+pHdSMhgIELmkoJcML1/ERxS93whLzMFSLJpwzrGYOUlt/4P872VliAtNGpOfrDo9NG
msIixrAxk2HEvo96QChxeapFTMZ/HLWPQ24Naw5Zy9heRvzOONvInYQpMmLcvLBRojdLQ97G9j2t
y83tLW8NdR/PMZooN+3BQgg3FURdMQrMPOqq0kLubPPOaAhsTs35ME7yc6bVZfWkTDWsTPA7QSxS
EtYSCWiUkEdN4Lxdk4N47gFD0fbXNNdBzklG3/c1Y5Y1KikNPs/C0Qk6s8hIsT5x9LVV1p61Xu6i
iNvbdLqi43KOZ32o+zsZdKSVXyrhTuiFuKd0oZ9kG60Y4ysdpz+xKYaa9juuM+jzzO6X+qlvC7nW
ToruS2Dixi1h0V1us/0flF4oK6Yj+ksc/ES8RHHy7aLG4V0MoegDRdnvFTXPWtBzycXwXi/WUZYY
BuE+YaL7t9R6gTOqE7ErFsX7lYMJtqPAU4EI+RH+M4nvFFph6q47sk9Fl2qdVhdi8LXx6e+484lZ
loZHHnwf6vBFC5OWuLhLWr6pVUYdZJUc09Xjx/amhXdsrgJ0TZXZd+pgWyrjQibs1soDJAQH7ydI
yRRp6jXAW/H69/M5HbVZYBeLP53D2dzr2kVIFsUa8swtZtIpHRoZVQFUpZci9gunDdCQEXNpx8fh
Wc0p5pQ3kMSZTJWK+lQkq/J4q4wLBUPWn9n5TvAyNtu6j68JV3vK7QwfEfCuiAFo1ZOxybPUqXC0
2oGrKp8qZQVuGx+P8S2DG/v///qpMtB3qSUfxTYmUibnxFmdxaJ3JxOH3VmSNgJM+JWL2rdwIJZK
yHe5hLUDFt0PEiKV7GfXwv8dADIn54e1kvEG32d91ZhWjn9ep+uTEEr3bIKPHNYS7uXsgKY/RCkR
Erk56BpQYcNYISIf634z+9MH/orB+a40KcLqaWo4HAstAT63po2p06STL2mIpYxefm4Yb+Rbq4lm
bmLFpafqW8cy3LpdKLT9iSIQ1OQ3sgGU6zvth7YGkoAGqLg65t/+rNogr+owxus78/EFe6xmFu3E
AfKigWexOKVJl/t8CwEe0s9QYNT6MfqJaMuUZkhZkC2BigrzsHgenLvr+Cw8e9EKrVYOCE52v1c0
7dj5IUxihibi2L2Dp0Ned0AFXBub7UNrwCPaK7HJgAJYxQpe3cdHYKaNJfXIA7198j5Kdn1vpvIq
EhHp4/JShY4sKryfyJKn6+iEyPCSaCo4b2yMI6eaSlvWWwwcQTRAqlphAzbBTH9Mw0PlwTtptVqY
oDTJZ5xtMNj4A2c+/vYxmEc5GGCKznfamMpvXRG944/9lBMNlvQPEbeB6UxOE/z7KBOdxAEFaHBq
7ecM3qMIs7LfOSdVnMy3OiR0Swl/xAFRiE5GdZoGLdThokzk9eY4SOG6KZm4B1GaMk3KtlOhYfuL
E5DXVLqHZKJBM4YYKLxbou+iTzcppSi38W/BCibd6s87hUURhKfVmqkT38W2KLY7HOmS6uDT7fNX
gLB8YK7DXseJP9FtKhM8mvG9P0ppDsoWf6EB1/AOipc7pkgfK3IaWJWk/Mb/BkYhI7ie7D5j+Iu5
o2Fg6qk53TdV/M8/hiVJC6EzT7YVm92NJPL4gsmRDJeQgtIemCiDKrYQ2hDsNNONRRq3+nR713+D
J40IfZosSfe6FD2Wv7hW9sQRAgpt2l4JPFptavKYuxzOZtndzKjnQZhppYWApeWkn5hykYzgdcdU
keUjDr+OXUrtncNW1vt83YI02x9xC5/y8371GV5/yBYK3mrYyJCPfW/fPzq+MoPUUfRRLUHZtFc8
7aJnv/vDr7yIwsYy5fgNAX9TNpksOBtcSd9OjLqjFIMNo3czyccktkDgDXJE26FbuOM1DFjaVlrD
fxqqtHF95942fW2UMWoNiuFBdAiZU2pQ8NQHbpDvUSTJEq9J0UsDr1WNdElJEnexITGj4COweM11
gnOAL1fTuCxzoWnac95zxa3dLTZd7fJkSHsi4k9i6AsWLp2+eNBzujhcURM+zp4I5SYNwZ5JxbKP
EnfUdBEaEU4OBRHVkKjg8gJvvPELssUipJc66DCQSlEIzFq213GbH6HIEytXbbnaCh9SnP/jAY3a
XVffUqBUihEzzwfi3nqhrz2Aurq94ItcIW33t5G4jqcdS9BoGgWaabryLpJn9kS8BbOGnFFJOC6k
cIe1vP9G/mjMINBFIHJ5LqUeP8Jz13Q6rVEbGxIb33xHuwjiYfv965m4ThvB+MbmX0a61xt8/wsI
Ma1CO2LAIbKQxn5nqfZ6ZHUP3P2CBWqQEL9yieAhomKlXWJwQqa2/HBA5TlOYKGkYqKdqbr5jx5o
Vaa+NrHvwLd/Pbbws0ggDRId1qd3/NIttRH81PaxkQz78SWgjp5x8fkEfs+LzUS9E9K8S6ZmUVPc
5HfK4jzRmKiwzMg6tCv0r67pxOQOSP09gvLtf/yaTNpLVG+9dOYdpLHe9zs+r4Oofgh4P1KamX/S
GdRrA50z2Nai4Dp2mPQVV16IBsHjJ89zS4IB9LxEVpAWyMXINakxpjDopR9pMN7cSXemzbz9eNzz
6JzjS3vrIsm6KIUPHMpWZu6TP+0PWIjR0+10uv6Vom4slmBlxp63xgcofH/OFrdDgYg5nWUwgC2X
T5kI31B2XL0YZADnuL/4n+JfelLio9JoC9OHePL0S/gGhIKhQPXsXPCAM/zTHh3ZsWgSA0Zu4z61
L+kkaG3DFAeSQtqQoIhe0RubtuEaaP6Rn6KHAgrLYoSC5jo2KFYc9jawLCJRjJOrr+KClRGfiWhG
CIxVTGuUqlGDGrDeUJJkIXfo564sRn9XeAmNWkI82HW0My09xQy1QP0kjKCrA8eFvAqHYdvgnBAD
1+YGVcsr5Hl5QrjqdPp5OAu91wRBzvcAY8aRJGd/3Q7e258ZJ8YbdC9pWsmqEgVzUyFhmfcZGCc7
iGUKHNCcNym2Ge8Ck5rNDmshnolntswKvy2T9V62HVxSZsm5hWo3WD1tQonS/ucwfPYYQBGcMFAI
VKDIfuml1kR/JKIaTH/TCfqt6PkHHe2iNJyXJgRQbHn8RFZZakTrBBPwjnwc2ssXJbxuKll0/rBK
wzC+41KhBhKG8udWG+Zc9ouEZsUpaPRGfSVHwGC1yQhtDDp6IXv+2RRy2he26zc1e/ld8HSMhhKP
n2n/LCFNQOJ975XNAhlHAIz0VlF32iTlFHnXzF97AJLxaew8yKlj/JvuBGNAizPnUaceo4ouKiKR
SL2y9fdSYl4dyOoM8ABZQMdIY91OaL5b1uQaVVx+0Ok5qmx+hIXcicLPHjn2tErlCH5Xn0xeqvKS
E1IYrMH1DCZQnu+T1ylIificwjkAjyJ+9EQ1H5/+i6OUHENF984p1WqrMRPvrjpbVDoGKy5pCHFK
8AXHXcxgwiNq71mGzWJRqWhjS7HwDNJvQHSd4h4+UJQ/nhLIDXwARxCsBpBnUJs+ShAzaCWYUDUD
dax86IShNprNAhT4tdNA+i4G628Ss+vAfxtMTcHxgL8VOm03ptbxZ/5BvedZHsYlCT7cyUWlogMt
MCMNkrc6Fmc4lGn15VXp2/uIVShoT6B45BsE5ED0/6lnSscvjOLDlJGj38b3+4gWnZbz1TCE8Czy
rZolrbTWhLZ+doYaiNi/r1P3lVe9oSWBaNc2EDKQYZtg5GgtNUFs+egXTk+M0xIfLLZRuMRFKt3Q
+a3w+OjmJLhyMlDYsieQNTcGKMEW8vUnHyD9HQa7uZhBP/hWogUkTUajb50DpR4SKEn0zJ4C5Gov
Yz8TXXk+mN/9fMD8K4YQmw7YfRNFPWtEMyMYjmkGWo3Ez0+g2jNH7CDkkb2T36ljHkkxT4KliT1s
OBPJl4Z+Bkxn0h6ZC4s8VCHTGBnkiCL5SB0gMs2xAA7HxqQZGGJFpXwhuYhureIXoELhdupIZjPZ
T+/JRuCiWuYKq+jmYxyIMgS316aXzmnoFYKz0pIoL4dYvDX2F0SEHg08cPW0JAS9kZIlXj60sEwB
ocx2lMQHwz5bE367TBRbrRTUDu36oMtNvXCRKgFvclRsqbQqeGFtWA5oDB2X1fEk5fh/W4nw9EKG
xoWuogdimUjof8J4nX6qsZaBUlKw+l+OwTJ1Gwg5y2TmYQoGesyE9PDzf09zSn4CsEpEgYbyyIlV
q0EIm/YMgestv6MXSqqwi7PCcdkZA7K1UKhTOhgzwVju8V2xZJeEDwwVecRe8YhTbLZcadq5gmkP
eB9pxoPvC5+BkUC9C8rK5iT96RMyMMmO4sQ3gLUEizZQUEEHOhZFCv97A1NL0QV2/e0CK/AXsrlN
HO8ELRQSnXtJUoBgomIys7KDQTt4ENammM5LCYi3IxDXwNfILdiBrsFSgXC5e1k6XAokfXwhdYB+
enreKni5FTnYMz+JJz54Jt3+642Q3duQ32EcrxD8XHgKVCwksKgYj94wHXJsn6XVkPww3CuTsPjv
50aC0ZeOe4zPl4ZdBOx5mdFVljZCZuNS1tyyVJowb+CZw7ncSu/YeMyjYK0733VSG7cxI0zBJ3qU
zKlqG3CryEJ4BsW52b95eoiX1gc4Wu+RdEzEss5/g7K3sgUbZS6U0czJ5FMPJqsf5403ANSsmc9n
kumFYfGeqANUwoBisUIk9KZpofjzSrf8LZWIkp6XnAuUJUO2SmMDVR77GNmNQejjytSEY4wjHAUu
1nIas+qnTamblIQoqVDODYXmkqnsBcMs0rIX7pa/Cx8tQuzMnM+Q1ZZ8tKQbZqH2KJ5rhrlyj/Pw
DJLb8PkDRqqEmGAYhfFlfE5Tae0LK3Rm3QvY3vLUqDD3k5wWirTZgk+AwWRSO+wRRrjUZov78XXW
RHLmbHTte3P7HRweInKfryrFQFfWdMHtGLrPfSL6jFQTfrSRsQX6wCSnzaWM+U4MjGWiQk9GO+x+
LcRPBKr0qdo7d/7tsiP5V6Us+ClshhNBouj7ij77VTPqELciHHbDGfTCI9fp4OJQW1fxhG1dOgl+
axPuUyeV2yGfRYRDSSFHeeKpuzyQBQ/btrvmHEzBKpjew4g1SmLCL5fvdXQSmpY7Xr9Wwdm5QmB2
1U78aZMg1/In0uAzK+yIbb+tcWjCE+7w5ZtokzkTF7oTTAPRXfohyNJkjyJQyZHLGyCf86tlM/g5
5O0s5OmXMiDyhz3ex8gGfviShspE5aptAiGn6j3UjUaVuw3EvS4kSra6l6QVzXwKVaB8Xc4Z9EXr
dP1suuKbaF2mgXHS4m9VjWy7eB4r413z7sEHZ8la3kRsN9DRKQMAb+pzcaXQml6WKsGmwvsg6eMj
kFHPhN1Wj0rxOLfiv81weyJK+HMfOh6YjTZY71MvxsxPxP2i36UKE30+IvO7ZluujBexkD6pe8LH
iz1Aa+qF1BXVvoujWe6m75mToDkSIZhDtbQPTuSb7v6Unq0cC4h6b/kkRiy4WJPNhA7rbMpJHK6G
1Aut0+V4OKsxT+qnEEaQBuk7tlbk8D4BgRu3GK4sPwr/h5vi5S/wpG9TPca1wdDpI2uE5Ilne3Xk
E8WHKEspOpuGtovZ9jkbCu8NrIsvAPWnVc+P+oWY7tjbt52AejxsuI8kUUQiRUivlzIWEdo8oIhj
nmvVJqMolx6QSEtHYppMF1ticLy8Q4fIf1tgKUQSogX+CiH+YqYyJuHHTIqv9OXfaTDE+ZhQhipg
UFquNprmGes4IAZuargsgcWD3GZS2y/2PbGc/m47jdQnJw9NdQs1iGqHJruJMzCZrXloZSRi98C5
+1nOHgfhUodytEBNBJkKb7LwVEV/R6jNnkWv528LarqyJShB0+EaDDrKdWFWz0/nWrHu9j3bXE1l
SiwT6XqUUDOsNTaCTYk7GsO8CxFNnhwEIXiuaTIho8wtWZgQkuJXQ+B8/79iM/Q69j2w+IXPbNP5
Z3poJSBu8162ShcSFhaI940NckqvH7CL8KrJ7E2LrdcyjsEfYKXB1auC25axTIQQFgpLJ9QTSlGy
g0vtx6s+4ZTQuRlmiEYfbGobNAjulj73Jz1yMrGyuffnoRBQsOm9QsAEqy3KVnmTYgGACPKCJDHz
C9Y0EmlNP6C4OAr9bLT1rZwfmdo9SeTCuKJ6MAeAY9eEZk53AfjjDS+kQwSyD619C+7B3VR0eSTo
wD2ULrp0xkxoWMVSiac/z33x1+vMp+3MDJ4mpPvqJuVjoyjhgCpxb6+yzW5LpVgWTZEoW7FodFD3
sPlMvoWAOkRYfg9ilkHV8uran4dxF2ElIdJ1SPpZP8s4pDMFtl4h+nFx1u3xFB9sabwzHQq0mM6n
dd2cwPDDaLz2BMgYe6K7FuQ22dkVDKyjcte4WZRqFZV56biQjPnaoOctDCXBKXEYhA9H/I4pM+lF
dW4q5BhkaAq56chYeOZPyMWIk+0z1ryouZOsIgj5cgNiAcjxrr9OiYbth56qgCvYVf/Vor8PSnKl
eKqK+O2eWaF1murfvr0NrKb2C7sOPbMXcMJuwnmNPUVbf3BFV4FnHNkby0qCQVxLG0vcHaOcilpo
HYnGTmIDyzbTrhlFH/6wNexoEEyG/KEyS7viqXoReTR1tojwL9zIWmoM3m9aae/9m9N2oC6RqCWa
tyMnXpxWvqIkLSCqZAwAKWHCuXXI1LY6hfVg0d2hDsxQfyyExuzrPO0V1PV4gIcDv5uaOpbNFAlk
etV+oA/EZqMYlVWCD6vS6bigYDKWQUTFvdmbYnsXYrnQTFN47suFO9nn6+gb8x5dAq96hXfWYmpE
cdOI7p+kI0C8I3aOZ2Jz0NhwyRnlqhVwcQpRpVzYTGtmoVfscwJcA2In8EBOPu/Uiv2QgrAWX4mE
1SlNL0ZboskT11fsYHBvAQ7ddvnXstohutLiS+yLA8gvb2A7pFAtOfwomNs9LQzzKc8AMGNNo16p
zlSYmzg2inuQMn2d8j8T8yY3iBMS1n5ZPHkpMXW54vMHEL0uoi0Q5PFvPGQrRnArxcKrgU61zS4h
xz8HvG4FeLrjU+iD4QEyHuIPFhNcbXDMlz9nj80A7gkSuL1bw35xrmxK4VF8+8r+pVLMJOphjnty
93+W6sr37ZbzUsXw2IQCMzfCN6E2BIdEdGgvrdXIOGkFbK2rcKFIXu3vCmmEOHI+PQnwVNzbOZ97
GXGeTb/qKewSyJ6lDZgKCkVuRUPiF1voKIqezL4IXgbZlBDDWTNcXoBt0emiStUWmu2hRXsW3wR5
+C4c48YQg5xFKPhtl39sWz3X8J8G2tSGNwfsMGa9KeFI3C+nUPpBSgcOLWe5ICtqRhIIg1G12NYr
UIdSs+cUf1eIBxLrWyawmb4ZgHZwH1NL3qjpRADPyBjyVK230xGiOqND9fcKRWG9KHyeEbwyV13e
56COqr8C2CdGoSpo49L+BQDEpM97J8m+0td1M3fMSKccynGuBJgDFabbiB1QGVv8gDVfApGmNObo
YEyk+NuZO2bH/ZSb1lJyLrOVAS1KOb60GYzinKJwT4eHP4mnU0BsCJFhBpbTzh8kaE86NFVA1E/d
zK9vGfnRZ4hIcad5wLnAHTjRHjxWtVIRPDZWSCTad2ZIqDdtSTnL+6mEAwQ/i5yU1QRsnedRY63+
Ge+lu8dmI9OtPkurZEbVYVEn/dNWSb3NO85LGxHKvwj87zsHoU6u/F9/BgOF6LWG+CwqM6qFhque
iZrFqqRyGnkz1+vSlIln+IjKMmiTlb9xzKl0QLoA4jBDwZF14CBoCiQfAbZpJ5WTh2EZ6vupguM7
cG5BNa5Hb1dy2HOmQ4lbMpV3KKbDBfV5axzo2Qsj5DPTn0uwNYkIlXsgLdIX5LgUROZS1YPBh6da
ZGJCaq+24vwitJCjbdBetl4bg9+gY67ZiuZhO+EOpRZYKDkGG0+QNrAtd2TNUl3ci/o+qQweBEE1
TFt6TxGNVN4SbhtEt2NXORSdXoeRjB/Z277MCdCDmSnJRNTW8N+4XzcEdkIy+eKpaYg1KFF0FqGJ
PZ4E+Ghsaa6vGPVPoSDlOzqeAEKf/CsXi9Hk5gUIprP7+K46xZ1pjrAS3GFYE88LXrECUCUNEaiA
u8EbrWouCuAHTZIn5kRmXWk1ATiSHseezp0lDkfEx/Ctuyct/w/SeZTU36nGio///hBSUwlbO9d2
ccBTaOFsS2gqU027wYsAw2KLijkB9xhyqGRXNhBWcyrCVkNeDmjbkAKcVpuWdlsVlIAEgbyIhitH
CnrtYOtxrz2EoSRJb3ZMSkAkDY0LAodBtBc+/AKdIN2bYT+7ziIZtbexp8VlQ4/Fykw/g32L81Vg
1qB2VX3lwwke8Gztih+JlCFeShGbw9jpBHHLAHnw8K5R47jvEVRgyzMh8sqS3xxQrHhXCieO80wV
NbCyh/1D5A8uPDGMhgtqawQ+At8eOvM30nuEoiOUaPPkN7dtHAwHxtqb84f9nVHGmXt1hMU1Wa42
wsv5prtJDJKsxBflKqxNpYQSKMfbx0hGbAa64mpkaWUw8NZFA512V8c9U4SPnvIytE/jvZ84ozkx
qFp/f0q+0DMz0DBwaBt7gp3BmcgRxWxmjvlDYFk5ws3Qo1T6nR93OZokJGrW757ZS4BuoxgPrUqw
qZXTN8sOwEql+3RO1GKUYgRtZj3j2iQnvvsyTOTMIsrshPVX8j9XTFNT2IUOsabb5tNIQG8C5XFB
eK7W5WHZPsgJ/DSqOgbyiQBB98B3eoP5IktQAsBZv2fVWTd7F8f30fwiYnFb2FX8xef1ET20mn7C
XnhbCZXo+NAQ9Cy+6KT6UrInp7Js8I5xggZ/lycFdyUouYE5nU7mq2TEXLFk/Ub5c/FqONSiu64c
Hogm3MrdaCUZHLZNKDwv/VVPeqyVLa0agMSXBEAkjCeAH32O0SG9Tbi7QnSFvUglXZr88dxJv0wN
4vCZmGxtEG2Kj6qg4qqs5gA1w6dlym2whPXmDleO6GnwcbODPSsJK3KKc7qaEr0ZecG8uxQLwmpq
6DZhKm+IHdDtzmhDmwRkAMYjRC3unfay7XGlB8viKxSLUlR/AwXfnH30R7nF6azqjcnaXuIQbDzQ
Oe/MRAN+zz7ljdte5wIwR4SvLAruTyxlEaF+PeOrZma2VeEOqiF5opoYDP1m9PM5W1tpfGLZ0TZX
8rTmwQKQeLc3hDeR8+HhqnGR/IGgZBEc5Cph1R2Lwlo0YRwOC6j/dEiuwyGuU0HC1kpDUZwztm9F
puT21fzCqoqmWCDl43LRyuz5Xs2g9jciffYjIW/OCYM9gmFSbyEtznCmCFHTCJmPy3h+9K/9KHpH
grlhv5HDkjfReLwqPjh9lHgxHbxl/lnj4/i5hVEUql+xJOojeBhTPnkEms8dFZq0atkoBdcPyPQu
BmgSaPucQpBnRC6KVxlWpsdR3tMrLAaEzS5kfauMTrVXRQXltdHHI0huJLXvF6J69oqyfu7Og+zT
nUmjSFUJtWgKQ/Id5qKy4JFZcEyZ2X6IcUoyP9mW3rWmfcp0yffGtRSPbRCsTh4R2Cbiv4qKRgtY
+typeEFktQOtNM8Ghn91FnKzHirQdtbXTt2BWEC6ir6QrCfzbfDdEqvkBJRN7JLfYRqq/3uyHp0K
rAFnOOM4UGvtN3eFgNL1Sfm5HndVWvZJ+LIOoGXSAEKhn6ZNYBXukT+mvrENQszEYlBQbKeWWD5G
szIf9WYgWaDEwOekVA0MfGEUSVTj7WD7YD/KHis3Xh4Easf7NNHE/iM8iaXmcduNUKT4aKae03W/
T7zDA5j+nRqc/jgsE7VkLeaKOEZ9AS84yFrZsI1EZcsqdqJXsgh9Jro1KgEMtngeuSDRZUwpV5by
kvWvZi7TU7NRhImdFQoiClpAODYNGxjznjdX4++8/QzaP6QX6lQRJ8rIWKYBc/IDuKUBb/d7R6/8
hKe9eTtEWYWgm96DCu1PxuQTUDfhgeIjfDZvivHFfADW7PAupcTTvgKdFDRHjnaEEv0wgsuMhBcP
piWkliGmmLi2GQfIKl/e6s1MnXeIOGcN4YLnfkT3O82SLmFoLwc7FvNL5iaqzfXFj2u3vFftPfM7
epwjj4EGzTJ0OL0zoW2/fSSJYXsoxlM3BVTEazCDvnSEqLIOW2Dl7hH5jAiJXP0KDOvpLC1Uw/2I
L6tv4yKxvrvc2kAZuctNLeqOu83sRgEYl2Ca0PsjeL0Vjhir9coAA3lep3sJ1CiRGKsNhozi4E2J
zTrCKDd7m5pbuUjyBBkLb8RoX1u0er3sIt34aDtqRFf0I4E1nkI22IKJtd2tm/fARaGtYN4R80bT
+Sf36QAaTRYveiZwZjv/p172wNuVddX/LWJ/i5/EhOvP2A/HqqqtEtAJ51SiFqiR0wQtwRsMhIYf
AjwVZg3cLR+7BPzD/jx6x04qQ+rIuoQSZhQ2t8fmrmcKxQ7l/4KZSa099xqg8XPptVikQRxfAFnv
sNMzZ9/qzvdDhQUhmmHmmt6U5tAHT2iox5ojt7epPMiWSCp+gM9hB+Uo89hHKcuPdtdn0pff2roz
oOa4ND5XI+EupYr5Z03RQG5Rar6awwWEUiSf4QMrD7qmsmUqO+gOigegG5DMvq9+uzQh1oxzpf3W
BOcomiS+279MYaOYmyl7Pg9zhqTcA/oVzcSWu22xPA0ErC5lTUoeUnF1ayw8+hramBtqnwwW2alp
495f15j07bmvmuXEX9XCXXwsNtrm+D42B1lPr8ytIkzfCSY1nsyVXH8P2qk/DsDrPhzpj/MCxVxL
njmLe7zpd15/BlVwCGB0ibQxXy1VQBz38D4surutj0KyqufQIoQ5FDuJYOttYUuFPskPJnXw4b6w
n5w2G4NyD/qpZT3TDPSQN3obQse+oZcHIhBP46sDIeV8iRUia4K61bp9YdhR3lGq+OCTdLz4FhWM
JdlpDqbY6bC5i41QL3QeSpvMrwn0btnDD89AWcyUYyRe/U8e6gk+MY1C7orSIV2mSaiYRWLcAYOc
l4MkHTJNxMiCZvskUuWHSmJSQoUenw88Aba4rlId4MkXtRd8u6OlPdgjMt14yAbX8U9M4FaUWgtC
MVh0lfN3ikWoVz3xqL408ZiZsNBmlpRrrAEHel5D8ssAu/rL+2DdjeGcFofCizjuvJCwDHa3kXQo
bn1DYrwp8lgkWNbCBR9aVK/Vv9qoTcn+hLFqwTj7CRwag/lSmAfpCalWZM0B2bYvcint5HtOKEDK
vS8RJYVc6CkWvr7yf8YeUZ/IQ4O6gyYB3C1iY3ahCUSKleemAZq7Mt4bs2OeDrqGyGXnHWXnBajD
qsszBG/zqS/s83D2TIIfnKC9COnBssmSTWRmCces3A6QbPvdWKUJOYf0j0aDi7c4eXcNqn85LNrw
38saokKFtSEMiUAJoWPSt2bpzDWaLT0EJThikQEdmjuSKF1ZlhRVRdmsupman3kOcQyvG7rSsbZc
JCflIRIeWx8IhaMHkA74O6hH0BbSDZ/l94Ffx9TJafQixyLcJ4+RMGNlozczYmEuGm2T+K60T+iw
X82w4utShWyGPGwrLYCY+dAUseJUgNKbWeW3rANOVaOlUDdVUThvWAVICMwz66CxLgtEp7pZoZUb
TySiQNeATtmQYJ6NMpxkat+Lk8Iu9U5dM8lOKeJSzyYwsxC3jDOgz4qOiUAkVaGl4Bfx+mIlBort
TVQU2rW/6jdz6qRmEVNwf1zQtxZrzkU6YLq+ReqWrOzmzX0VXdCkMaDliLGaOcSQoXAJvw32OmU4
7O7LwF7F7MuX25EqyyIeKBlgFmSC1IToEqq0WBOKhZp1ucL1jvLtqXtBMiUYfY51YHzRSQGU8Elo
uJaTHurMwdh3rzKyTtwv+wyb9wi3me67hF696vslIdZhT8fh5dbxG0XGpblgppox6nMdzwROyaYh
kZ5a/q2gplENyoBfIvwEKfi3TJqFzcLwl2yOhmaF/EWbLxy8xiHMO041/7qxDyxoaNOsS/UeiB3q
OIDah9a4ggFmCHHpfH/Xy7qzVbJzUJY3jhlD+zM7BsrmkiTaboIBty0R2esGY3u2dbyyYUDBVjCR
AVFFV0Kz6zkouAl+leKmtY35dyCsMW3o0Kjba6KiqFphWbHHmcZQd8AVNkTjwdOGMg+pcH4kV4X/
1ShFAP8axaiUkKx1IKsEtLwhVlG84exwcb+qeF4uPm1vbZXEuHjVVyN5J5OwwQi4WgGHJkro85CP
wGMrr/Ja7w7Pw403QSP1i77R5BuNwV88OaHY+ME8ek2InLrds2B5BgTxG3pNEL+aki0v6rptYO+/
DmMqUnHOcbCWTLEXFdPOQIEW9JuVAAXXplPzutZsYPw86bEDa0pEoICshBC9THoh/Hkgfh/+N6XW
ejhPPPelFpwWY3QNPpOWdQU0UzLDdiGV7ToUU0o+SKpicNI1VhR3DbM/xxASqNYY0eL+BAXEHDle
gV/HHm+Nt6pBGcZR6pzYmu8f6aTXRlI+mBcInOx6Mc5N3kmd3VYrR5DQUxtDWvmoyYLpKiB4Ur6t
2eO6R5cdJ7RYN4/MIU5lV/H8R3YsHgMp7UPrArmJOKS0tPIsROu3Q7D4IngzO5mFncFjuIyBlGGK
XnojTqm0PYev6xhF1zEEhWA6HrKxy3qoPXij5dq4bRUVwmUayoGiZ1csyeMFCFlFzRqLhXrBWgY1
UhTjbS79UltTsjV/nkU7OqHGs3iPMzK1oLgWI7AHwqKZkyif9zi5Ph+5UiPvXxEWnenhoGsTejQk
aXhx9qQfNIPJfewiSPI6ss5NPbGEQz3DNfMyfSOi9HPmmBIEV5x3oMX2R0ay58ZpqKbxTCrsHLYk
LqT0abvNKLy4aSpsorNGkk6DdagdupmgK3gDj8Hj63yBlPDYB486LHUzBZymbiEmQHVYb/Vubu6Y
JPCTLeycISuXJp0r9zRypZm2xdl2rQxy8wI1d8ZYQLNVfogfo68vo4q+Zt+bG9E13/iqXyO+A2WK
vzubA54L3RH3pkUNJb3EHo/1u7wf5JiGc1fnHSz9CA5422xdtVNhVRTiOlzOaQMQHKKSdu1dWjE/
mp2lOTnso9RU4+m0/7PCiGjVAngp6nxVw6cgmcrvoOqUbRC0H4jJeCAeVuTJ8V0UTVJ6FTCzpLmY
CqGHPmjBISfBZNzpT43fFZ4fLVk5vho89LPUPR1cCbxJEkXS6LeGD5Uzsdc5ufLSZgYMj1ri6wFm
yKkfkhv3A1j967aJxzWYhunSM2NwU9xJSyUzr55twyNVcLBMNgt5ZyX2LzkS0OrBBPPlLipDtEu0
Bb+zt268wG+FNc4VjUlH8RzujJ05ZjkFUrR3MHkjE66x7XjHnwR0DCCYhXu3bwCUza+CdIa0CEOd
unZl0JDEzKGcLMiPIgP1bPvSSMSduShKUclgXPefFENzRrX6MDXKDA9s9eC/uCGyKvy8zK6VYvz0
O7LIKJBK7tko2XkuN6NeBYTHHqgL6iU84une2jT5Z9d7ivyKfyFj0GXfXAOrCMOHdviBs2C6fxf4
rKu4qGrevN4S+82izOflK5sM24MtzMgnIi19d13TbJqmvDqVlBd4QTXimmpT6qhIPXDQAmHkjf4c
I2aCQDQ0oGr3jMrCry50UHibZu5kYpFa1ylifkO+d3eCnznM+ylJFhBTTv8CPkxgwLJLd/TP76rg
OYqZJn1cr5pTg8b/ClSGkjl2lYkg+iaog5VqOPuMdcaAMylXuEz2lFjm3upUriM3Q9UYGebAoEYb
hPWYUCQad8fNp5tu+3kJq9VFBC/nshdZ9CdsuT5Sdm4r9mqwzx5GnwZ7AbExf6C2g1zFVCInfByK
pDjE4+qXIO8kKAhvgW5As5ogA2BqSfW/xEt3ogPCoEsYS2akcDIRI5qD3XfdqwJVfUZgAQPqXlBI
nPYZg3dw9wmpxXOismoE/wy0eQtCGiaIIYHtr1dh4vTFuRIE5Mc+Jjh6RHpY46IhuFZbfNcsVcrv
RV3COxCw/r+uNhzOjXIT3DzFW/CZPhF1oyHBSYop+sIxHg81/sCQYvNJvZcTVJxNIFf5B7kjRpfL
EQ0lt8KuvbRzEL7LoHTzJ5w9hWhkV+sDZDCcsaM2oPL9sKy83FR8u/Ptyqo3JA7R8G1W8+jOgCX/
WMxp8q54JXWANd4crT7jE+AB/crChgZmMaI0Jk3wswZD7FiUC0JyCD9E0iQfEVBkSsP2+6GYgeBz
iTTcwVq+jzTr4S3A9jg+c24iptgq00PZQQ/zJjnNmqkxRAPZqVqptLEn/JT22vPz2If93XCr9L1X
/EYT13CraD6GbnNafbt/cqJrSIwH3jZIkokUqVif1S5CsfKSaRpffPwzkN1gWb+y9ysmuTXHue1A
IRznvlSo7QhFUWfKxBkSM240/sTdUD42H1LWdcco579db+pnKsZm6Ch0q+8OcxRAHDUSropZzaw9
RT5tAbBFBXTyNN+PHzODGjm/SLUbhAx7R8RXQEOzDbF5tY4trV9OcbQEOVNISIq9Qd3/SL7FrzFD
98Zr0onxmG5XA5l30fND6ntgs+tGMNxwsf5AKcPFX4vri6TEr+mFdHXwCTGPq0BZrZnrRsFtg+8J
Dzx2EsEK9/3LgvS+VH/INDQ1WGT9BkKAHgFxKnrI6+tx8bfDaDAzc2pqomxNqKU1gDtOBjOCEaKK
NzR4Wd6+o07+fUnt3PqEnVoHFaU7+heZBQFYZf/iBtEAMESrx+P2CrakYokQHpbkDmZfvHPvfHb4
u6Sni5vlnn54Ey9IJT2+qtx0lbOw9rGYsbcO9iTg/WcLEGNUlJeMeSMPrYu7WeZbWJiXsY7JYcU3
A/nO6m7gRvO0jTLcpQcKoMBgNNTlmteEuuo8V+FWHXv0+mNkU7HkJYAWLWIpr8F8cJS/2h09YD4h
kxjo060m5xdtR6jZy/V5AEnj24bsE+QX1wbsgEHHtXNGtbgpVgQ9i8z7ZoUNAdbxG/DyzWjV4I+J
1fA3I0N78XRlCRJ1z1nhleX1tsttgahDOhegkqCXA+6DISu0+QHXFMDXEzVM1XB4BwZsIRasYQje
ma1TQEehE71HS08BYPZadJyYZSqP6YrGBVNR0wbHXGEulGN+rclZA8DL79dGVJzk8/4uhxUuNuJB
06rRNqdbCjbv1ya+DhrS/Bdo9sXNXeazhd4nQ9+FsC3C++BF0yaxavaNwSdbOXkrBx81nBHvuZpu
IiqP3t24AwEtowhHVdQa2WIYojOgv7KuTet0YfFe5Bn3k1wPXKvOggAQuTRESVjUbiOBW0g+X8KH
doFtpj3lktKAYQH2uD7PMgfqZ8aqBezuyxGcj6WQHEIQKMMPoW2A+zmQKCOjoFlTOo5w2IqrfWmN
lvUEK5rrMA1EcQyK9l/8O0jzgrUYXGfHYd6vJUCscD1o/XPHaalTuCJpXzpLm0+OKTf0mHof+jRe
+tkw5lT4Czec3R47b8gr5v76CnZIKSA8mU95mqll10i09yNFRjPkwuLMuKQP7v+tSdGVJGa9skLV
RjtaAa3Ajq1QkODPJ0Lk3SJRDyF8FrHJ+ON10rgplakckueIAln+foBoMPCME50jPIcZWLTyj5Q2
EEeM3yB746fYXjGOec1Z+gIoF7CzZsWbIzkXp+WbP/Aw3uX02FlYAAkVFVM7DNr1jnWVjdftRrAN
3sYwoAiRh5OwKRrxry40LPYQlDYLals6QUSva8otzXhLqPVBh4hu0Lo7bX1puTKxqo6h8FiNJu6Z
iCEO5s9T8nY5wZOoLAB4Lg70E2k/MPHdNiCWKkmGmo9paKAt4APf7n2rKTjLIVr6Pasuwq69EXsY
DSIDgWb+x3oAeDjiOv6mmnznEkpX7moXd/hL48Ocusy1kue6C/1nsSWzcJ942O1pYrdyFuzNeqgn
HVH/zki0/V3tj6FsYSpCgVN6il6pJgOm1Hacc6x/s18MqEMP6abo5pO2phfHi44pQGPFGVv1bNOq
yj3fY9HLKgcQvC9n6MlENb6fbNRz9+90QwG2KYhCukUsarxa2m/m0k+cRD8flfBU0DM2uAkMqHEy
hkttDNFwXASmXebKVRjLGffTp6eKK7mPSgSD/Or2LvZqDvLxIrB15jXQw1DRXkz1YLzwbjy08EvZ
AwTipMX2vMznuReX2bmPrMI2shm+9TMl8ndaMHWOic056unQgvO7IQ4MAK/qRh/0z6+6Fce2cbv/
ZmCkPXFIJJVhNjem8Y76xMEpEg3tbvTNiyAxmL9m0dcxCpX0KaKEnQJAZJIwmZPLNwTTu//c1KMn
vp8S94Tz3Wr8atm/C2wSB94c5T1RhZk/VYXDL9E9r11V68j9OBApIxruOblLum57NvttUI3dXbSv
mM7KyLxq+6AUkOtxxWdWbk2lSlkeEwGoyNJ1sNALalBhbmPn9XmJdIL6DMVriOsinGY6mlVbi4i1
ITY1hg8da1DmHIAZVUM/q1DRLDMZ6kR5UZ/ajJCzD9lA+Yry4FqQ5BRSdw/nJMWjcNW4PbqHgd/5
1Ka6mSc9JieZI36Qgh4TCX1OSUvnF69CiJVWa2NF1iMSMkjV9u/eYjGdQlP/jk7gf+m+VaXYA+Mt
Uf7LEZG5V2QqFUtiBrjmXW0AQ95SxKV7kNiz6FM0wNU3ZC7RgN6Z8CcNRzMBPBY6yG0zweW4g8Nx
IdBm0516hTMHZHSWuU/hkJstqdGtQ7+MDOWsGHeqh4PWM+MoG/Q2rbaLfYPHKSWFZPFcDki5YTrN
yfbtzt0BXiOLuxcTYyZk9hOfsnl5gPFElPmI2cWJwvu7DzpUq5M1N4cPccYmPWhBMXu7BQF1P5kv
WWd1kgZTlWQoJL1pTwWbVw4qKGmqBpMxU7b6ghC3dQ8tMya9AEpqNeIPq7guU9WxmWx4WP4bioGa
UwmAWWnmMnFI1jGLRMx4+gyrsDiD4Hmo3Dk1XyjGWCDEqUwC12W5ScnTv7P4xSxJFKHS35iow2+6
Ql+cne5O03iRk76Qxx+pJtUkOqgODqZDOzUvPNy7QCUXEq3gVXO1YE88vo3JmvXLP5FSlgwiI8hf
jXA/g9A6hjfMobhOC641ihx+U+HnkBFD/mw3pwzfoLYGZtQhy+k3okYtaWbWlgSMQnH8w6OgXYo/
xD37Eam1al50KDyck8/MhFfoqF+g7pYKlSaKl7+ZR2gzh89WuSkJ6dYtrr4ZNR0d5Kwyj4HMNuFE
qmsOe78rcT2Tj7s9BnLSsFOJHUd4tr6kzHM0OtxjXx5rDykpitnwTW6+MYdl6+JIHstMyoNIevEo
jUxHqrjHEAJhA+41TdobiDRdjtz7Sgod8jQR/y+6ZAsolywyD8uPaKf9kz4+rvish76R0AoTVukH
BkTG5U6eA3zCoZsZiv7sD8HIUgX4/+nZB12n7S7GVgqbvS9cJh6ExVvonFgdDxQD41XEqskKzhJH
m7FVVHWi/Gsmm/eFzXOG36JkIbkSe/vZy/apbbRMuHyB/DmdlKp6MJCaFD2B4MJVHbUeGezcTtxy
OZj0/OINRVZIQ7HV7Bq8KhLROocduHm6dO81jTYO8M8Mb1dwlSUut0/g9IC6bc+mrXcDZ9GYSl+n
Wc4jyPH60QImuFQyZqRD1MnxCmYQ33hvxgiy/AQKdXoo58dybDWfs8rSWSrZhwqTwNNHm0xrGJf+
mr2evZ7JuFx9N6CVyzy5AvVWig94djmbIg/jMqgKn646gKs6iE5ZvaPQfp+6HyLnoffBkZL5tAF7
cB6KNckSHGTjcWxBXP9LVWdNJkAJLkWKzzwSfiQJMfO/htS/5DfnnRvWvHmIR50UxghPpfbEW/+e
db4WOBAfL+haIDiVM/q4GrGnwKOSBuxw1icMZcwn7Ilr8HawJlRXu+zJvow6oGiQMaRnp19tF72t
FMLoOEa4mjOf8Wya4TK/35X1Q3tiOTgRuH0r9JXvQ7gAdnA4WecCmknvTv+mDCNzp39kqhbweMce
qEZdTqGrQc1e8NIiOlXkIJdRiQRq9wLafAj3KoNRTMWAkDuvSfVfBMWnqZqpgd3vU0gqnVrCJ8W+
RYs98EmwHmV9xGIMQ0zSBhSqutvlaR+nQTDqwfyRQEdzDmtDwWmBR+dUp46pSSkg1JLgPQR2E6cX
tyYuvi7v3hGcYwtBmP2uPq0f1ruPcfDQLRM413geBa3UxMm+1wPLzMlSNg/kqtCqCrT0jH1bZ8WE
C2QasR7S7d8asqY5Nx4Lyt/fhuhM+NeUvulALlTmRhsPsJKvQzckyxRbqB9nCIIHsvK150IooB9H
zWZXRiB9sPF0g5PZUq0ISUzrQcMu+c8q1FlYTS2LybRDJTPYGXg6ZIvalDO25OR4BjSOuh/ZpbRh
FNt5HxLZ8k70AvqqKpXyf3A8ALu1F3ydLXFDVpfD/awVyPVRRWUDwKrZkdKoBkVO36vUhgJbUgsZ
egB38+TuIIVT8as6lqEY4cr7Av+Et7rgHUmJV+wfiqePjbLrXW2yyElTalk90XijLiWCaalAVgXA
eyxTJvcUEE3KnveJYkYzDnL07HcppW/8k/UFZGdPIAplfPQMxlm0xYVdFUadzzBzFl3xgGsCr1Kn
o8CV5xlAI6b3cu3pAUml10WpbdN8xXkARTDLLXYRDQcABgD4oBbuOJMsocvXzjDSUAJrQDFORokC
X9NMHs6k3gWemlZ7656j2DWpHAyx2xSMdta0ViVmCnIoHpuTv7gphlY0eBjGr64NuDYPv9RasKqO
UsTz/ddRJMWEuxbfg+J65qNHRECFDWWYUglOgxMfVHK7OenJdC9/ZfUYopqOyvgu6sw8/M/MV4sO
PQ7gS9HvTcAPZz16lrce0tACwdlAIa+iUQGRi0uC3J3sTmi1ahhfUtGHYPZJBKn0f2FV1Xg+tTPK
vTKZvcsNUooevuFCKedu6fOGAxeBtS7oQhg9pby6OCBV4YvlkFBtmG/3TqEMoK/UxpOvYVGFDCOW
va7QOYgNQB12lCYkouz0oCRI3VhWhOjjSc6mf/VMsBqxkxTXNZHEi+8x2MadZOM8f8pDKRVflSMH
3bnyt/gChkyP+E8854QsvACg7XqOg1ocQoz3Hxc+N1okS7gYpT+PF4/Xcq/P7y4OdEjZ2txtR4SY
TlgB1/6aZrCcI6vJadoKWyjHakgcY/y3sA6rNK8aXwNS2KhPp6fFQEXLuwO2epXxMOQIet+rBABc
a2G2EqnVvUuUntFMS4m50o6B0VKl/Y6wr7Z9Da0FbpXoAuZ+mBX1ZhgvmsVqB6Tub6M2AXUdjYqq
qM6yvgzWVhjGvccy/A7POPBK/Sa7DPozhno5d5Fo53EHC4b99kFqa2L5neQa2fbwHUdgZ2FOU0j6
JYlafzs6BTPf+zW+d8b0o2nl3tsVPqvDGoojGn5WoHlwDveDRD01CskvQtYOgLEXXJU3WS3otkaV
dbwizuzPqTVcSmqTGa+la7qa15EUGPIFxJeM3XZMf+LzDH4vwgWE2h9r1K4EThu+QoUeGxRBXFF+
8M0Pq9yPXpbY+1O7tC9Hkw9fU5rrwz7IHbMwwl7ZlNcSg/44KyQ7QanT5HADS/aOdCcADzeWhtas
ZWmfcpPceI93l7O08ti518Ly27hyucjESyBexxZ2Ma0mZ6GJrvgU6fvQ25ijqz8pSy9A6ozl4R26
jJ+r8kSMhyXkmrOqT9nWPSrdMBuX/BIaFma2NB+UcuB8WQrQrEaqd0ZZfbzSQji5RVO7aMEfwqPl
mol30zxT9HKi4Xbolx1zIBo7nFm7z4ORNvOB58+uMDhQW+L0BujsMNoryE7sC6uG5IeRGo7MQGfB
ooOXqutJUFLC22qWPEqPOnIyelTqRjp4Gpi69SRdyvGSlw8IE6ui0Wg1zNkKIteRCCJVb7SnnUOI
+Xla7mgYiLHA1Mp9w4+bQi/8JTtq+PLaeAn6bTEciSzkDs3VktPWI27Rp4Pd7QqQ716Mdfdlnm14
2GPz4XoTIQ/ba+pHNtcgWU0QfI30DmX3IUeEHx7EQbr5jB5SjHV+tHs/ZxpfM8pjfu8yRWYYEDvx
VqwAlDxSbgOHD7q2fWDNhMRsdui8Ar5BN10mm4FMeCHOaFjVgXckDcv57Q6B/55xfaTr++sHl96Z
0dBDm/FlrdOLyXF8kKcZvBBk0Y+/9oSAXYQuxqBWG/ZaAjY+Lxx+oVBOGhd+fOxYtOMAGZNzu0c+
QbkZHo85VX6Qdm/nLJPxtTJnW3DePlr5vpzfCZY1ujagkpFX+vC0E2x2OCFkxa2jH4IXb6qwQeO4
s/gSV5xe9v0pR93Kle1Q/AsM5VAIWYYZGV7mmlhfq76gAq8RBD7g3Nqa60yZ+JrHErtuwpNz/tkJ
Y14sHmu83uEDdrWQJ3HQDq+ufIj5zAijx0B4OH8al9EvCbG1OroMReyyhHqrdMUL3PGw7q0rjj4n
A3BIugNY2iNDND8/WWwZWv0gPRkDbcMZ43hgMTLIqS42fY9imXM0vKR1oVYZIKoyCnEgvL3cQc0Q
/QYDAPT6qLURmUY2d5MoDtqPi2DEm7F1jkzh0xLciQOFmFUci7u0PEFoqgEoG7Ru/xSRSSEwejur
HOsoZjJn9Gf5SG8QdCKFpirib3Z8jOikx/KzBAcPFHHiWWbRJ8hcomK7DPo2fX/ubjUqvgokCAZk
c1Z2yPnQ5K/NF31mmqQ6Z7rYSIsNpqGvFmHg47jI0ZoFL2RCoz6Mdji4QCYLnAcYUGLRPFV1vTzV
vh9SYtEABv/Iv6icV1w4hGbkTM7Kmk8336fXy6CvAgLClUhRCMRuK0RMQSs4c9KhkQYPbf1VLg1D
Na/5PCjfQSd7aN2jKKcGy09zgvgVDF51VRVtGDyp8xibTek/TKKK71jjNxcgw2zGBxGCuFWJ96bF
7dEehwBSys4AkGPIWNmZuLWFCYQ/HwQWynIaq+wRSJlR6LcTc93XfXK0or8hXalQBoFikrv4ls7W
mZICPPx2JEevY16tIwy+jQaCdxGNUlU1Qt4uXNaV8TSu5vGKI8q2mGfcMAig/dvNTL/vp89c0uMu
ij+pbEPCRIIRRKZNbYkv4Y3tUSBkg6EsfHr3F6fQCeTCFhHN91SGPdFPIkwjnufVcl1r2CqoabxR
lKZE3JOgFAKjPg3N1jzPpQvlaS0B8cJLyW66dwUkGBq6nQEVrU6O5fLrb7/Xr+/acNegkGscq3je
/3dAqKwduUFsT/gAYF1RTiLW2YllPGw8TIsrTEZLrG4hI/cIEZ1GRk+VwOUtbbTVz9xca+KKiftI
u2JOdfnqN80sFxU/GOnG59VLTi0yJMG1wi14TQTdHIOyGQnLO2k2I7lG1Ph9Go2AT62R6pKhmMrv
Y6VRhT2yjmQFeMsE4KK400HyyVLNT8mtocPhVP36XMk0Clfxyl4AZAZGS3Qyt1bD5P3PZO1XwJ/3
SqkqiCiEaDcVqE76U0yZDpkga+DahkoVuFDxv20Oq1IK4wcZGT4H9wJsMItocz6OvlEA/NijqMXN
uURcpRxCe185dZ3HLsqYPEjj69aOIG4S0JsFg4VzAMguk0B+Kg/2ZMuUZgfulD+p/e36KBEAVf7J
X2sUY8Ex55er5TDuEOsdLKvq8BSw8Pm8/iu5f8cyF9EX+UAsn8j5O0TSOqeAd64SLfzBUiEwN+/N
gM1As71q82qAjO//8MlQHoIr6q/M2/mVPmIOmTAX0n36g4SaPF9w4RcQ0W0UFvpShIsJTo6QbErp
90m6gPkAFYrqPg0WOg1DOiefRnA1EpByyTh91ACvF0lOPYVxW/QD3yYiX9D4z6oOe9u/9eD1aSod
nKN1cTVM7WWNtobfPcZ02mXav5gl/OV+zoZiPgcQXYIoNgQBrUu7KCoZgg/xoEznuRfBMZakDMq2
HF6WsgILF8CVEN8u9sRuE+5RjmedJ8Z9C80mvIeT0fjtBpK3sGhNUH4h3lw6HwrtZQRzWAYFWCv4
hJjhDXO+k/eAKGTTXURiU5xpGtSoXEWE9lXzVtLZqwbqqECc7IeWlqSjJAaVTVcDSdaNxw5g6YBU
1UyT1xpYHNh6MLvKCO6XDbrdeeYwvWkjU48OmP0VLcD8cDqid7qPKnVdzoPra87oChqT8wpvHCc4
3BjFcZu8ht0UyuFkuVBpZoF9W5CqfuxSJv2N3vYeEZxhAOhFKe96gKrygKH6+7gdU21k7Ju3JMe5
ZeqOIqf6JcnH1Yt57iIQSgqb/r3Y+fawxd8SyX94sXsrxBT2dFmBO7AyUl/LvZMXg6LwdmwjpeEJ
ggP54A5rNNG5wqa1EqOCM54gYAQwwXpN1O+XO+DWFzm5KU8whjh9SFcTG3x1IjO3if+rZh68BZb9
kY4KeBd8mwYUutEyag3mJHIcpoxUKt0x8gg1WpeUyLQvoP0rcmr0BXbWdFP+uNesmNuxV1g72IWo
fJlLSghM78ujMQB9tH7WfoW4PWc+DmMP9RNrSkcbSmTB3imRW3iVPuhOHDQltbN3NBmlOPoziAas
yoVkdWpHU1kH+527Yt0nw8k1LXsmrUTL0yz6u/jYLTeHb0U9anF7f93zjehuUKCsWdVT+NPhGzfD
xdqLXcj1IzNfAZjvaZKfgs0pSLpI2CgYFBOC5bSZiIxgLkX99fEczHLchk44WPQbTcgQZFLM6RX/
rkE+kyqWVNq9J7ucftT0Cpxklen692MW4Ul1U1kuu8b38CdhrESEU/nVNFWTdPenYTytcuW02ek4
hDERvt1SQpVkLMNVv+knsF04T6KBBkZcVGa8URAGcEfC0O3RnENVUSDsl5dDqamyVVwNH2Jx6mGw
9SGYrHdnQTdFBOnKPG28yGNBmM9RPbezhpfGvPljYxRd5y/4vZYPMRbmFEA6SMAoERX7alU3lC81
8qImMUMZ4lmAenQMemg+WfPx1ycBmOtdKp1SA8FfypcrmYnATIdl1hll7PnC9P/0SMn4AgGWJ2DP
0RCIAmT6yTt+yna36Do7bBOxEB3G83hs6y9LWfaeY0JWbhcDiDRSAUkKlBGHE0NUsKNdyLojEReq
Ehr5h4SCyz6SYTj3VNGbeHEZJYjhnCQI3UQAviNPiG+K2bonBQo79Qhl8X0nvHvgdmYUBjM+7ZZJ
diQQ7FETRBbs3o2Y/sMhJHsgzMKwsJ0B7qS0xDxgHuXQWKeOvodeJiWrz4V8Yxd3joVZ7k32iOaL
TaiRRohV2D5iC+oLVs4XTec3bLEBlw0/KjrHLiq2eusT916NzyjlgEIM4zxQlvb6UdtA30knqeCu
8fv2z1ZOrlCylSZ7s0lBRpbeQ7Amqnfp7PaKw1gwWQ5s7u4QvGNagjuwtG2f86YdLziluGfmlp5z
/a9gE0H8pC3+wwgAinrLymmPr8mStAvQ2h+JB7hqIuwudKm+aGlmQsYVpdHY0/1Rv70Oc/Iyu3+l
Bm7MorbzVKsS+KMhF0ZXdA5oCJLpVVaBYUKbmNUYfiavWxMrZ1W1wZE1YuKEZS48E6yFIfEHTSjv
vvDd0AuvefcwaIM+yzdeXc6mZkoIbcw+papS3zHt8aEBjy3mogF+87LPrGLYvWbhyUiz+48tHoA8
jl9iQuykxIjd9NDCKesRljeyDv0vUTGHhVkFbXfhll4PivcKPOFSpIcxnlKFB1a/3KYDj37vIUqK
ykt53ualN2JLLCnPWerzYKtXCtqm2R7oUlJ1BaRz4t88fch/OXKfCYsqTGkM9IU2/KQoYbewTq/6
0dz45pjOSRMlf85yBusZ14MologWD5G+aLRRRnBJDJcOgcnC5CnASnB2FNbmVBzrG0zEsqBEWciB
eGRl+QZ5QCSUt4d4BlidimSReJs170x2Ml7OQAo3FNR5aQFRaWnuGdhxHhbaAFKijxdA8p4NqYus
aQrH3ml17B4yeb03asoBTJ8KFXOBmrFSoGVnlg2Y1w9zAoku6DHHw9W5ta7Mk/SPfVaLIup3O8kt
xrs0m9LaqOI0KX4yC5f3m39gxDiyiklxWzS0U75DfwwI7QdAoPZ5PVB373j0Ag4Mma9aI3vPssdc
VmOuZV6YFwbVq8thRQTOmFcwnRd5/fyI4rstz3UGIpUkuisZpSZJpXVn8ZzuxWzppvykBHuD/TD8
qw9y/xOl3UTwe2hzWX38sG2pCxPzTA1+KxsgjPV6kDTpNOtv3mz9Ah7lwEGphqnXaVtMsKm70ppp
ZguQ4gbxixMf9CMeo+SfnQj5wM6fO27eBmbNV7VSZgnfoTPCeTqdTRascTc31raRfSycbRIVvJNj
l5NNpRW9+NBcAwitGccFQMadPounngAwuoFJOiOYQo/O6olt1fJdrBFoTVeKys7JAoklRPlcUZIU
PBdJ6G4WY89EEh3mTUga47PgkXrZ2UnqzpZqcEEhyivLefoVAZt3JVyhCq1it5ShQynSgh5J37r0
CPdZy6HbL4YEpLWfvXhEhJ9hiFP9GqJ6s4jpcIDv6zUJH57DqBO6WjB3hEJyC4w02NU/iljz6+Az
X/3qGsoUqE6oO6TzTt0AA21D59GmIqW2cxENNq6lYqjeoUqaSNw5kKXl5RqLEOPiCg2SnI7Yji/a
WNMXBnxCmIDslveGBXAsYmuppDkKawh3/kZWEgEtc5zLtvZ9rMQPBTgDftRPsp3wZnEja3TCmciY
X5IcHvSOIjD8noxsnUpZeRG1sUuHUIlzkRs4REMjEtvYjHJB32pVi6kQOW254vdt9w3lp8YijuwG
3WyT9oCHMj634ETdcoeYD8nt88fjkhRZkAe1l3/hidwtxiCVtqN0xc81DDlVrP6tIN6ziKGIjRlI
MrA0StgB1r3kMyePYBH9VeYgOl1orFL5+ODRhhMQl8cOFiuQoObMOMSGLImf0yHZ9GFlnl0D2ck+
9ZlK4PLVKnojadyVpKZz7Q0A+AGeV8K/aMV9h8mIZjn5ozd/dsEFjrIrsZpWCn6dlmRMO8c2HADC
J53Cjj44k559iPQKfGKX5xT7MMrfXrbRq2OKlZUoC0LjN/oRxpG5M80ydmSu9b9ug50fw/qODqTC
qiXrxHZTooJIf8UtYtnhq159ad1gwJTSh47EPG8wdtlODrdYM3ADNjid+L7ZoPzUH4iqZ/nCcFcS
oms1r2I7sDm8s7cRuAoPIX8ofWLA7TEWpBXf6wd7hilRTKcfEfpOKmS9TdsxVE5WsM3FdZ18rFDA
i3WNoPzSbNTKJYro92EgfoqX9IqdyrUFV3FgaXMZP+ZjQDsU3lD2DgOXZVzQUllJrTEfBuPyhblm
fJTHba5O8aXgtJzdrfGQhoySeIm7xsagkONmlfsCZ5mAqS7+Z34dENtAE67ztLKT1dPfiUxldqrE
wQbll19a+nfm0XVdeRzdBs4eXswHycSLsi0lirCblhl9pA9jtbtlxj2igreeLSV6pOxxjwZg3BhF
SMxizORYrXr22GHqA6U+17WzsjVmkECKKw4xqO53/zhIRjoO/awosjUfyphgLnsZl0geckghRQYC
aWdfK2GI0A9D8KDMcdpvyjLKCHaCkursOqkyCvCfuVDEU6U0ISjkmKyZFTwAnMe+qm5/ah3Gjt1F
Zupu9QZ8XT90Svyb3z+6fHpjF/0LpT/rv3JArK/1Hsf33So2w4UqjINanCquZYJpi3zhlzEVaRT3
PowtYomlA9bu4k5HaBPathimuUGp3CghOWBhgnq+w+AdgKLjNsrD4YiIxLD0jLw2XmmgZKJ7vsmF
ubfJOJirGpqGzCx6irLvTSSHkDLBe4/BXmeRKYSib/aIMVeyIzzJe/bWqIi2wifII7/xZQZIV0SK
GiFnwBmUhWwLCeTzYts6B/jqvGcbfOmKgwnvTpWZZ0vWD89E/k71oM7ztFn0oMlavpLhjBDwbVUv
MkYDaw6h7tPxzE1R9WGBkA8H88l48OwGvGF/vYQ4hzw9cMxkoftkgR2R42ifpBpNzH6RGFzWWc8S
2mVuQSJ0F9d6Fwr4dsYbcdf/Q135mpHy80HS3neNfdf60LfNM/6BQkv4SEwPXNu0KunmAND093yU
Yt7NL9EPmacfmULMMu5AoSNcVgveOiSyKXVU4lWGXiY2/CQgpZyHPOlY6fc9GGQ6/3Obkhshli8i
7mUv+fpZRMQuVwJ2XkjiVfvPhHjbTYqLyWsKYg+DAgunYrzSyJCy1b/x9wf5CQQEdHJxWJFph8pa
7onje904EI8xQ0Hc0cR0fvpgDqPRHXZSuu/pyaU/nbRwGu1ll+e3JpinquVKTQJvbJN1C0rl5TIa
RCDi1n7gCU2k3cqNKZUuQAVvdhd9VwfyQ/4CDzj/pdWmvHiwhI80queCpgZHPrWq25kWfKTC09aY
/M0JcPpJVD2UaxwRHCbeCmqfyXb49OPkx9pKtdsEKOaV931bDIHwUZZxVCddmXjJJc/y6OWy8c4+
Uc+5T3YVqpUQ370PuXKGLPapSUR0z1fMES+0w9XiOziVmQUixsCBBuXnV0yav9qr9z2b8f/cWKvB
yXcaD0GOYm9q7X/D9xp3aiE8jgnyK8NkPtppqeWeF8MCjmzH99aRA67khZxwqh2zK+J/W0+GRel6
YyuTobrWtLW9mysO6Rewm3RI3jd9h/g1cGZC7q11nBDSK5zD1zTrYiaBGSKd8TN9SDMj1wf8zlNj
mIehBAZE4cFgTtaqyZFxXa/OsvyWse42hOTt5VG2X/kn4Gvn5mbkihAYd2OcN9befpmdG6jUpbvm
66/H3ApCNghB31jBRMZ9Ui27HGTo5j9MOL8Q61894xmpw5e8nCOQZEx945bV4sA2/W4oyktwyc29
3kXYkRtSx0k4wP7qoQ66frs69AC+hDHs03+d0NMeu5oPTfm9vEu/E9HNPBZRoYvxYPvbwxNl73M6
5QghjbRGlX4w0PWZVa9+8gSY2qKDIVR/H7R8F22TMul1jJpa4T/4aQ1gzHhrbsnAZtjJDx9JEk37
A1w37fNzPQkA58/q5Dw/jE+81biuEGwSSu21e+C0Ok5BZjsvcjcN/r5M98ZtYtSyo5+JBDUf5UDr
2rJL+H9OCY1FbaEr3YXnOgoUscrJmIPC5eCdbG4Ml49OjJ34t0pR1BSUHF/7sV5SPuYxe9llu5bP
EzM3aJT6eGWNsYMKJiy/VMW29qkErUDKgrCoxi6f9XxCqilbo1qucjvtUyDhfN8vujQuFKQPKjSK
tZZgOP5gTRO+Y8vFNO4+XFSoW6odFqnfSuukJBJrwUWUH4tNstR18YlpGjg9zzOf3qxBU8jgsg9v
HWhbBdfXfirsc3DrbNt36++fh2rFg/fURY+UeTpDZ1bo0wX85fg/w/2ILwjhgmBju/L4rpjz9WiW
uv6V3tINl2s6fnUyjLuyCFUwYahrPeP5vJR4ZGgV8lsLo6mEOq+7TucqTcB/iQbq6iFg04KaB9Sw
lDjgSW1COcUPWXLJ4M89SbL9KFUy74mF3POft1N/Dz1NK54oolqpempgpKnR/mvdTGQ/UheVGuEu
7wfeeY8E67qWIzXyshOEiN3nVGM624Ys9moyOxf1wNLzw1QK1ENy197QTZw++cKA//Azbd6QDK0I
SUL6eoyyMtIZL9SFxmRICtYbI9e2VAOsBz25dfhB+Lw93i9D2BpwaDosoJQV/pnLmy6gesm1FUk2
73ZAcm+FqDziYbeOjuD+lGc10VjnAlAXfYLHiXGFebD8IkoIBMY+dIqATwgyCZV/kYWckDBxVqzR
PNsSuvPc6Um7Z+PruKMUFnDXiBQzkwTaUmyV1acmzzQvbt89SHj/1YEqMMPorh8KIfLjee7q3Ypc
ROavnbMO34u3aJ4NUDKggYYHswXhxpnHyF0y03TmIbg5rQ1FDH3Uzt9OfrvNa76+cE7DrneDPl5a
S7BzQDzHyYlvpHZ34C1vvCXmz2kMXnpxkut6FKU5bxvS2Ek8OsN+wY5mGu8H5JSBD7FzK3oFoGlk
aGDaSAFrEymqLXANvNBMDxdayMDmuT0RUytOtVYR8XuL5EA7PQuT5yCu7OIGYezkx11lEJMX++O1
2dkQOsLO6cxM4h3NW8VRz8VzSnjJ6O33vWvzUGE0JmYhCBp48IldBHiNofbIj1l3Wj91RqDyjzh0
jHKZR0/FT75/XExIKgWhPeQLHL0L+pHeenLh3MZCgbEs5HT1kNvPUA5Sj9wkWbsRdtj0CkzyLIXL
O1zDoTWST0z5SESqclFCvz27nJBvMPlMYOsA4q++054OmU8O5kyCfC9Cm1XXg1CU7Kb7Del6bxl0
EP1wC5GIf6WC/1F9GWqDbYoMDagUZNYQYrZs3uOaMdhoZvLxdV6s9qUNZbmb9zhe3C9UVyY2pnuL
CL4Ym3haJKt/E3z9fkRIKGERCkfjnvCM+3FOXUiFrSvyLPIqrC+PA8/eNMwHTqbnl+XvSevARPm1
TXe992DQ/VbdseLNTM3D522GsdmqWXY1qqgKF9XWNnuxWxXRZkf8i93T1xJmdhGqfu0KZDqp8zsr
+LBXlonF+vo8kmqTY7GQq91wq0WI2Io6bcV77tFGSoaq0wgZ7RqZcqKXH5qa0eIs8bmRQqdeNqUC
3CO/xxnjbu3J0b/DgFvwyIQbghzA2uJzpP09J2HVlf1N2U+SxJP6bo9E7ZLdrcHvMc6VdDMnU41m
xre/+ZBTS7q5dsCv88q1oswhh5sAFd6T2eAP+a0epzTRSj4cgUUz6jfb3aJfmQzEu8sUVp0+CnFW
Qm2xsjAFcZRJtcRhEZjE2z+I6jeyx5tVGsrpAgTFjcwY/L6Cc9xhhjfTI3PvLWIdFldI71NM9p0C
oVfLW89tmCTRG4dbkEc85XoILYMIneNCykd4+NbK4L51kgxAMorRayrf68jAKBhkQJcRjVxvazSx
QPrwT5YDt9+I9hF5VUQHlYjGiq30edpgxbu+gqb4Rd/2kebkcnqRZ0/z/YsnNo+/YygQud+pGhu0
NZAovM8bNSfXjzcIU3WOJKMn0Vc/t/h+EDOz7h6rEAvBpJAkU1+UvH7rMvos+HnuBkrOImA3pXVa
GIpjshwOaxl6yKrIHl8TvKJonBG2pUMXYQPNyVG3e9REH+En4LqeXebVnjRfFu6KzgH2a1mrgDi/
DiA5t8/Syo/eM7MtbUkleFpePRG1r0482EUCWZ/dwkg62x2IkdHJ8Ty56bLWCSMyEtKi5M1Re+o6
IyZAoaBHI24L+guYMGQAozCCnNFlqZ1aQaDWW0FrQxPdEvN3USnuPcqIZ1E0aFMBHAWx/j4a3qji
8uGyvAiEHK7Lytu4YYab/+FDmuPiozMVl/hIKjo25AtHKIPyu6bfViNEK/IiNY1LCNyBRBgWnQHy
9KeH9jWyupHyeHTye6zOVQYqKY8aGXXCRKsWBwtLIAfOQ4lgaBRYONWXCPbr5RwdIgR8AH41hS4c
pri5Ie7bmuRg2DapA10/Xdxdrevm3oSNcrXs5/P7RRAjz6VpRJgbcr9FK5gc5Zl7I1Z8iUDtaHKP
T+it+4QHwFMKMY0FsrHAEMe2N6jiNIqjAVdv3Egz2hzptABN5eZdPURsVPZcsagZ0g0K/WKEHJSE
6hq6w28OZVYEyk9utKnl5h/bngczb142JNKMeMYlG/hTxUisNRT8b+i+RBSqRQV/lt50sBgtOIa3
hlxQdGY9qx9wIp2zvD+DmFNi/QMBT0FUIsnajO2ixEdgXIr32DnaevttpDocsuZ15cmYKdbLi0Uq
WRzAfJuUKTLKpt8zZWlou1iTLhIu+ydZGUIW7St6g7fk90BDtJ6T3RTEuhxixN/D3YbmFfZegUum
zYEoF9Ra7kZB0sLQUNhoq8khuvFnJVOjJEaC+DBPmIq/BwVb8UTJjEKz3noW8S7/qZcmGMITEy0q
uBuIiOuHA++K+q2LkzYf8uvnflBoa9IQfBv30AtjqkCh+RL01ZXt9atFXs280Aqn3jfDZtFQFm3s
wXiviWubWZjnFU+t8ck9dYhsdrk+qJ0HYAgslepQfHEL0Sla47I/X6BKO3FRiKeIWY7q+XjvrKR0
FMFl2q0s9wEpIZQ74mR4Me23mk8NPh+vTVmnl8l9lmTxDP9NSeeu8gEwgPFRjVmqDDMb7UmPCEx+
bvbiBA0sPFpWmH1gCZZo1F4cgkF/r0NF76jLVd52Mvjx8rT66KNKR8yspTya8x2NtmJAPknKhYpY
AxD5MrYK08LgKGyyl7919iOPFXDJtprDyMbFA014sdO3sq3JhwoBPBn1MyU4BNoBaVnSmDeTJxGk
XPu8LKWHOD6wAjvaRAvCfa/vlxdROs96ZAL8m86AHfQQZk8TdJFJ6WJoPf4uUqqWEzHlWoQjxtb1
kjRDVqcG/+Q2X2PoczuXpn/M1oLxzf3A8SySojASqhmpfx9XnuwMpXNa7eddJOTF7f94g7/rza0E
yQepmcMAyqAFE0M1NXAuGWSx7MNHC8mc8BEYlmyVv2K8m7QhZLmC9gBYdkbjNGLBAxtdRghhjOKD
6OetaaMYyTjEDVEjy+lGndoFZTk2hQuuC9vhjszbGSNFaCoVl0dIqfP/i1maUp/VMNx6aeSuoaFo
W08dwUiOeyQgoq96zbzYTxxQwdKAV1RbJ+QHsxJmJ3vnO3tZvQvdnqQASJhF4dCkDb001Yeiw0TW
Qgb5bqbQpICgZNtzKQCWHeyzNOTSla20uEFHYtee5h77udwHDx5blODP+8ExHCFOhUwy4/6wCxv2
8mTq5MRkG9CyMVRNWrSpaJfU6hJNmnltvwjRtpRXAv9VaGs7b+R2e5Ld8T7nQ8gtprqA+4XdE/GB
xMhvQ/TDN/Ny3f/d2jMJh11UjaF543MGholGHqjgG3BTE7sT1zrQ/x5xnFndBDim9FfUKoHSYROT
93SwGvsxC+ZMF6o8fyBZrcP9l9HKFjoOAk3dUqAi74mcp/HQoPmxI4NmpWwnly//o5clQgw0ltF+
dqEPbRC6DgHOSoVd7COhCRolyT6WASGpahjsjB+rbFmnHSxwCZh/dU6k1L5GMPKJdo2LVBglLTvT
OSViyWouLSeZnEhqf/Icu8a3FOw5DUxgs1RO6as1gZ+c3FYp9edsnlqmegrYJn5c2mZc9J/N3q8i
FfkTA5cY+BPKqD1ncybYRCoN1YrC4HqLVeY5SBkHuIQ3TsV0Z6m+HTyTak2+fPSR48U+mN6G6gAk
SODgzEPbEVzf2W9giWhZ/ZQTg9n+FuN2hG8fk0kEhxn65vmnT5/IbVoMP3Lcnj5GDSjN6HN4yRgx
G6MIzcWRJ350BhdGv59Ywd/G9EzO0kfP1Gq1FrmtLvLuT1YnyuRi0G71OVNCSrgVK2Nb89nF22PD
dJAx8gCrc7DaVvuwVihoPGPS1JbLwXGEDYQZdip8JJ5Z8KfqW4O0E+9wDa0Z4VSw1992cnqJPQuJ
d/VVdmd350W+/yk6iI2UgAlNdV1URdtSIMtDEbo5yLCpnPd5UHeUhZCqlxqB+VLCknI4GTeOikl6
SnnA2GDS0w65ZK3jlq709Dthb/DL+iaPPyBYeBe1bOA1icdiMwBnHiqkvsfQnZXzoCQWUzGO8G2x
OzWX70Oj2fwJGwURV3xYi9FLPcW7BY9YGmxq+BHUqHuaYyVABYCIpJiUfDdDsgIiWFtk539/uXHw
ZweHYDkShcpZC8FnWXSXzX3h7A69U4T/M6C0eSyoWgdUz0j/wkjR4BsdgfPtwzJ8aLjCFwZIceCv
kFjDJwO+f8UfikuQKvFNqRHMy8Wt9vq/8tfwvKhA7IgTav+0W6tdFb9Z5W/GniPQwUyGrLIw8kxY
aDZb84mrXaS2eIaA8RJG4B018lIS5YpOBvpgrif+WaBheKbuos/2tnbxrGWfL+K0wbGbZqKAdJom
QPfKzLP8CdXS150EkoclX47mA8uBqz+WM/HEOPjOLaGh+8TQWoWwfaKk8CGQgBpZzeVrUmGD4bTr
w0XMjkawCxQ+yK//D89ebChgNf+UUTQY+OW5FB08P2flCQNro9OL6kQrqrOrheqFqmx6MEJZPYG4
/CoiG1wXmeAgI+gecqBHTF31E422TD1TR8rnvACs1nwX7xQHfdaGWkS3bg093pF9X1LL61E794gQ
AWPlQGGHAnKFx4HPmzUDNSWM4B3GHuX3OzXI4xN6ZnnBgRomOWnkfQU7YfmXYzchsU/sLBTxepug
JOEIgShOpf3GukcJ1ihpYUA596oJdtpA86uBirInK7MRM+v1XfZu0eRrnKGAx2iEAacXBv/EArX9
QbY93hflrIjXpo5vq73Xoq7E6vAMcK8OljL4LuzIsPweq/FjtyTrshMRJ9HJAMz8UGafKXQfA0Od
MHBD01Y0ku2GiHa3itvNfrRcdMi1IkT14uyB4dGA2P8AtI2RubyK77EVaV1zmfSOuDbCyuSzLBCb
AUnNcQgA6DGKJf8yiPsO6ASKsbvGYCMrsKrwatYkRDOeZgq0Ae78/qA9w0akLi5DQ8zTvbr/i+8H
+e6k7g7X0kkNO1ncBag/FHOBSPVHBbSPGrNiC1otkY2CYVzATOxOCWEFw4JfUyCPdW6M7Ui1JCVO
qzHbIKedtURorElfBruhtse1bXMO40C3FnFHt4SqfWf4g9rCtPP9amLsOehUAnww+Yz66JgGXsPp
Lq6NLW6lDQQ+apjcK4oA3pGkFMaKlEDaQTR1SY1zqRhc253HZfBR2vlV13uYj65/Xf2PSVc0ClEK
IDyH44BGE4CB9UhkBILRc3DQIhlLvKz6H9QSB9VO6pjAyCjbswtEE4nKuI05HPG7IbDlfzxmbIO1
t/uCKDCCCaxEQMJKRgX8ttTSCuyfDMw/UpjbJWyuIF9aNs8U7g43C8ScbUUoAngW5ZG/GBPYhE1r
ZPKrSHr5xuQrVq568DfR/lW3gPqhY6LwjMDTBasKEkNDs+8Hyjt0O6cro/4ALllLEKGlIaH+kyyI
NnoLm2T4v8URlQUCHpNzyYB20haNyQ9eWTGQuRO01vnf1ab11gDGhqls4PODvhZ3WexopCLdWqp6
Tf1alQzapHA0HAkJ74V4RWjoD4/WR0E92C94YOqSB8W1Tqihcrs77pi2ihKd+KGK7OlaMhx7yNeu
Ry2IPKhnHQpicLytkyBAXvPM6JNRkYIBiSXYzd310BxGEQdxqjs/+joj0cmg+TxqOfWRGCAt8IL3
6seOtM508kitIvLRm6NzYlU2vYvkkj4Vb6bErSjPGrlox1AZ1R00yqQmWukbFUdstp3zFZJcQrer
hGgyow5rXQ2hsZQTBaHAShiHloprKnRRaVMo/rdxAJ4pQPsY0VBv6Y56kg30wm8BLigbzC7rAtHX
vypvhEqtjQOwB4Gn/zJU//zDSwWPFXthsF/AG90UMVQIQQSP0QY7Two6oB+90Pw3PMiRu4qX9CfC
m1vxODt2OUWn7pIv+CTo75/aSYsHi0DccNVa+HzgRoVOUweQ2b7aEW971mIv0eHUgffainZ/JyLm
4uLQgOdA96fV0lNwVRc5+B8B2z9fRra3Rn8Idn4+llzHiPZSjo3NVYYZkBGXb8JXv1wSEij/7oi8
VmdF+2M14/zNJB+4nV7JtXB7x9b/mdCLOX8uVHodiSydc92xO/+1WBkh9cZKNdg8z68tmHBo+4Lf
0BQe9Vm0WxfdpMP2QHwfUYCtHyCPENvocBARfZ/J/S/6UAP4M3Nu25uFuJU1eQs1zPCQBTyMjDlZ
OD8dinS8rsPGeBYQpK7qjcHJfYI5birOAEolUtsNg1Vt+CkraP26bNHgFD4Xd7AwooXcHYV8h1u+
+db82kQHbJEhGcOfbUXhdxbvwA76gKr7MAZevln7TwG2RqmRNra31nVWw5Hhxz76p4avs27ytowz
T1axqwmRhIb8Y7pjd03ot3yvb1TMeo55qxJ0qaPApIwVz25P2rFKeATt3gdka0ximuSZlapJHEum
ckV23X5dNfebaXTYBDceTgjGCJpnZLQ6JrRsKIduKNBQHD+NHQQOFCkcbIqPbEWR2CuGZOe3nFWf
O16H9MKbSbk832Hxw31gysBK5FhpAzVcdj6DrRLAdxkfp4FmQhmof5JSzv8P+L5G74DPdmDcpHup
yRLf1LXdVvVQzu0Osb/qMi/CXSFOeFurVAm1gVrto3jfbzBN4G5E6ocHBAXDj+jnV30zR14FZd+h
yzhzl0VsuM3LWsgepJ7rlPMPmcETsyl19ezh4V+aYD+Xue4gwUkgV5ChvJ2/jsjHXQMoFWarl2WF
UIuh8v96UluBOSd4NqEXh8MCElzabmI9CNvglIjrx4VF1OzGj5k/wVi9K9o8QeJyQJeRiqrsDKLI
ksV21wmwz9H//z0fgzVTyW6PUlubM+nY70vHkZ3J6I/MJBxOp8S1k+wmMQNMiajcpUb/kNY07zAi
Lrj/XwA431jJHxO+jilXy0jDsHnqCN1d1lV4KQIlFa5S65UVYsyMLvujHKmFOitSPqZlrjqd+4Nh
+KpMIlgSuEuj3l8F/9TzMo3Wp8XEDKGnL/sVvcFCwdU3jRd1eM1GtR/0kjIRjEcQtk8mc6NQLheL
jjE5l5TWAOD9pDF+x4AMMUUccFeabzd5lwezWJ4+UXDDjNeAZ9VvL76i4jKpZfXIivajGBGzWk8O
riM7nROZDebdC67MNXAbGoBucRel+iO2Sc7YcHjQAE4HyIHjaqqpBuzMRCGU4rs4zRYH++KhLkHM
78Gc7ugdi/VIZznYywgujXaj1IdUlKnQzNSk3HgGeknNKdHUms3rWm31bFdzwq+igeB6bsZPM7ES
8lDKb/JhIb84Umb1BVM66sMSI0AH8/pZ0JvbptUKfkxmnCAZ+F50ygRzTSGvsmY9seZh2Bl76k70
NgGUjI55fsZlIzv7SaB0qX1hNrm8nScziKmrsjZZO2gvaXQUXQm/XyJl1URixm94AExx1i6n6aqb
Ku/yXmkYk5UbyDQrmq0N5Y32iv5pqsRhUrJos0MpxQnt5g86knC5gp2C+mEl5ZAqtt1oGTuGpPGJ
FCklJgcuLac0U0axQgH4s7dZGQ+i+sSGIk9A3VBRj4GCiKSPLZR9+wtHU64SdVbKK5J1ZRFvAzNj
w1SMeHUQkidhaG8nNDSFp7HzZvih5FBprANowghZgm5z3+LS3LY5Isax5JSuDWiEGZRGq7qURq00
dNRvOGltIIi1W9SAM8IscAJ7LUgeihskSTKV/1ytMbd5TzJ4ikDvLAEN085n4F1IjwBeqEyiXZIl
PIzT5s6IH2fOlR2w7T27bm6efM4o2Hp+u0SGDEMdAsVUWsKudfSSMX7VIvMITNhP4TxeXclRMbpG
jNeOzC0eX2V4DA7SZYCZepd9KWIz7yeGUyGU1m66mPxPApV5YtS6BLuocWjf+xS32Xr4x2tNIa1e
nzrxBiQVynQ3I3fSaSHzP5gAL36TPJtN3M6WVlMjTachJjyc4gpzb5jTjGZ/mrOhhzDzO3U9XOBV
TMbRXFdhNeteQvmnJ+BheAGlwWUDs3oML9aa1Ae2nji2C6uBMUXREgVNvtrk+e6WOzwO44Ux2Lu7
9ODx+su0ElIbLquGv4stRXN/M853isSojnvbRmIzuXb7SFMT26sBxQhfWkWGkeUo4eI7hY9kxAI/
F2Myxz+9zCuUcWDugMKN/rEUh9GMaLnv4+Rnsc8KeFR5JJjHQ4x1HYfAwZ8TOW2/37OGswvfjZp/
PzAKBKQM52n3RK1eLgZLrIJ2RK/EgakHhBWmoXST/+Bg2XX0GZXw7kyENNnZN5C94fxbm8RwkgEC
8QnwMsYeSMLFVomadXbjq6xdUxyAp/3+2UJ/Yg0UCn1RQU4LgWW3ykCCWVWPeayx/02C2avoEyL9
A2kPMtft6dmdw5sAJISKl5lAMCctSWwFZt22DuOSlzJ44A6wGZH8HQCzUxPK3OGSAgP9+r6HN89l
e+uwgrU69uqOVWn0XqJKehNwvqM12UIlWtQA3Y0/ngfOWdQjw9iGl1rG2h//Qc9TY3M/SdP4hIy4
cCW8jnMWohd08KhwabhTIgnr5eTsLBQXe8KwgNeQx+xpIkMSIV6mmQt5SbRvsL7d1DqLkM8Ef8Bx
bzhlRO4lduaepV7dusOkI5GD84UL5HltIB+LobOjQ9zziNpHf+k+lW/DXQMMFRCduf872TtgNTah
w6/5h5iUFsO0yDYBk0lq5KRoRto6nWBobremWr3rZ8OMHUZ+DFYr3FpZ3T6+xR7J/s06VjYcUfB8
SIye+QUFjE2/UAU4oYIzc5BKdJ9+7z96S+PdsTHwQYFJwynx3jgBqp8wDFEhYFXGuAeaIajLW+7Z
22zkSv+frs/suhplAL1WAbTZ5CcS687gBNYl40ncBSK5UTP5GIB4wVkX8sRL8CoGzDFApPbcxirG
uixbt6KE/ulHZvPuK24j6anEykiiLGKwenV1h51CEsOUApXaYsy5tXIPv43np9paCDfCjtXyjVmS
cWfuWZSTFIpTLgml+Sbp6NF6Ff6xbecUIZY9hkDBNP6M3nM1TgRXB8pE4O9tXTRS6QvS2Gne8Pho
Rh8JWRk/5I7NZiZcg6Juj81NBTXFWV9fZ8h/ec4m4nmje/C/+JtZHWN3xIX4MwDXp70HCnz8YXIH
IKZzuCcroqsc3uFzRqJNDcjLJQhJGhJlwaRQj86deCCgHpnbgfdYcsU6aRsSuJsQN4JuCm0EZKAk
7kxXvAIqKIrCKWkvvRy50a0rVMwuZ4xFiRZ/DsBdnhy6wTL/gwxZpkwdNf6H6B35Cn9EgJwFnGLv
IPGAOXOIXboWm52gLWYh4+OED/uBcbM7SM+7Mjk2SROqdbzqn/wi3VvFQcXCwTG/WEazYSWIkuk8
U8UJGFb0EPKZb74xlcpgqig/iRR0P0OPxbDtpJE4JtJc8qE8dk7IUUPdX1Uj4FWjkqafbx9jgFTW
TLmmYg7ed/oEBF8246Fran+41Ri5+GlgpNZOpEH9hxKYg08S2UPXG2aeeKU/cezNbRu3ywVfkxtg
9LpqIh8ihaD73yUWougNx6PYKGidwcoSAVdLssXDE0ADsfSigXMlddwIKFS8gri7YPxSC/oLzRX7
bvxtB/TsVPO5jlZQFFgH6DzrhogOmy97BLOUDyCe2AWuQJdrO/VbdC1wWv6xU4eQYBY+k83LEEAP
rD6W2HJdYN472PP895d1+tEhOW53PRA/aEVJtxEXP8SOJ22ZRBUpho3mzXVLaM5+Kz5wQXvT90ZT
pFh91RwlpKukVejQEZ0RC7HijySdEXoNlGClZsE32Eg45k8NvVVgJZOgn9kNvAyzuOQBzkHy3QCP
TNtDBEKk/ouAPI/CxrE0iDFpcpJ1nrXWhNuKMPLD+gO7udOT/8wC27dnFCI94kSJ2yi7dTBei4/b
oCxmJ5HwgmZlbYQJaBOlJXpG/eALXxYiGsgWNAMuFPqGmGknKyCdgdmllFUjrEPGCZtGT6Xob8DX
9AHkbO16lLOGdSNBTRyKv2Na2SmT79qH3ojuXXGmaGaZQXKjjm8S3XFfg7C8EOCDTcUeWuRASO9R
Sy52cOCVXpH78NBt33Skczf1idy/Z3QEf8emKqK5lu8/pbJsREK+zNwIEr0yvn8QRhUR/8lmGMBp
W0ZVSRFC0OOE+XPeMZUIw6IAMjSxB53ErHZaMGJ/+aJaxrHZq8wOqtNhE4xYOwPAB5lcAAD8MaTJ
g/7UmwKywP3xfszFZW+sxGkRJ36UVImJOotN3J5c6ZPOTwqKrIDgittNjmwLFTPzrYRf0daCX5Pv
fMZ4fhnqvYPcoZp86g+vEb+/p+80fl9SBjYqrPIYl3k++GvU9nKAfR4zPZWD11CQ9Y4/g64N2NwS
fdrt7FPx2190cbAkZwldqez5THYSYGM2dq9dMdMzAet9/6n6h8eecaQtB7uOESv0GLKRDr1yA3UC
kVjcKKb1BW2+0/2hDKvocB4GeNaOjRW8bDs6qq6UdgCSFdu2uvssXkFhm55h0hzG8yzKOQhoHPIz
iPp+v+w+DMwaYTAbB2bpZZwNCAvRrZdx2eCNmQxlAjTZ3tBydlOvq2QUX/Qid8Se0JV89Emp0wY3
gwDAkBv7ZMABeJBj8b24AJULSq40at2Je6y2rnPaD3pq3FWP023aCK8P3CmdlGWnDeV022ByaQJZ
k8+V/DQOjE334bTQhWX9fUKslZ/o7NQJqOUEnD574GkMaciSLSkMn+O3fnLODI5skPo+LshKj6EE
YWwER5dPM2tnaRKkSF0bzvlKQbgZ4lstAmK+0JhPMdQ1BgNcggAy0CJmNx0dhjvwnmYeNope4QjJ
Ea8piCMEepVVmig95WCv1Hd3cP/qaseI+HFEErAIdG5R3Vj63gkxgoHa2GGHhZa31zr1ymLciRwO
+dVZk9h7xwFaDpBFA9Wb2zNHQBhF8DVLqpsqSE5gs1pb4/TRgx40WNzrPx5RR6EjOf/RMp2CEYlm
D/1no7/RJdfmPDYYGGywvdQGYGVQ2wVW6L8DQmYrCkw6+8hyj7CnIJKvwsY0+1VaTNMJkwxc4kKK
EvIeTV5JjfqSq2DTov0NCu6vIWAV8xqyXWChaoPflYRjAb9tM+P0Rqtj1RVKvaAMXB9k43db07wi
cF0aR1YEjBKBtl+01v2c8HRh3Qjsa8NaZlzM/ZCXvvlWdi+8aZ/awdtfWnDCwRG7wDhs3Z1ycK/q
VV7eJyGXhttWU+aCP9tkIPiM6QrY0/8Z5CM7N4fVgt5gneH3idFPl67ceNKc8tboKgMXE2Vc/0O5
TAzePD2mXsouMGQ59FePh2riD8HZqauw1Nc1C7eL5ibIoiftGLzirkfgBJivwJBDtlnmAR272h/I
qejlwqAl/w/vHa52kq8BgZjNs5KU/5diVPe4Hp7f33Ehe7EVN3mtR7T7A8db+V/qurFFpwnaOJ7g
H2HnCxDfl34a0jP5k1Vivoj7l9UwV0UXv8urKDDUbF7pFedh/bgjmU2bMwz1wimAWXZg/eW0ztdX
O6wSgq/6tgprSsUS6m9qD5bp0zJqVZGAxRAYyShMFqud89Qhw1Fs7/W7O1Q/0xp22OmKC9VZFMms
vBtscyS5fBl68CuB+kUm6pNmEPjp0Il715h67/kteOiss/2k35J0MhA21ut8DTobZMmqDpPHeOy6
f1+y80k8zlAQIZ7y8P4P1UWT+G/PY7fAG+zBmjjgieN3ygFFZPBsSY1wrns9cYpPTcHeMZQmqRQG
RjwKVrnMR9V17uXpqfFnKfl0c8IsULXPRFk9rfa+7VSzwHL27zcJPweO36TnOb98yhzjZGDtkg0y
FytT6nBO5TTyLrG1zOfENpUJJZgQpo3qRb19tXwUbVh/2YgQ+idDplDYrGg9veovyZGzMWVsQn+D
I3/plpuXYvKHtZyyn/N8Je/lLWAWo48Nw1jkmUoBiXewcQe8bJxosoZ7kGLNrJ0WecDzbwRDmv8H
8cwKpjweeqYeJjhztMlHvcEVdDI9PPQsiUrTyjOt5o2f0CzkbcjQI7cfH5JmgHMf92XBnXEpMFjZ
8XMnGKu4H2fR6GYNbLR2JT2+X7IhEC0uNg/TvbpwCTEa0YnZoNSpYPDCvwdeBVqHAijbIFu8hjOA
y4KBUJZ+9UDT9zn0M1y5pPAexgpVa48Y0sGPnb+cpYZQ29LvxCE/QJc/L+7pm0SeQq7nH/TwI8fD
EFJe1HG9GaOO9qtfINO0IySwxGAvAagAEOqf7rgFD6/gSdlMfbc0ZWm09hHuOHLznPd6D5EYTayY
y9Gd6o0IXG2fMBMVMn/omhCsOKN964tpPhhDHT5j1Ilhf4xAAKMgk05lEjSSOK2IRzOX6WpQUK6i
LOfCXNGu5jJFW4iXrpM+lQdaorlWifXODGB7vp7MzvAlADWdnvwqA4TB4A3dpmBbWQPcA9PNWzH+
UCOXO77CFun90GnrY8hw9p8fHTNn0PTfqxGSVjvF8wmztIUhC3WtDn31JAqRV9QdO1YgQdMvRN23
C6j+12mdgJi+sbso7DYfBWohgC119+9P3FRA3wqcgZYgoD1mRdHU8dXzwaxsWilXt7RfeEx78s1m
F5p3Ih6ig27vVOG4pvgqjg4j5C559bE8sIjUreQe+TAdTxVbfO9OCIo+VAuHnsX8UHMu4ED/YgTo
+7jzkpMj1nKcUzO68urRipX1cZV/q3UNUP54BJ7oX8lURQUvDx5rMEq388IjAYVAkSvFZs1do2k2
MdjdnA0+CEyGe8Z2rLcvloCuah4tnmmg/fXNEaV3g14uWhw/hWoIcfgednhE+YmsaB37qpE15Nix
CLx0KjvyCitieScZCOZZjzya3toIJmtbhTq91E0CRD2a/HwWl/dis8CnKW2Rj6bML0jkQHgNtCT0
fmNrylAeaSWjLRQCzKSHxiA0WOeTv0HBEEeiPWmBoxp66vajE1rX6SKy6KN1q1VnvLEicIOOHWpJ
3t8ns6pvir+no1qmEOyDwIgxIihdtn/0D+IDWyQKZqRgSowrbU16cUPVoESVx64nvqBd1RMGinRI
87TCBMU3g4dmwhyeF0FKqb9d3pHzaotKrB5ygxNuhSUcyNTc1eMlv3LyOHGheEnFApdWK9dEBKfb
VYjKGOHVKeVRlFDgSlCHfHwnDvOr2Y9vUQvICS6PcbWJ79LwmIqyas4ZbWe9Ct+QehA03vFzlyT/
4b5x0SwGAhv67LM2yRW1jJrxqIhRc+93p/LGzmdVZYMxOb+X9298egWElKiZzPRatJV9Fgu/84Dv
Fda1Iz/eiH3DEGIUCF1zARMj3Fw5nNppJLsQ/In7btnj3KmLGAFf4OIiejbcPqKdzvY8lkAD0LkV
K5nvlthYPJolbpVMRrt8NJYjmse3fel0QMc9UXoIMKyVUMSHueDv2PMazTyS36hsoQwQkLPwz/e9
ihl4LExwZ3dSxf8eZ+sPAZIa0UbOspjZ57cr6vVYDJRsAc9Di36AzIGq87rHAN7oBNmHjFF0mWPf
GiGvbt9C+ulDl0nHKuSg8Wls4NijBpxY5bE0FrwiboG4RqoschPzeBMeTu7pkabH95QtbFSeYNEn
hHUbLW2TgqD7jbaME5CGYjUl6I13H5gBS7bsPfO/+q6sWO8dKmD2AFhMNoRCZZwbfmAebcEXB7CV
+Jq1qxQC4d0MqvP1qhgtHHIodaGsuGcYhRlW5MHXCtgEV4VEyxEM5ZloZA/SLztiL7rXziocFl25
dNQguqP6jncAkkuCOinLgbujE+uVHAtUb/Bmvy3UfPi478tWsdmALjg+Zwik/IS8ulHWXW9q4sIl
VSek/Ukez6wrgWdP3hwDBW1efBrGKrWhdfi0fK+GMFyN+2ay/ATA7WpneaR4L5b34zp9PIag+d8o
yONmYxGanHqzgfRFk5IpQAroRBXV6Ioc12hbsMPMwNZAT5paqi4pkBQBYmF+iqZfjl215BRNa2xN
qMEi7iH+vSpq4l9vjYM9L6L0JHrSRsHjxDK62z4liMjfy/oMnPIyTuEMp+bPAFA76lTyEWHq1OXd
K2v9+orOZfIWy3OJ6v+g6Yt9fSpBucQQ/vr9CazER83axECRI14eQvQcnmevHKbtcoFlww7X9Fr1
KuAYm5TAKIm63QJGASm2iuCznx7Omlom60IdejOu5hZbJkxUO3miOTa4IG2V+pFCqWFjFMLkbUhg
amGOcNUwe2c0ht4oPyp2cy8UGUX9J5RduSM4N25Is6kQdKb9VKqkXN+P1gYO1Wf34rGdJqotZusw
Ch3qGv3R7gyaZX4chOY4NyzL4h5l/bwuDhiIKdvTV1ifBljORRY4w2YTl73KeedJ3hb9eXOmMgww
FLHOnhpcuaQpnlmG5Z4wJn7DktYr1RV1nmUo2NO5HPT1nvR55C5ON0XbuZHpL3s0jooQyXJ35W/P
LP37KjUNdToRLe4RTnhQZkDZGgBKpdlFEzGM54pBHlgKy8LF6v/MTPIj2qw9XGEp2V3EsJAvOARQ
/KejU8tEf1GIQS3o4P6MWM2dxCjq+p2igFTsFP8AgIWWbZ2GBpBW6DbA9I7BCh/nxcIMIwKWCh/1
Wr3k/S3U6Bk6iXnbHKMCyinTQGUGsElKUN5zoXK+qiqGReGBx+ik687689QCBdnp5odKxc7+mPnO
A6qLkrV/pDMF5q9QagvMTfxg+WFC9q6RkG2X3xPLdPH50CHlQk6wK7drTy2UwCm6rUT8aOWxvN/Q
4Wv7ZnoEmECqK+i6XfgtY8xJEIVEeVyQ33UqpZZTxOO93P1wc5u06o+Tdo6R9q8kApF32J5XBBAt
MeJFcCD8ej/RZIwTP0xy2Icdd4THZLvIQrdwmbzfN0smFrxZ1R4Y43/NdtNiQcE5vNhw+IAQOTx4
bKbdPhZjr9j/1mDg3E3UUNHj9XXNnFC5opWiof6idn3TEGkD5F4tsfBR3XYk362D1EWAG47J5WCi
5hswNdTGLZDkRUocH5Oc09DJ2npr4CqSI9zi0LpvuHmX9U+bjAaT/LN2ohCeLE4YXZYCoaXZeJYc
26LbMrkzojoCwezGCDYjKMCp5Lcl6QRFF4oeQ1XbvM87JAXRtJVG5+8tLfy1gJTBmrMh0rO2YDxi
VmSZgocBYkGksh5QhEmtOr82gTc9aKorAjLhFuYmE+vjkBdY9kn2DDCGbU4DUg7uV+NqZ8iqLfZc
HqNeb04zYVRr69A51UizlBv2voWN32xYEfLQxuL03ncQAJ3DNgCm2A/GAbrez6ctdzXAF3EXRK77
Styu7J9VXp7MT0V4WmJaRv8Ku10hIsSggYHnRUom9iQuO84OJARJb3fAO+CNYFC3DBq8BAV27eLq
UGvwrO3b8A6eaog6hKL7TqssvzN+8FvuxQAFK/R2GyRBsMkRDshDZT01zgrFTVdqbeQ4gr2Wqxhw
Vs5OYvj6aNnd+0+9VVaE8K2edcCWfCe0gvLAMaM1czBj/xBYR3oyUh/JDx6Pev2JgbpWs5Py9d08
6a5WlyyZgXf+HLDBAT9j89kIRGLHjH+iJERFOJLPBrsWn00Zuy5QLAX1lj07rycfbV9OpAthyYhH
1sSe19AbIcW7EmrNyqcpPjL3qeEeJxdF7+jPnvXpjREcplmPnXIpe/bI5zEfUrftkd6vohND1W/T
2h75tHO82EeiEUo5/3zzcQuzcFMBIJj5bWp7o70D6ssIowmgKKvkn1A0AiSIpykwikKD7+v7e5Ff
XcMGWNJeKSuKfBdU5dbAdUnsbrBZszclxvv8oXJyUduUDLsndHjYzXTF1paLIJW24gKzxSqgL+zg
2Yq1RpagJm9WxbNed1XRchf4v3QAP5mQXm6E+92OOUhK7QbvgD8+YkQDT8Mi54OqKTVRx32BFV9n
WrCftRLq3IDeU+Gy09+uhhe6Jj1Rtdtt+wBJteb/zhKORi9Oofe57F287TuoibKUqOXpo2eovvi4
ZwOYSmfpadkMoY7KskJ4nuh/y1/eQhPl7wA6KfXTgDlGamDBTHWLkqrNJnVg4CBj04vlEy0I8bIH
wpe9/aCsOWMLQoFyKYkfhqg2ciQV1vinTgssICyRfkEiZ1wMFYSL5fuzWwMxMcrhAc8Tba53LUgL
JL8WoAaXaQODrSW38GTpCK1ODuff8HMSfWgNr2IdWdcmuB3LzVL++SJ70MfVQWIUqRFXbdnmD3Ev
aKfV4rvThPIs+VdtmUyL0y3DIKaXxL8sMZAeYFR/CgkARJeGTckUZ0ky26/hTP/+DSx5+YQOUsFl
iT8MbapOqpOApX08+qnoPOBDAc0Vzh9/qQKNMIltR7XFUrYPD8QfHqs7zp7IS8W9PhdZ2mwiHyux
nKhy+y46hKyH/3bnLjpU5JmCpFrNPoI8Lg1Cep5JFrp06bUnO23Jugwsk1gNsdFK+CAM4Lv5UtD1
3qZBjzTUyTXDdvCjBBPYzSPf0RaVUeFeBkjs7MGikKwOcX+ly7QpQYR11aZkrId4WEfhJKXlpJXL
N+mmFIYbyFEkRr/pcpzkyHNpC7v28emh1DxvmaTvnHWRIkm26D8IprMPIDzXTEUWzPS7uONIbutq
Q0KamWQcFrCY4wQEajuqIISXu0x62OMFSbvBHaPIKZLMVy7C85DrwL03gBrGbUxZuSYLcCoYr65t
FaJhHtBh+kEXex0UuUh9rIjgSzP6Rd/p0q8uitNSI8XUOsoacTJ2Dm2DrvF8yEfK0Qj02PKTkvuN
k1r5IR1IL1VUcoMsMzJrVbLPaIh7b6VzLXRvqm9pCO2CyISDM1yieytzHN7E7JWNx2+wWMJ4527I
psD+ur/JhEqhE6LqNSVP51F3DJVVZAYYfW5aAHjYtVsWxBR+6Men2RC0JEY4BheY2gMSJR8EVvsL
nwSXyy2GC+o6z5P9K4UUSb0WIgfBypDpeT8iVJbiXqCpMPHhQqw5MGAVWRKbQJrYkRMWWnWolRZd
vdhHpEY3BF0EheTNXOywrIs+VHQHkSNBf9RWOL3w6xpkyKtIwkGc25sQBATNwsXX6g1irO888w63
E3aGd6X9cslo/GeUFu6HHP3FuLnVP0Q4qkmQfTOZ3o8o7EuCNqeA5oDlhzZL9Kj6cq08awLquZfm
JvsbNOlwVegz35nYUpIaozOAL8vcNKQ/SVCld/4Qvgv5/HMM9b3EuUPCGESKVJNsFCSv6FsiTO6e
xpWGRPhwFTOvZmUgIviQvdN5ls0JbHwWjPc41m2h4h7dTQip5TIyI5CZBcnwJsnQrOVW+ZkqhgXp
5OQH/mFF52vMUvfG1kmWdWanKnz+zwQCD4EbYiE4i86l0tolRxLJeMlg8yGtih1qD9CwBqwE4GF9
MRtsgGlDqwksbcA4KOU7jTu34/8XOD9hb/g0HE2L/Gza2LB5OWo55o5oEdMq+dW+qAt53H9/dVt/
DfNJt3DM865eCzbXmk394QyU+34sUqNXLe1P6wXcxD0lJVebKcm17AtHHgo0qbdkwEzvMU9JceVy
OerH333ICK7hvBvnVkELIkov55jHndxQYVU1qbHBQMYxYaPguLzrCm0wNVNe5GrHUx4SDc5q8u78
npj0lgfRRmJYtU9efZRBLWHuHBLjm2So2GK87bfg2YvJcwHG2kg6ErXBK9cvkRnR4a5HOeePiRJf
rlfPxNqRhKVeiDAUG6UfZjO9HgRQnvnNsq8U7x34QORHk7/2ZodSiSLwe+tkLKXG5zTvmzU9Guu8
fjHn0GOs4JqFWo0MnRD7KdEMymnM6OksiXc2LI7VdNNvz4ZwaUy9Ol9mbivFHtLpk2jn5h6pf3G2
OGMYvKx84EhJLoDfSjzxBRDexRCXuLFudOMl+aNOISxnKD6i3eykAvPxCbCciFjzDhZZqug0ei0i
ABuOP4aD36OEhni5MxqjuhcDC0tdONVVwbao3KIcKJkVr7URlTkMxI307kfKpO7WYn9IenLYQ8v/
ETYchIkgKx8i6ED8QoLhULWWwfvSc/PPGf3adNjkvCYB+dBI5ZYg+71Srrnb9aUu+gKftvrqd7UL
Ac3NK18JgNufGLQYvYA2gny/Jw+uGaXwjj5GeC+PoTwTWYZOyO37RdeOsMOWaZKVDk+4OicG61TL
BxtnrKkJzLWNYITTTq5IWT4dMjYChrbVUSYePACpRox80PgqVaiZt0q6Oulj+A9eN0oCuz80uxl9
ZJ7+c2UdjL00aZB9BFqdMOvs0ufGacGBkczIpebAG8ShHoLWBKBJudDqD508xXMyWsT5EROFR5oG
3Ptu9JHIEXvCA5JYGjix6p0UZrxMa0zY4avXBIDR2ZQyiqQoPpN7ySeTlZPQfqabws7Jxpteht84
4EsYUcjSGAcDoMYxdV/yjQM5vbrsbbaSTNIz5Oc+EIjuyG11tO0reoDGiiiF48JnuWjocZjNfNhN
YgbV4WCxLe9ExNbEFnr6yqf3stBQT2yiQLKD4+VrRN6naf6WkCm92cP2zp54ytr40gjcpQhUsdPQ
rUdcxJ1+wfoVIohH9Xg7DNbVVYrFdEJpTiSGnyTSAvBuPennQmNtm20A01f8+u8d1N92KTUCkxzr
XATOOpD+d1qewkL7JHENeFH4ZW5CyKEyjTRtLHrqL082UXL6bTU/1C970ZvMcP8JvZAJKbf062dx
cIq+/nDWbDgEluvw571gKPnRBuvXkvJ4rKinRAWIr7uT2fKC8ivMlWB7x4P4DWLLw7fpaDgSna72
W6t0fercyDpSnh0EAhrEP+r1VhgUj3GE3q1Ob197DF26qhR6x7O71XZ1r+gh9efMzCqMk1ezVzuz
ayQDCsOEILMcKek2eXu+3v+EFw/9VNRDHnlH5sni/reNcDFO25slv37LDfKbGfHe+xi6YmP0giAE
xg3RfZh63ciVxDnHp1KH1Mj/VWxeNrA+u5un8s7WRweMWg32/YGhzs3tKbex6ZCYy52A3V7Nvsct
gREMag4Fk1qvKFXil8jq//Lh7cU1TEy06U0ueVUWw4dpChYi8f1N/uAmOh2/OeO7Gymbi0jV5kLG
+i7tWLAal5le6zFmEwAfGvp7+DWOAVZ137qK9UMQ4livKOlbCQp3zfJRD/brBLMojNaMvC0GK7Au
6m8fYdBwfO+W5JnYNOwS7UhvYDKyyE7yTPEyjNY7m5styoovblU7J2veMVbaXLROb/ED1RjAjT97
5eiptdKZLN/kcLsdDt8DxOzlrpSu/J6pM06cJ01uov/mZGc+fB5l/xHWNAvlcFdIEZoQuHW5q6k0
ddY7yNof+eu78QNh9dUltgFO6GT/f4wsxOvt2zhTLcND+dAvIl8Dfqi6FSHbelLCkaqfZ6fNMumQ
8KQ/CIs4mpksyv6J8Db4AgforAW5xi9qOX7NR3uP5bzTPGUnHLNXtE/D4CNW8WoVeGWZPLVs8WiU
dTXe0BQMOv6rt8GNvJqTyldkytd5gvTf92BPirT1XqbZWKMxGapQC7BevVNPCGWxBAuE4s1nXKWb
vfYZHDxLBbbOE8cawvAHjOosxmH75GEj++QYiLZ4/BBw00ZT54f0Qt1unBMx1ObaRAUki0e8LNe1
XSeMnjjAL5Eo8DuGiUtSYNZeSqlrTuXgxsFzz3exSZAG7IvCZaDxaFXkiZ8hQo3QICYTaNROXa8U
XSoRlrJCzDPUjfcTlJtyWRZXNP8May76WFkueYmQlkukgnnlIMCJBUqZ8xenBCEv4HHqqwvP93gB
4S9v4LrTAmVLaW5CUoIkFBJ853fNdg7qbCYa9RZho/Jk9W2pDTi4CGH7SK3H6QTsl53FO+Dl0CWD
HKDHSueiFJHfGPobw4Cj3nFg5+/RjHkPYKiLJx+k5WyuklQ0jFknOkeNYzYH+wVOTd1mlr3a+iAg
/lS6CJ4uj4VnFQlOFrWQzelOp572Jquy0wXdtfKkGikBbxiQL5DmMg9DkJdoHQavoK8CbVlOPMNF
WKoaxJ1h4pfytWNtz73Am3q5a2lBS5OflqcMOASBrfhPWxWdLgMzvJ2fSddNTEjstYr/igkOEv6K
swcsEbbI2x9WVE/gttzU9B/+D2pFY07T0mG9RiOrbaA7pQZO2fzkdsPKRC/5zLcmcmOikdNMzwnr
n8mV4w7vgHLMP//TKNVmT6+5/TihrpwFBQy/gHUtADEx/WBuvGGE6WDiuWgkzoqWRQiUT0ns/5f1
jCupOs1VHgkdZSffrtKX1+UEjUsatpIJamYxeygDsA+DWD131C5waqqsZcueNplilydE88+B8gz+
t23l3cefTwyCbl4mGyiqpFrtl9zuL+nY7ML27NIMTSE6Xn3xkWSxKWN/Le9qaOFL0DKbUnYb/IJr
n0m0WWi/HMoq8i929jww4EgISn4eSnRaa3cKgok1vb8XvL4OxdHXWsTD4rka6at/mv/BAFCmh16R
SDuGp9sttC5Tct4mrGKfqbqRlUOxMoSJHqEL76Qk+eRiq1Rq3kT9VmBmJCpYMTGW/+xCvW7UT0zt
dfkMbErqNCpzHGFU+GsrHVYfAAUqNiiBUaDCGcgGFrFRhrwJXIqMBHt105Zj6TCXfGfDjdEBRYZG
PDjS1LVc45lhlkR+BV5mZijPuyTv49KJ7WaPKKdz8ouzxf5bxI7/hjT4otex4AoIQD8FE0EJI7Jj
mWMSJ0ZCHfijgdDHebSqRfIslQX2bHJtW/VI7yHy8QOUZ7WR6Vf+92/z6kwoIUJirrAG+MUWHcfz
q9h2rWXGHRCdg19OXgf3uKHHZsm4HcRLc0aKxgXMC1NG/u+2JM2eUMLzDk5ChsyQ2Z0lBy6FtG19
nmFS7kz2zzhC4eVo1vbs94SnT3rp6WiawsXvfZ4tuZeE3/QMjunY0Jj6rggbA9k92yUR+7zQeVaC
GxoXbvRl512OIvxuykVMh4almC1RaZBNKwSR+COcYfjAUL7f9Y4mGqHco4HGXVLLztVpbNyuo0mO
aNK0G3JFAdwM+nZFvNLj6/DYXBYGxyniGtjI26jhubGn1DS04DyEbWnKoHAxh5cBucGXAB34PRzN
WnvcPN5KQqD2vewvFRM2qVWsHY8VzUbKOGJMdh1OCTdEqy3ydrhAadLQ5jzlAyp6f3Wnosrl7dJL
892HBU9qf7XkVHmVZ00Aq2+N92Okbayf6fNNVx99fSWGLckM0OEyjCSI3lF7agrUnS83jvMcQ98Q
H8QrZuHK5zDMs8YD+VWfo16fsT/hUjRyJIj/GN/bauB1aLl9XdCQdjLoq+wHbYcrmiLruI8Eplrq
SAZqGtETCUsU2d1hXW6ZNk2V9w2XZ2XNKXXYwGi1jibh8iLmRls52LMiHCTcmKfCm+zlMXk/WvAk
KxpvxNKR9hnN93C0qhWutrnpNihuxuxEHZ4YwfykovG/7XzkypOQdBJdH4+EG2RghY6CHzKozcJQ
lnpSt1EXtmrkvswmyA631T7aAyvZiWMF1eWIGzP9D463nB/kJRb0ZX3aJXXaWzfCQNytPvIuGTp0
OON0mY4dqr2POeCCb4vrAxI0hxjG9TkNCJM5DmTpekHCGwcFDsVAdARrsO8THM++CKPbJLsb+9tD
9H20h/rtU0vRYZxK8f9VKbgBno/dUV3kTVRupFl9kui9FpCHRk+ylvBlLX2kqMSw1A/elsx2sUF0
rd7YWNJsNi6Y/Db05lqmbjsBQX+SXHFsSCB5PMHzOaeDVp4B6+HN9GC7rTy8rwXbm0TjB1RMS7sV
5z0RrkBrYLYGXSY8e57wTXsR8NdeGmZ3O8R1xj41t1lYQmdHHwPR1urFSjN1PCLVnEiIYU83h5Uk
O1NMAwKsO8u9GJdvZv+cuZbHsYqJzXvsaNSTkKG5Zyuvi4Y+R1Jh04yxBTqj1tmUavLYMI791k56
AMKnV7JM5FuJlZgn8dudqoQcvMLdxsdvaKQG9uQmAzOykhCh3PiL+u+SBWzkvcHsXwUJZlONd79+
loSP5DNXzLdI7324c/mP25oXcCIaLcCDstWVJbQD4AF54JZ+ygG3cqCzU8UJRW1EgWyHyTsN4e1S
Whhq/dyZ8nqiY5kN36fvoeg3GdlAiC2TtsMxIWFrNA+y2eRRt37K2+0/TUxlH1tRnwGhiJEjYOne
dkYQAf9KUInu24iW4A2OrKOGzntmBWUhCz2FJiHj3Veu/Kqlems09mZyc+JfKybXcKIUWaw4DOoA
7QcMbSCbjboxKRHLYnZTDtcApLzAyA7SFt30sjddnFcsjDUvjSKFEQQPL8uqFHIlEK0u94BHKsGZ
wKwQSYq5NzWSRfxrJQXOz5L5XdFTKL/2ZRNQKUupZxvstXi86aY5mkMdptHZYYeYQE6WBk3UiGtT
m5HLOO1MTZr3v8sfraAoYqmgdvj9uUto7kFiuvRaSXEIgQCmK8Y6C71zyHIGC5Q5X7MttPOnYbnK
GbvDy2e6/FNmY/Y2LjVIr74b+VUzQd9VvVrwxfo4OKVFyaE28AAT4h5M6FuXF5vARt25xiEI7fxw
IePpF0lz09NB1622HiSK8j22gNnhLkw0EbbIgrGXmwEKf5szhkx333E+grslzDABdeBMnC7JzO/B
ugNxMe24LfT6g/Cu+Daa3tUlWHdWzeFRR0owTHaNIq2ARaHg7eFUqNASaab4XnrNq15kNazQPUhk
GD9cY7/2oJBBYil9pMVJXbE6t45kHezTjdV3SnxTUAPqCuJ98wWIiyDRJSkbosrJpQBf1PwL3rLy
bPWElpiifq0eoNlIFiJ29udRxgTod0vyqruz3j/OAvbjXba7bI/Ty00wqGHlrCCuI+o7ri4Zs6wV
/ahAkItkcjhiGEF6opsRsoCLf4Hgs8mYqGscZ0+SFvw9mx7ZEHaqi1+AU5bRPprjOYRZQsXJCtEy
SLg6zjmTTMwjHD9IohcAcSrvjSuKXwhZ1m2FwkN7WxRGAoUqUh1v7mMb/mTCiso0eqxtDJP3oFl9
Hzfi9EFRNOJzz9DzcSkzKuFxTVyylIi0/QTeHnVHv9UDJNwHqCrqsxMd1J3iOXVOyI2MOCW21HC5
nvVVDRSfjNJVAIVUKKkXCNaIa0jUMUMd8ytkrhWMjKFyZsIUe4AtCfDy9ldVCo2UHWK8SyYb6kMa
XSEl4f46OR8GLnYY0mvS7n7l7C8Cn7xZQA3Wke+xRPICKkxCAc3tRJnHxno9MVSsBGVnqDy/S1wd
yfQPEFrfMPBDo4Z5AZ6pZeMz3J2hbm5j2s4SL+UTcocRj3WX2JYvz90gymUbSGJetcNyRslomLxA
SjfTeKP+4AJUvTJa4+z9Kq2mDH2/6xtJVpJEIuiyu2Q4LachRED/HzQw/x97OfF2hu2sWx5U0SMg
M7BwyctZlgwqOrB/BIdGBUoZqjCyTXCbeWqUbtRMTr4uqVXLTWAaox5Ndx+a1Ad1GkkAuAgaprVa
XQCrmU34LZZtyn88jAnlUbivmCLgOSdsxZqxq9N9Fl2Mf+LzIuxEZF9BTgJz191WPlRt3vmdwBvn
MgCCeb061uuRENVztI8STZvdV6iTxCa0f0x0EZBy7IgPiVVL0VnQkB0gnVs2lsl4UkLjiw0NLzAF
sEA62kxlukSYEJ9VexGR1kCpUhQndeqyKF6Yb5ASTeV/nppiIMXf2l9XIFK9WjPUxk17NtnZi+SE
y6SOqM0VXeqsaNSs3xxYCFImD3ToG2O+HEos/a1fkrp9yOpFf5yHvoTfOUteX7Nx0dLXScTeACxd
INFHDZHx2r5uiE6Zc5RQ50oyIZQ1lMAcJ8jauQ9F9TwdyCAbX9RcKeBoiHRHL/z8B6KVEIQU4wNi
Unf3VM8EWU3oBZZBPKHmpjN2Fl6ex9E9bwzHMhI0xjOTJ5pJBJ2014cV8IrmnQpiuPEYsouLsImw
en29HA1D2TdihNBm/XSXxaXGHPh1jBvL1LaZ4mN9D9fCa04jDRTgAWcx5PYSEHBDd1+nCof9R2vA
Fao1wDr4n+eICHY1k7PH5RD/QCW5Ghcb0uAcJi8rfIkGUnUb/xk8FswAfkOJH8LBorivzAFoARFe
2pC+Ojke8azi7acp0rqx7jn7KUHhuqNYWvA4MHljMlmyDoet1HPg3bIAtsk3hIRhCTWnebdiXE/1
PKOwAsZMzRe+eXhhiWSZM/Kq+gKOohmPyXeL5OvyKsVZzwXbYsLXjjj/lBGo3MTwVZ1JfqnP6Wto
A6XFdcTIM84RjzYJJdduh1uY0cO39PKRBJSebK9jkYhGRtZPYuLRA8nK9J1UJqkAW3vuMILZxfj8
NOcl4jbJbs+uWkwN+VLYyWgeTfegZkauIS1BLc4ufUSf4WcJJCCIOc+6LA7KsNVzTBkTS1zQKHUk
D2aV/r+cpw+vcjJ71OmCgKH46J+BKI3wHSsS6OJHcTthRwZq/EUQWWjrNQTsPk3yH64qzYqXLKpo
yc7jRdYRYv3F126UhoakvTrjTe7OmNgCwZuOLmIuiiCPhj1Jec3aKvxbbFkmgLR8alG432rKTNTD
ieJlUv8K6iy0qvCpVsqwl759cIyjKWEkMnW256AHNzypfWxWg37I4MXuVqqR/R7855jwkZEiz90e
C+t86fo5hQpskGHy3Mx+rFiGxbup2362HAgD2zQSl98AiO0QfMt52qae4ga7SLHb2inr6CN8bAgc
BLZ439aeQolvWzz1p7a5IwJqCHr7mpZpSbevYTUW7N0o4PQYEeRd4kh54s7f22tdMM2sxRvzwwmV
lI8HsEJmUAKuCKTFDEJAnEsD25qtiCqPfmzWy48J+CpdW5DPIhR7lseP4iKm2V4HsZosPifVlLFE
dLbedD4hsUB/H4M6sog9aFQNyNJxo4fcENst7YrR1tEF7ToMDTAITUhFiAiOJc5ilX7LxXS4Ky4C
0WWEAuNWM/kADx/Q3LEHP4bNtH3Qh21JpD6Pk76hIaixqvsqr8+SAOFN/DHEd+Pf8BfdzYgBnXYk
MzjFaS6fPMj64O4okuBX0a958X2nyEu0rqkONTamYtcCxfnWSlaRSlrLl1eG9C27MwgfJ/L6y7C5
nbpooRm0hSNWYV5L3AJO2hloQBZX3P5KBIpnX57QSfDtiI8saXbvM0l3nacRpaf96VIIKZSUhCMm
wqO2niDDXdCMGve0wfNBtPFscXbnp1FBPrPx1c93VwD1Kbpo9/GB2Q+qtzxbMsW88Mv1MvHW3Bzg
wz+ZbG0HFcLgWussBEP1J1UZf6Tn7SFRnhgzAPwGzY26fiEVSUsWQtpoPcnixdUAdXbBfOAW273m
hLEYENqpIMTu2QAONVUS1Hm07/8ZpS8jUvuD1J9xi5FtL6y7RvE5obmfgYxwTT2LIfk1REZT/GIC
wTJc/GDPalBxPob3t2Q0WiQGNdHVhgt1YqvTE2oStnRn6xy43Pa4q764LlVem/HqmDvu2XxXAdXk
URTKF/mKgsDt8pmV+EXoXr1PVoCrS3gvyV2DAvtmXq6eKHhM7mc0nFSEXSSdDZIRMupNhL77Fenv
P7QlQMYhQsZo5iwtL4PpcvoECHNePO0Kg24JeVDe/nwWTOr0ScEJMGzLLxrLtTPUpCfdUxxByXh7
TDwib/ZS9NHZ+71lnoqiIxG0KAjCNt8u7JKlC+8lwLjN7KauJ13DtZuSe8cJjxs0IrzMSFUvK0P6
JW8eSa7h+GbdF3XNpWfx4JxGOB+GMvVTvyV5gFzF/Zr0nx/nsaGY8EbYbTjJz62FsB0gyKb8v+0d
7fRnNawEl2EA1QulEsosWJ2rjj10MtBo0ORELZH6PXWWjbzSeqRtBKrOTozHZZSn3vm2kd/9arCD
axeKVqJOFRRIU7wbZgYgPLC1ed8O0w6IBne+/EXhvmJJV9PwTG7H9RJc5cuFby7Zelecw8269daH
kO2PuFI8wpeEnN2uWjP0SQbQzF4OSxuEkPsO2fYD1E5jDMLEtIYICGpq61UjGfRgFBxeMzl5iEwM
oXoqcxW7YJBwHD6FkTaWsbIXadoppeck/1/oGf8Zm3/mxPU+hSqa7Csdl3ZxvN3caaH1tAXWynDX
77AKlYgE0bAszEIqpeLhwlTNo/l+b0VxnbCH9bYb2xFiKDvyq9vkxXBYqvUP8vB+LqgBo7ctrBG+
xeAaKL6P4NoqjHKzp682uJMj2HxR3HThiKmrRcJR2O6Iq8kVHRuSVh8IfCgtz/Yg6bB+qx6bDtnZ
yM4ZIR66d+WqzjIo/XWv1GhczWK4wAG9p2xlNiIAMIb01IigV71bqKVe7IXQUXqflGOyjTlus+3U
43qE/nYUQd2ZnxbeSrQOQmlZWlSvp0AEYbAAIgVIgz2VNJRsp7jcztBYq0FUabUOb6qoqRyBODyH
DaUINpffKta5SCSrBvD4vmYVLVE2LTIIszt2ld9vdNDWHVd8z73mnlretjxJiXGHH49/+ipgMQ+f
cn+CcY4xBcdr8ha6yrms+bcyL33WEshqnUJYMgzH3BpWP8Q2jbP+2URT+oivRc7AaxW/S5jeeHRJ
qGBfQ2BaJoKLWnRmuAX3jm7NVRf+GORHaq3mAVXz+XgyXsyMoFUXH4GwQAgzIbdv9gJvoJbaMFEN
SkTbPLr4TA4Rn9p/XFA3J6a2Ui0yOTsVrgsigjZVrkGhPjBPZvIpO+1/5N8HOfHXcGGRjCs2cY2e
6ueFHBCrEAD+NkjKkwXeFVTQPjcOABnN5XQqvSg/wthQVMu1g5/HaljoWMqtON730YF60U4cGnEO
9pIYzHHOatJLzDSSuHp36SiCzDrGEZDBVlfTD6lF2zQA/8et9V000eWKaQ5H/7MnGd+qJybBRvYl
jtyKdax5E4mG/B4QF3n5ERXIkwt4lzRkGHCWz8Wa3aIeSjsk/23J9ckWUDHdxBKvrVlpc9vWhcGC
U5tDJOxzzmC4ozZyBpxF2Q67c7e8JbJfsiGVE76Hz0b0X94fcbI4AT8JNAHt5urYlOI4ZKywPwSW
6okKaAz6f2cOKP5Tu20t26MLPYuIngQqhT1Xjxc4trhJGoAXWZDv2U4Kl1kJnbqoQLyT6qxZ5kTw
vlWtv4L6/JBiqIjgP08UTrVzcMIqjRo3vxhscxJO6tbJLImokYzCKhqnyNX7jnT8crCsfN455a5h
NCM2wdTJqKERrR6QG/wgJm5hIk6e+0MrjlApZJ0mkjDMbh1V2+ZNUz/tWxjRu6MefA1h3kZAVrBt
legg+YYsZfiDQt16EXG8Si3WR2+cSrz0RHRuksZ8ZtQW4Nq+FxzAP2x2eTb8hBq2gTY/AJ9KS7Yl
cArtJpO7vp/SRobx7wtf8PGO1D9uCuZtpsZ6jHmSQ5FZ6i1xXxcqsbbSMajqz68XfNrOu3pqlGwK
MAF7dbQ1gRUgOKY9VMpTq8++SigYoPjHJ6GL/Z8RHzxdmiX47CowyV/gZE3HchN9xBiaOju1GgcO
0RFBiM1bMfUqEstN4PrpHWPSqPif6b9Og8oHmm5qosLzwmq4J/ECirOay87QYqnN9Pm4bFjLD4/v
plEm9Gkcpmbrnpj8qrShk+bgS6jMDSsUHMehrhOFgS7unje8qShV9SzOlNiTpQcKnnNDiXaQJzQ1
bbP/6sB6WQZ7TRpjCU1FkrFhTy6rcyZcbfPoX07PUpcryvo4LBmP3RFE6DXVHrEP80rbFokm0lEh
TU/mUrzvMhwAaGh0yujwltE0QJthsKv9bwvpxcwq4UCSXcpqSaCbcj2GFGavja5yYQyTTV5YNw00
EkKBzGLZ0pdUUwwrQ6SOpjG8sczNjMUUaFvBsNb4AzxMN8JlyrFSKWHBVQzoj25RueOV6PYpP0p4
GESm9DiOwzetQdlimrlRxQUllVP7Ud0rRyUf3jcDlHakroJdmgNisr6Ps2WM/2H2rMH3NuUNKvSP
5RwKnYVAMyko3NpH1jvn94uC4mHGadiPYI8ngKozeOgYoK44cg1USTIJiuTW5s+SCFSa8LmunRia
i1oX7QMGrkd6X/yUFN8Chumru+ZTlUBGUP6vAbZGvGLtO0oPkK4tasvncbBivOQ2smXM3h7ly0bE
DIpyVpf8rTbL0u325l6ficngMklGl6wBJS/gh0W2QQ9khudrEdpuaDk0ZZOUc4eSxa2XebNefHBN
kcJnZzVhcR1oAOSOlMjr19PfzDdrdipNbTtT6nDS2iImzJaeO+D/BYU53BavM9Rv4VHWhVYcShpZ
L2kmCQUxG60vJ+28NyJPfn2kNUK4cZ1t+S23lHs0uBgd/pDC5SpGdqf2h00aiekZgWs+YL7tYFHh
Z3ArCJLhjeNReCGe33imkugdFMVu6sWf4nkNN/xCLM04yPQevHZQEfdkrRN8h0+F6AJRD3vjEFm9
NapWK4BFeAXx/cE6Wt9UxzSZLSQlrpymo4bESbHbcxj3UW4KZ97UskRKaNg9veaZ+3eEOuglVr46
IotSvClDPsVuw7L+TcRryDDu35q0LO0R8FL3GgMCdAN+Vo1RM36fzneZfT3K4iy9HTLDf6dMFYyf
jjuDe8zxLj/Ss0SSd+upauAfkpXMC2UxWXlZXo9qEOI3bbOiCAuEJKmvKqN3R+bvcehxsnwNSRmp
DPz2vTagAPSfBgX38IKl11OFpaiVvbA2BMAOcv6wFwEko6tFAenbKEzQ58jA+j98WGlT5Tg6gB91
20Z94r18gfH9pYzHUUFCadlg0snPgk9EAu3m2XsT7U/y0629o5YKjjqFtZ5T2WZP66AwJUwjX2P1
5FHOGva4lOQkGGQ1rLO7y6Dq98ISyiCkm+fs8+B/eyDIfLoip9VVJ1+8UPCeKGYaJbMN5c1dA+rB
ghCRCnPw71jIRy+GNy3Abs2yjx/On5GU+8oyRrEqGHfoQ9+xgcPBB/i686HsavdETqb9LQ1nThpj
1+j8H1l3/cjH7SCmay9lwcghcPXCTxjLoLY1J28JoQBtD71CDIakehHqGKIorjJFuRaFX1GNBk16
jpVqzlvBT8BxXlMFMJJmx0uaKGPKFpf6ViXPsVVDLbfNRUp498w5sb39XJHf2e5ofOg7xhb0/qX8
S3N03ptLbfRWd5FeHs2X99QpnvKADgU9gOzkAjRwa8GLEa7ahdl8sJO02mnisTEXP1X0rsl9b7y6
dwMREC4WE2lJg9zx8DTJZ7ow6ORu2xA1nV7kAGgHlmhdyqzJiTgFbNumg3q6v87TaSq+LUtOX+dU
itHaf13yOLHGYVLT+Utm1xpTXCOxq358q7BVpBdBp1AdiDuypZCPJPEKQ5uyWs7TKhHRwFi5aiwx
DGXOaohgrvDyVtI8rYf2T7kE5XQxeuY4a5RMHcbmhIITdpp0Rtfvr1/CbKYaPxfBZncgSVMquMoX
aSmA1NXZ5wGlBNQCwrnIJFmVSR2lqO6sBcFa8jri0OqClbzm7zb88Ip9xK7MbOGy+M9qgiJIwGeh
5THKWduPIduliydSqWlfMS6QP9gmAt6EmH+MJbzEPrcXPXeMgK3Qp6LCppuz4E+9TqrHxZfFV4Yz
42DsPXAI+D+Jc+gS5tb+z5Tl/MZyKwjFrTvQ3v1wrARD+ATv230EwaCAlSgzM/m3EoFe1pQ7zj8z
7XnxvT5u28yiRh22ElYWye3HpAvLnCer43QQPvGDXKvLBmufX/QY3yu5rho1rn9+oJcMolbJAcCS
FrhzSyA8zquyySflvfTqjno3kh48zKi8T+W9zYjdqlk/mp5+jtg8PlSEf8Oqtr+wklZaToBQgj1U
pwV+Vz7Cez4cLyhKpcsl0aE6Id7+q4nSdwfvbi5oKV3P6Q2HAygeuvgOcWwYzjicrppuO4ZEwfKz
gx4XjVJ6pFgDtgeG95ufctX3tJPGYPlqWTsJcaHjTHfXuuCZcp6mIRfz2ll0mFONoA2HugBxO1M/
r4j3yXjGraYfJgggUp8ZKquND9jjNCIy3Hod611HbKyh5qjpuRMdOPDaZtlrTCCaRWeZs41KRltW
5/EVw5mtsOxoXKG/Yo3XsnKHCOHdoBhyBS9y1hV6AJjrWOsjsE2egVfIbds4Ttcd2Nw+SL8Kgclq
6uAax3G0Y0OXAC7to5vjQqpNO6jF6G5Xc6R3kRzk7EnVqus6yN+Zouq7gwzbOGltFtQihpvXD9ho
oZNU/ppWjQyEKZrLW7PCiBoUmXNhEB3OZ1Xtl7GhBG+6+g8ewnPIhYmn9uryF9Flzss7Tb2X2CNw
0mesag9vSbASGp82dKj0N3DYM34aJhQ+9z2chusRSxvGLVcakqvB7npBnelC1k/3g5XMac4gXRZZ
hTtjQeOLLv4Qxa0m1M+vD+b3xHl3++kxGjAP0Zu4fbgEfkE/bIRkUatsJCA4sGznX6DCz/AkxBsi
uy+0RhTeb+zGLg4/igUwTJ98H5xAsr1pbL77zfQNlKKFBulD5VVi7FTakc+CUy/wr3LSZuMQUQ3X
ARCd8fvTRHjEYieSPO4N59VsntdvnBaTpQU8Zp92X4V3a1K8CzGBtQXqpRnJKo3KDKgpzz4PL3XQ
gyEL5NaxSzbRfYTa+rRwqiqHHbfFeUAhZrpyuGwK+Ays3fnXF+4EvoagGIlgyeftH/2UeHAKY1WE
M1raUp7sFn/sTnp28a147MR/dFSiSx5CRaOHyPpgH9qKtgctUvnRRX1krbI+lH8d49Fum6c9Rx3J
99icdPyIWivsQuKMPV7VrI1e/QLWGGB2MzCjmxvW6PWlqRwh68lgB9pTeouyAHmpOC5kpomqlLZk
5sdKQJ1zhayjD+LiVt7lCd9fasx309xKjPFtox7HhDN9Qu7nZw9AwUAEtLV0+xPydfdjrGx59ocY
dk3gE6zqOR3Oo2KeExYGFq/VyNJ1CXTAwoyY1DEriCtBzUgk+3L+8xG0s9Ra9rrMbsi/YnCrHvTU
5PpuWdtjazUwJg5K9aa9b2QfJlVT7hMFa9nTpYEhXeSg02sXFtxnSDKGEfB3CWfERooX3M3Imaz5
xWa9Y6AVjssh5FZIlBoOtnzx7vVTOX148Q7Uh8l2HV9dRikWHbpQu1lB3A5b+7cr4BKTFefOztDp
L/i5bkZ9mDhBCOUHGRhCmPbJnSLsQc3CYI9Icz7W4NBK2y+scf2t/p7Ge4mLCUegYTEyXN9NvNN0
ODfx2Qzh5MTTbQZPQsqHGdxlb+fE13A4j1VI02j0eHm6fErNCk2qQhxv1V/DRqUACIIhKtND5P7y
daPy6X2Y8qo75KEJDe/uCDj3PMT/ckM286GxyQIZSTXiCwvwdxf3nbX5SOaoJSUip2t6QZni3RO6
QYnrq0NJlCqW5Vj9wWvK0oAzU3G7jSfMBWHGp15pLq2Dt2Yk3vcjB/CtilRh17zjLb3ebSSCE8kN
PVpZRGXdSO2Hr1zz84qbmYuLR70LZo3b2gn2GUnm14ZctsDvHyjkgAs5g1oNZtymfzhsxXU0uqi8
fMEL3mdOVZEGS+jIQ6x6OtMzT3RtSP4UgI67g02TfT9Am4zibCudUChTGdXaZoQJk9RL+1yH2W9B
TPng56oAALGjuOn9hqWROxlIqurwpw3m7vtZSLAlyawkLNq28toPTcSTgfXjW1wVl3skDSwnLZxc
YjJHHSeIvYJ5Et7QNLbe5ZxCjOeYbCJnLcTb3qrO/eMCrF1mGRoka+nbaIRFUFLlyDzoYV/6TnFZ
8w+r4bq8JMGNRFB+Bg8+NIO19kOfS7GCjYzgSReN0uLTJPQcoyQsnL1TW7q9XiGGWn+NNdfhIWb0
D9rh6ghL4kQTOP7Lt2yxaW8EOLxTBzgwUVjko2RlX0GoOJDpQ6E+YyQutaMSeLdHGPFMOwwNUw1b
cVw4YysocceKQcnrG2D5iYWgAa5gmNM0TduI8rENfXo3dQNlWaeAk9lxWWGagv76eJZHYFlJYOzV
vLUl0+KyAhgXi7sV7Qd2Z5ooQoU22ne1ezUppb2AHHDbTE+m/oKxIQ7rUgdEnwnu0VI2PObIXD7j
AySfcXqWcVqEBVCPIc6mfoIUfDtxEK6w22Jo8GBv4gj7mTN31+o++PWacjgNMEoC0hEI6D7TC9Xv
4oXu4MsLXopZbzh+RxbVBv26Kkh+GWik0JZS+YwSzT9uGBdcvSHaTjpcqgflIPt9cXBYs2VdEHyr
k323WnGMzLssVndDnLi++cRM/L+ntzvNkv3KcSVnBzRHgWE135abY/wogr2VCZR2XRRZDCQtw/vK
rp4Fkc8iJJnlFthEaCqjuJJLWea4TDJRJ2IrvIvtpZNeTagmcPZC7F+iXWs/vLLiuozrtQIQpgNj
m1rPymTB5o5Fmdmxdly6PZC+KoS/iBe2nxwYoEu7C5Du6it4TDkkiv5m0VDgbSB4P+VuKSxVuDlg
9z+d+K86mrEH47N7x0LcpVOXMY5UY6bk1FG951fRP/l/ZSgaOeGUnCuoJnykiyylMR4Vp0UkGDu3
CSC8BzzADqsRxTE8BgfGPy432cuIwk6enX2PbAGy8QEdzJZcxPq0SbSYrbfE2hefGX9bcyJN2GdB
SBODQsKbM9q9it+cuxFsn212XyL1RrnYqrKn7bu4EBInGDNntspAezrealZsjs6YqO4ANtL/HegC
g03ClT0M3nkwZNi800LGybdVEsKreSKyLEdjAdgRqNtv+reslGzFW2J77nAs3vBaT3JpJsdH3VGv
cvnI1NvKLkCtXtex8z4lUqd0KhxtzYZm52z05l+ainfFV75VC0/ar/XApyZQOKbR7kmHY0HBPE9p
xbUzil9VxGALF4CCxHtCplf3MwSPF6qG9OphhnmBGPdvKjazgLfwA+QkjUS2eOMHmcMoCKfYhdRx
R31hL2eu8FORgo3R5+1Fis3Jt+tvJX+jQlXxyiatC8gdXYcRdZsMnIklTsUn+bzzKOGW8U2DX8JA
5d71TGPkCffrfWTjwKcVEqlzea7OfhithedHuMWFZyd+QUNr4+1u2vUUAEqz3mBZ/3rP3MfIG8av
OADSxbV4rq/cCmD8QlEiaz63RJgM0ohfgA3iM06Jnbc0Yytn5nVwTYOYuyo3UK1S2fzeOOe4L0vt
86pauI8F5GI8jMvJFgpedPDIFgrCZcNf5Qfq0f6r7f9PczzCTtfVm/0hZUejzDhseNv75O3z0MLw
uIcxImcivpKZrgCscx663FQ2JxtNNelPnj6nLJaFrH40/UTI6GnSyHNIo9BfnL5H/9FK3AFeZWvj
RWMOOh7dNBmLNRJWIyk1BHCiXK02wPEc1feJNCObTriq1+8PiSukwAbMbXXdm00dfMWEFG1jJhdr
9zTyyjpWfP1yBTXwcMT/A9yzK+obZ7ZqCYP2vYpKW1/BIPMb4ffixVx3/8c5iWf4Q0To6YUMLBd3
Ty5cRiApc+qjh66RCpf/T4+gUeQnHYhRsrDm1jboEQ7hIctZtuFI0lsNGPrQ9fXSmrzNhi3Co/Tt
A5OpZvqBKWtWZx0PTgo7rSdZ2Y/lc6uybBSHFCcLr+bwqcadX5CxjCV6c38FwwFcqA+chT4mmwpz
LiVgiiXR8rUlfCzrG+W0r+yDViBNzA+OYxskP5zpKYDqIxQPfY6lDXLaWtS6pRtTNkfMp+ayRnM0
8BybeeGENsoMzM2zmg5TYX/YXWyhWCR/phaE28ZlpeESoQzLCaZ/VbNGjPmA6vuTjYKPYfiLyvMP
t22uyMRPorm5p79b0DUbkpzibqs3K0b4EOAz2eUv8lPwHKJ07F7nvBFvjnZH/StNo9TN/LwISWGG
cz92+L4AdM0usYmFVk9waV4jK/prAfB1D0C3qQM1160g2NcAME5PuBpw4nnsVa+jbZ1TDXT+elsq
FlvfM/VwPayzV+/WizqtaftdSGSdg2vd69dYK10NF6hrKUKBHF7iP+tXNfMQL3P51V9yrDNXQJ0L
vkKdF6EC+Hj37Cl/qUMNVZBePJA0+fC0Ih3xPReieHJBRqhLrwruNnexjts0FPw6oqXOTo0iGv66
ejqskPARq8W4t3x4BtLOSFVyzvPPSDCSvwiWq5MmHkoEXhfmyrvpTCxqJMOZMrmjpeV6cTLJXOGE
w0h+8lY9M/3U8AP0PYMG55jz0HJUnt3e47kyz6hSEm2ADsQ4SNFpmunw6RROzIl/NA8/QJRLin6U
e03X7ODFTfc2BY1P8kzjttVR0hazgREcbnceoMJgdKsYdGtE0xFH21w1Qxv76R+oFX4cXcN2NnOY
urQgII8d+dhCsgLGTaHXLrmEExx3LVecjjxDQzeVJurSGiQLmtfn4jXaS3vYg218BBeADom7ztLI
OPcswiYiRtsCQSJQykyTnyAHToMfO/sfvI8JAvxqS4y/34TI77r1gd/s/u7X8kljmR3qeXmr5SvV
qWNmfnhUnKCPDrES/YbwcerMyxyRvg7w4e0aMyYXsSzXRtwrYfghrbehRkFt6Geawj5VwXsME8a4
m6IGT6gIyqX7Sc5tSgAgD8BKemMMZGTPJZjdVnS+QYQZiPFjP3C9gD2ei2w62BV1Gf8YjX6G+Pzz
CjwaZfODbFzwGAnlLPh4ZViekEfddv27c57/t0vampBn9+Rb5Ex+4VULcWPi2rUR1hQPSt2bqn0B
7TtM5PV4qcKT0cI+lWunQ1tut3ML5BFgtniCB3Jc5WMhHCeCA7T3NGnw9XCHNjS5rhIfDH074Dmi
mskBUwP1YUFv4QUVihubGbb19Fj3huPhej3ieI57j4IgT7L5jOaSVVYpfvJxGw4gXU1J1/WEEtAL
EUQoZLoLp9vW3UbHafOPsLVzVgcONbET1vKsoe+RIhCZjvKmVSf+j2BmtVbvRqYoF9QwbWXoIxHH
CPGeyPYv7Ea5WH0P7Zrl4Yn5W6RYVlo1WKKB1yc4Y4ZTu5jvmg33uUAxpqp4xqEu1chQSC4An9P5
eVqv8D+x4ZQ94/MsVOXpN/6zoCuA/8+3orL0MIHr/h4RKPh2ESZLYSO/dHGnwarf7UCa0sTTRY8A
Z74MFDHssyYY6diMS0lUJFf2xI8XGyiirNbMkM7mmpM/AK3TnK7uzv+h35CbpYVCriuo9FU0e/YJ
WSmOTbpq+gg1t9i+aMRtvlgSwk+VW2PwNNQxEH4KpQQD1pAuk9O6dQsBWzEJVpxXE1gMki1FHt0P
kB0+RtzAJZ5gA/2PIkLb2p4h5teuRWsbQ4BqjySyrIFN6vsY3Xqjir9C0DfXdabxLR/kJ1D9ei3g
4JvzCjwb5VOeE17DbsQQ9O7+tLecf/scsfqsGXPXXH2MdtWdnQVsz2puBt8M7f8h4Q9oRxDeT0x3
6/dUvHSYyT5EKWLz58yNrcE5GVR/BqE1SPDxUQ30QKDvVg278KdxibTNIpmZykoNvCz188fHP6Wo
/5OseLrPHMMm71TuHkrufC2Kaea7dvWgu9GT6lm3Zc88UFY3CX+PWzg/AXSgdDFox3CmGJNu25Nw
a8SP8TkZOVE8lz7e9odNLzyoenVJKwC9PPpxb8lMQyKMu4MjjS54bedf5ztdny+V9j/jLC1Ijqfd
xuKnkXsga+TwBf3rmQ0FFdBdpjJDPfCJuoWNo13yilkDhElG2X7q4+elDqq3f3rNwKYVN9rtHPHR
tqPITT8a/RBf51Ml/2KK5eRfRZvztafRmKluF0aF25VG0hR4Uub57vOh7Gb1k6AOVu00VVuRU+w8
Kqr+QqyzSSdh2V49hpFzm0/HM36/vBg0EnNvhkgfoJhJh4bD7M7/SbfSOAEm+7apjAwaUl4liswb
cNzbDeO2zyqSQZ1H2GeCAjBLLW7O8Bd3VVJS3f+mo6+UuBZUNfGmp3NmYbbumrVxPvH5xej98fRB
c6TEajjZ+aXrK9t1f6UJLDgp/0AfGqbGzn6+cR1xq2ZmKoq8SnwWdB3hdxZphYr2L5iKHVpiGueB
PXOE6waIGeekNae4fOZkOxZ37NzGBz4a6GPRcgF5LduxOsgVoz/k6kiaJn27FZkkdxuoKrGD1a1F
oG7YYiyhL3an6Bge/rIpSzqB82lPOAdXpi8iUuwJw3So8hmGui+OFAXpMhgzGB4erVSR2BrwIcDg
NB+k5COVE/zKfeADaKPB05sazbyZf4JssKfOT62b04fTFLVZSjeMJWMYNxpawsvwwHKQia7pGD01
hvhd8qNZRo0Akgwehtg2kZkzT94jpbwcxZilrpOUAiIXmVYXclt8+KUNwVwKOshlJCGUZoG9OXWF
7qMmZeDEQElX1vcdYrQFPbaw2dycmJtGrm786MSFp5UBhzuSybaCPw/ZqAXPLGG+recyYPWEfaVc
nG2L9lqSsjEDQ2tQqNAT/Lf9qG8d4Te3dssDRwi6fRH+94HNSqrkCxuHDQObxQZV+Uayq6hxfzEG
Psk3EnqxU1Hw5MdCCsYR4uEZFgKfbWmSuX3s2lpCSrhZ9597c3qix9WwwDy5cOOrV/GLJ9uEsI/+
+iYoZGrNtEVoLcVwy4jfK0Z1Ew9fP6FFtNH5B1OAw9jJmSQmw6/MULof0ptb2lZ8cCILN0Ulw4FR
XO/sWy+gzp5L+b+TS3ci8wHBA8M1+Ia9G+Ejp/RN+ul8zKhWe4ygq6YxdB2LZ1cdfGegPWCIIxVT
kWVAds2FCNg0oCaGBsDjUnvb12U96rMttvi8bF7PLIFxm4RCXZ+q9jAfzZsHbvOq/NLHlJiMFFrn
gugVmPgAK4UNio4jEKg9BYT5eWKa320EXw5lEJa5SKtqr7uo//e7cFlCUbGC0e34RrVk7Cl1sYKz
kiHtTQp6nnqDOSKHMBvKHn5hbGRoKPRp5R534VJqiyZvh/ATcxJ6K3pVO7/TKopoyLzAzgpH5k7H
4d/rorpkAS++e4P5n442+GV6MHzv4ekxapWEXzjDz6lOrsZXSBjPAY0gbb60LuSEw/zBjjzCW6o/
6mpOnOi49mNDEKDvg9kWpOqeS1rsJA8YVrFTuzcFltjvZ2WeedV2KfDklntwwpH/YBRrU6ULBzyp
ScJgIXZaaLA+dUp+Da81R8fZbL3XJK1Ap99a+uudjxP6vj6GRW65FYNCzSbTpj0Ox99G5OASLHGF
jD+QRDBL40cOb8H/WZHodp4JJhmpnkRyM8bADjsLHJGVZbd6GH4DgxNSYOsxuu7WsXwrDpxD2Bf5
AuMyq6bla/iaRwU1ESiWhz7umsf4ypBuHHPs7y3oDaU6X8jWlaL4M0of/R3PefK/SOYwUZxrZLTi
FxSaWgppsGG1UGLj1Y8NZOaRGMzXoR6VvDzqv68qNgdDlFNK4GQlNbA9M645g2L1c7nLJ+MRSZLM
WtRTAiWYPbO20R7VhLFfgDH/YV3K1XI1lF6wpWG5w4duI43CxeefRW2cXAEqxcFAU4TH1r+OpLTd
TWt9qjox/vZTzGQqd6hS+3j4DJCD0DJ2ddLlx5N1BXFxPUMD0lGTrmzIYfZwhPmOJjvU2oYlqYvd
CwHO+AA7k4+5fe2MU2PVXFjQgirnb4ctStuJSUDELDMAoqV1qHH7HihdLDA1xaSWaw0IEBpu67Bd
+VEEr7bhizJ1HCUE5a2UQhs74D5dzvpF4cVKp7k4z9X1wJgPlGqmBtuZpm+38XFP7BDzJAWkQ1Z3
hFi0z2DcGONbhIYm1OLwF2maMA/gOIreJgczf3LnppBD9sCsnZrvNH+Jhp5fUv8GyZrFVSjzLsu0
x2yXNPQYHvdcrydoQ24zUebn6oWvNeMhjfbD++Wb2x1K/wWBdUiRoEg0flxGN7FNesPb89mi24yV
ZvWZz8wG8v+JWpTzFPHtqwgTd0WhXGJGVpVdVRhTCMwZ7JWeL+0rVeFKmRIa/WOAzqfGp6ojyjCS
w/wXhujufp5Kc11v0L1MuczXa4rWWInC98KcTnDlkRolnUg69h9vfh3ZaCX80k+3kYWxHOzJKAho
0VwZzcINTFSKt9N0tLwRX62rU/VCC0Jn1fgqSlvZB5F7jrUI9l6+0QjWGHYhiDZuSDy/VXLclDoD
htK1ph+v82d7pXFX6eTEm7KPPozRZno/4NITMU2zOWK/sxb//QXpgZYXp51b+7k/W4Ia1YKOxp+8
pUtQpvF//bGC2nI8QcEq/SNmgbkbs1PsjqJBFP0N67DIBTw7PAESYIDw4Uu3s7xWl9+XcPNxUp3L
Hk78avyhxJ3mm9Wqtorw3Y7jiK8+6y14QL+BoVHiACzerGPNkfCqScF36ptFQL+ZW5pzNF1dhIVe
q940gjWawK2sLcDBzAPsnrDaIoFu3eHem6XZKKQRVJqCK+sAfVotJILQCHwroqd2HziVw2LlOZUK
lTv5mKx9IoTxeKuM+LI9UMAVi7R6w1KarU1ZVEvlcRThN9HK58TYhJJB2T+frRkTriesQw5O7XWR
wS2OIK3ni4rd0ET7MH7uTcZXd3NBmQ6HOxbNv49OwcIux/WJxkratH8g2mn53meicE/y5xBOTHZU
6/csyaznfMVn9VqhZqGlbkAiNLp6sC0m4Mub5iqqqbcfykuPUcKR0UZc3N738VwyGGD/ZNK+wjiI
YjWfSfqXCWHOU5NcYwicbsqzdx7tOmFOZdwLnqQeHMU77vFQ9K+GzHuIbYGqcImc6eDA+V/tvAJn
tsq6TzU7AAP2cJN78U15n0dqvkBJyB5hGBpeASbXg1gf2rn1rNSnW0LfMjxjwzOOiqkpPhMWxgcq
+QtnZbbFFTA7AmVviX0eibtaIR3d81XgK6RzDQu7/u++vcve60LDmbMnkr9NSFs9l5AM9XYStHbS
YCwamOP7IdMcKm/GkeCGYCikdTSW5z1fUK/7bydP2LOVOulOOHpN09lFuHyWq7wXEdemUdjPJ9yA
TcrlxFJgq1xUDEJynBL0DzuKKDD4DWbPZfAxOeIZn7zY1pt1zvpAPa0gaR7xwFtAQVvb3QgZMv2i
rPQ9h+wP8pOPetazq19Jh9oHF92qfSgzBL2qXL4vNw/uMpqZ6wTfRb3aFq7nTTAk+OiDWUFkjQui
PYveH0WDszY5DmABQPDzGyBWjOhvR6b8jGtBDWfelcmuf9W66RHh85xv1QCNQm0jZ11VpNt6xSCZ
17KgkEDyfVSNIxnHklfMHpPNCvbdSl8+XSWyoGjBYo4ygu0KWQycVbexV+me1oL77oaP12JtZgGv
PuSbpAesjEFxYs2J1nm39oO2qKt3Tn5owZ1p8mg8KHsadgcXxqPn7NxavE2HoKUxzTbVzgHSSdNH
oWsZ0F0ASFh+YZs74B9URvjh1zGPKAtTPz9Wm6/RpyN62RW7RhHnYSOqw8YocDIKTAdu5OxmZU4P
Jb2JRQsxKSot1xHUBGzK1DPibsW80XS78mXc+GzqnqGX0FpMOnw/FNi9eMREyliqBnYdhqj1XfNB
xj0RYZDhIZzkg25si9cpNNJ8oLLLq5pgIeEmyrhH3jNIMgz82cxNft7qGDNyJx6JFJZkDePui7B+
gVCZrtwkvy8scGY+dj0vP4g7qbYTmHFjN91cuE0dhHScZ5fOmkSCsLTRteo/uGDa6CVHpCcrNGMT
eY+7tV4QTfkynzsjxFLM6o9K43MX/RoAXBcpObljy1zClYV+WDWEfN1CTCR79ORAWsLIxqdKu17W
S/5+h8d6vl3YN7KO23qlpOv+uErfcUFfkVOul3dg6gAF/9HpPJMoRVhSceYTo6poUineyV18xZni
wcCYn8QFbD6ZgKEc70MJLgscl13OHz8FNPZRKft/ZjgnS0RZkI4NBw12w4yMTyhrx4ult7JQ3Kd/
95I+TCw4odoMVHcKq4hc+3B3wwQfa8tqvYLB/BIJw3xS2rArrnkUjBP9fEdxwVcyaUOLGscvscC3
U6J9+gfpa6CjNDA2vqAwfIKtT9zsT9Lri8jPBj/y9sakUfZ9o+PmxZ5nvPmRjzCErTCELCsTWaKO
bmaxXDEJNYQxnhpmiLh0xBauLNkLpOc0UBySlxrpKwfNR0paLnkh7FTDEvMBJS0fLr6ykUSAaF25
mFcsDt/VwKwWmgrR+/S/BBCFKoCe3M9yOl0Qv4df3uUC/A7iDms/Cj3Cr9IUByd+fBbQ59VT0Eus
4fhaiqnzeGDZx1FghW0DpgtvgPA1XB1XJOoeEDmc9c6NySr26I3Rt/6YTdnfAJJiT/LHfgo555J4
R79o7htf5CD2UayMrYLAO10FW6oc/V4SiFIc6EEpbjgzgGLVF2PYNYHd8fUzDCY6xpdqQuzjruar
trOzFAkDqNJy67NtDdWbDU/Ey2Nro8W/fyphIKE2arrzTEvTAzaytZF1wzfSYih9sb3EygEupf//
N7Vl5604ZYUEVX3/W8LgQtJyM9ddVdugMUF7NfjwDGFgUaCXywJilFJQzrURLoHPItTOJlnrx8Js
TuHE0zWxJrADo0bHYNy6dXIZhUiBhWBRwojuX/yaNq7JPq4DB45xRAT+u4IFY41Fcs6f6HyK/jyI
oCXam3dhYEd3ONPQlVdf2imEnFH/9KQWXgD7cyN/TyMtOmeXrLuN7IROX+7gxvcVgAUSxZ5HTmf0
8YnW3416+zt1b2m8E3N7oPqY1+2tkIw/TaTU4wNmAAWKGGy2crYbWTMS4ZJu1iIeeoJcdedvyoB5
AtIWeXO1kd7JeJXitXGCzhe2vVboZzhQy5DkLSbDgQfHnOzS0tA4LnADDsr/rvxjY2bNaY7rwBIE
4g1BEh1tCw8Ak9CF9doYGxjp21kNTZHqu6GkpINMgqvvnePcckOX9oNqau/XMAEArs5xftlaGonl
m8zus6vgKw/gMxFcFYaniSLgEXkhywASuMoSzUWgpTPGT38sPc2wCJ7R3gDUVlJW7afF1lrbu8PE
/z3qQGH/CCNUarP1gLOgXfkXOoqLVydZyRooocK2J0CFll6STclMNsTx9+3gHDLoT41YADw1HWB9
Y7sVjNEN4XzJWhlPkjREhZcufAiR5n3XKSvcdjOJaE8apDnOQP3EkvcOyCIHmYqzIMLcWeLzmPw0
pFQE6wZXJYnF62raW2ASLnTOm+rHymsSJ+gCbuIHSJ6tAPjBD4VUUS0tTwf33cS6W81mPPzfx35J
sR6a1ftQ2CBFPUPRcmq+qMiLPlPzK60Gdo5J+8quybIsyN4hzGyTmdUiDBctQhBJTnbeSacr6sqr
YWg50MaKbAFdoMP3KkfFXcf8HDV+ITeekxuk8o0PwKqgOYKQl6Dm7+5uxLDs5rsk1XitY70M7OAm
rFaGTsTpPR7A1lLfAQUC/9oDCW9OVgZsKO0Ph+Jhcn8rmnXo5DYagc2J95ZpupqIZyd/49sUQrqr
wMBwNThgIPOhXayC08dzJEHGoDLxiwV0sBmOA2fz3x0HoLaJJJnrGxrrQXf2CJqPRp64gas3prjr
dGaeDNPn3Y8RGYRj0f8J9RR4IeOhFlxtMvMJV38EeB/nxgC8gc7gLKpqQOB4zeuBDABeKwqgtrQh
Fab+L6rVhBJWAybvmuAQvDRXrp38WinNPcyeAEYCCO5CZhu/nBus74BInucdLV4+BbDxQTBMHe0l
J4aZyS9WMujeP3L9teKjWX9g72+z5VArJR112E8NcOqgrKo1yuK871mt84FJtiuTcfqxmIfjdWtg
j0ia2LG0OgKPR4U/p3Xhesc2kvqmNachrTg9U70AhbeazSYnyH+qX73zwYc2z1Sxc5TxAQgSeZ69
A0kZQ3UA5DKPyhxZuu3y8coJi5D0GHVQDmAcdfM9KgQjfh3y5zbYDm3VddTlNbKtkRd7uQtgKLBJ
kLQKGaC3DPRNU0Oa0YJv2UELIUDxiVwqi9bjAZI5HNXoeX7kfmfvvMxXnnknj+//5v4IVOlXnnMA
Zb4GQqPJUA3NNbns5hBQPCfyp8Ow30CTfmjbb0tdlB0Q3BrHgO3o09repUDZcEGhT5ijfclpbfDc
L/0IwWjeFcFWvfddhWjE+atdfJ2hKUT68rrBMGC/rOY+XNQR/5pEplkAuXcvKHOL4I5sLsy1NDKZ
2felkojpg7qvoH4jwTHsGN07a3/58HcTj8/mU1YXl/djrILOipSWO3cyS0rlfruWXRbNPPqoADtC
jnJtUP/X64IpsUACad1WsudCF6cHpSdgDsl6BgDej9bm71cfvqjtGOOynBHjXiDDT+cayyOjNOtB
zBCzcmHuaDVZuR1h9RD6/6RA7jtqhJlzUnV1aZ5t3PEf2w1e6JZJ2uKvXoNF80Ror3ycvD6Pmsck
Vna4oYx9LgJZXlA1XMWDwg+ixwLPpRhaMP4Ekuq6tx2wNOq/VakFMrkc3RFA1L9fu/GyFJ9o8qXH
YufqRBACOMuwoavYcMCa5yY7queA7iLWQj2+QCXWeja26M54lHjE7AN3p6Liqpgs+WUqGVlXMbtf
l459Quch51PyRznS1m/63XFUFhgE2/xcDSc82LMAx6zxArQYucUSYZJ5tUY21znmCyNuFFv+G2Ai
nYpR23OgtNvN+iv+kJmQwoVq7NDAivK7nqmjfANGGBdcVVqGuD2xx1bvl6C7cwRm/9lvFAVvbp+5
HqGUvgkYQ8BefW6X6+GnK9z3JG3V7v8jiUog4Mwp6wYrim+1LfnFnr7MlR0YDjPazKYKNXRcONu2
dXhx577dbvn8FYg+uFhT8NZudSNkY03tQG74fRRCSSYOVfVgo7ehOmyCIdnNj33jLSHcm1SGSBPd
K5+rGHrGY//xDKHqrP/vtcxzQ5dJbGTfgbqyFBVzu3L0TLmn+EhHVCMK5F0jFyRcZ9/6U6SZkeoC
MFH4boyZtpBh6WOrj4Tb+ZQ5YB8ThQkBT7MQtP093DD+JjMNXyIvTw59ClztwMocIAxV9VbNxNCG
KmvjOTuUklJgUyLnzTK2cEvuazgXZ3mZnIRLQ/12ao8C2nzTmxUoulN1FtKmBL41Io2/GEn2JI47
sFQhqhXENJFt15VjaEBgsDBhvARrZMIB1fDEiOZdS+wux2cYNRjxpn2d3pHercG602EXRAeZZy6D
mmQmfld5Sjed+nao83k5kf2DWmbpRahwW6MkcPnQSplO7Z6Ng5TMOkmYPkqHXPcYZKWIMS/sGx8f
3KhOX7mcRGd/9v00dgE5VCliH1kWp56oYCwVmbW0W06pBDeD6QAVaSI279rVZj5WURlovW5OiSyz
/2nk96O6RT8DW1Zlt6j4AkpDajk3B/kzz72BzsUT4q5p2Haz8O8/bUXp57ouQ2jf3LAaJDRVVyJZ
4jnQKh6SmY1nSXZj6E0SsUnZRd8cqsvOV6VQ1ItKmfJps80gMpxT6Dt9Q2LqWMkD4AkzJj1/f/N5
Sm3XmSYH7LL9d1PzvgQ0OvkFBkblBFYY1FyVr+RC2bf+7nJKs3YkyV8nH0Xxf/P5AixMF6SEWdDf
oOwNvjcqalHqD/w3zYAR+8LS+BhuxggdiTZpGTwN8o24fEuXmS+Ln5Zun1xISOjNGesBGwUsaf/X
qnt2mdIWXky8zpFviAa/5l2PZxS5llucPVNTdX9M6MBcQnb+KBKeYHDKssClFrU9zRKX7u62o4Lp
X0JEoiNZsJwpbUV5ow6n+5unT57W6CHjuhEqPPeb7E3brWHJ/SXTH4DJLpm7kj49rxBhGxgzsHbr
s2ISnZPZ935aXH42AzuQN7F53e7KzzaaP8oEHGBybQGmL0amfPSTBqAh33DRHui9Z3iqA+g2Xp/M
TJasvLx0kVvEHklk4eJe3QQkWyYBarE7LJTqpWuL2DBQKMuyM44fXj4EHL3lL5Lt3cBU9czlEgYP
xJRPVFbLTWj2m/UHWZa4AEOMyEH4Hktii0hNrtS/2UKjTFfqlw4b+euMjpxnktLtPGvaewQo5KzF
1OqX5SjOYpfsBjSzB+jwfB0my3Jhf33QYDRzkS5qoZ8yILvRvLfo1uC7md2nwdvMXwZ8DI940Smx
yIq7fzoF/9jhqrXPPxltElrqckpGsKos0yv1C99xTy2oj6neTIILgC15y2IXZgh9j7gz+VQH45sb
YWoB9CSP7VKHLSjaRJ06uSim6PIEkColUDFjzpfTCGzpXU3X/R0BBX77YhYKlpoFuG6E+jn/4JkS
bVMfV5CuS9o5Ds1x+8UaY8h/yGi1JYfu2bwBhS3W+fBd/+3lMu8KhTGaVBk9aM5dbFJzvdLibTKI
MUnO2ZpvJogBmkH1FfHuKbBpy8xK3N97Xtjx7MyvE3cJBwlQuZiWiR4BuKyDT6nmcWd6qMm4iij4
dDMT6Ib9tpG1e5wIPJJVPl0tn3XOoNWevzvZV2DOId2ul14HNc4fC+kRXpi9VpdZPSaqLSjYiySl
/0IRytmDRiSyInq77yNmdpIn03TIoYnVxdQgOs50cJEaad1WQjGv67EOQKUqcdxrRg50O+BcdlQp
GcHRxtJV+olDQmnOksBE2Qm674WjA4CNY0z7mczE9JwLNDi0j6xq82BTyFvU9f4QgNSJ+MWtQyn7
Low10osAo5mJfByJhiUMC4Qj2XfYJdBanY5e0/Pdwnb3FQ5EkqrBUWnjcQTSA8Isoaispq+A5P70
9Zo9HFKPkhIKuxll7ZG0OPNMqDvOmno6w/gVz6FHLFYQVzNzs+rwWn9Iz/4hswmCEEYxB+7lwHgC
8nzv/aUsCeexeq1OewJP9DVCWajXdaaVPZ8g98TJ8FygdZfJgmd+vmQTDfUsP1Rjv2L4FjkuIlnY
UORq69E6LGC6HAGfsW6BemQJh3DCq4Worwu3Y22cUgK+pwTTz/jaOHayTcK+42KFqGaasfWR7M0D
HvLHZiNGJTShJ6mkXoUG61JRbRnVGy29TEfcD+FBhxdmLF8NBx+NntHcbm3grpqbkWqk4xflhNLZ
Lf57I2bqZVKJJXLVsUDDPoa8HlOGhMkJ0cNRi8lR4Q3JeRRt5ef4u7LEWuwyfDS0bYyKuIMzR/+G
gJbsZghn9/SWXRWWUMlKKrP+90rKc0iOt4NOyNudIwJ0JTqg1N5zinMNcVhoXwXTaq5gtAMSAbmk
BPjxaLKrbt0JT8uI0bfuGQoHUi3Pi9nEPtO7C0tTgqQ7cPY2jqnimad7uA/vWh0N/tTFfqUD7yhZ
y1V7uAYbNdFT5P9lmISK6uY8/tkhndGg/6ksrrNJzLgYv69WlXam5XhmQGk5Jr82hUNiTvebJf13
lAmZMEPS56pjqanyqfB5YpH5IWYTbADUUZlbfbD7dyN3pGwOvaMX4N++MGAe/Sl5Yd1VxwnGsdfW
g8/DOoOrK56keVJcJ2EdsoHAvaP2uXbvOplHolMHBM3eIXy13UgNrBE0sBq89JCkv9LkxOIXDPpx
UONY5tvFdX2SBAMUKpEnu7vZYexgtemSWfZSUNINl4dOJSNPrfXx1oS0tQjgWmW437GUrY1PxKfz
Vzb2DCyxCitwMadPconrUqR+BopB/c4HfINPEZRIGvuLUyyGyEM+e/L+9L84dlErE4SniAATqN4N
Ip0YGYaA729Phg7cfmdWl9k12itEW7yMl2BdsAagP7DcqbTyERz0ZKUSGJGpfVL6Pi/VsL10/tEl
G/wnAhyTDGj/p2DkTukecxbr6QaZfZgz8/KAOTikpJXZwmJ7+rXI8/LskEYodqhsS8KqeqhN2z0y
XApNBVOMpxq61cfWCTMaPkKN2Z9XWHSh+qcVDLlXlsAxSrt1CQy4wd20BACxrCX1S5B5Jj+zrxWa
cV22XYZDs1kdor0hnpL+Rj0qSHz9f8/iVclXhYoGndtJw7VUNE1stZ749bC8WCPJEUEJxkkQU4Ba
ZHZXOPMmhWDaGja0n3WfTQNdN3X/DqnT/ssnuge4mBzTaTy30Gut0+w9sDkmLhVG1cIHXaawcPjW
M7x8uvLORLbI0LwLLObcwAWnNyVf/6FDwQypSr1i1+fj5kBid5BH7RvGzJ/GrIwDNuBQO3hhiTUp
NlMPnzw6AO/b+Ou7riO+ZBmvh8z/6yxzb7/4z2FuCm5wbJGyacMbvFZeHybdvydTJ5OscgBJtTIR
AhNdjR6t1Hxx6F/mAeDWtPwvl9geq+0qZg5CyC5GGany028tkP6Pbipm/pG9+NpkeLQ6g5M7Hqzd
/rAdae0E+lpiAfK7lMkthv2LEX/wfNF7qwD7PzGYOsDaPX7Ln9/8pUW+HiSpmmu3GqDAgX45u4Tt
bmS+CNHa8r55sNKpnpEz+2+pFA+ZaN4dmbrRYxvocwW6pKFm6O0feXHfq6F4J1wWT42PXYe/v60T
X6RV9tkLW1TuJ8ijAAOUhT6nonnLSzhqh7CAATTMg8RB5gpCN1voFhpVZ0tYJWRDnbNMBtL1KE/e
eDAZxrJyD6rgjF0yRCaAUxEMK9MNKoyNB6uEgWX5cEQOveyQIQOSiz7a09QlMBRw81Stzi9kGiRF
6RYVt4HfJs5LN8N6gpFBWF9Lu+YURTyhuEKSd3trRdzHgOoouZXEtN3ym35xk/Gyq3VZpeIl3Abj
b9cC6TD1yWf4Hzth9hZPIeHdjMG9WQ8Lm4XiEJmNJg5oqpoGYwTDWTDsXtXMe3cln4EZp1yYVPJc
xN+kd13JDljlTMmoqFSX3O+FEvdykC+tkxwHyywJ9ZbpXoZhw7cWHKBemAgRFJMJL7FpcoiQJIP3
UcGFJkWLzvIrhQIkceoV+yOrWH8Efwx2YgW9dpgmvdZo99hMArh1opbmVJiI3vSpFaC9MgrrcBLl
ywlAw0TAf2LRFD+NFP8qZBHwJlfAyG0wXHwRKK7Hu3srgstejgAvb2mpt9Ww4+mOR+uaJHZwLBB3
17OiHalz3Btrpc1uHYoPY0F7rDjJ+CaEMismAI8u2/6OVl1Aht/x+GRVFC87L6OYyVQHyteNlILS
UHy1QzfPs1VHmB0bLM6Z+W2DXC0gv8xgrvGs+8IKm1NXNCYSSGt2BJ6/mwaybv/6SLkGg1GB1/ac
jPEYkpJeONIZ6Kt0QAUUIbe4ddYUuV4ncg804fnpKxEsvmSdtWUVrpLMjDC/7QSvqxWIQRGZYHcC
Yxy/CWZ91+6RcLYPLGk7yjlVQvFSTfH2GpznokUb9aSArhvG/tZZZ8kMxYdfpSSVtWVTifPslCpo
eoB7zROCzO9IoW1bBB9YbTbSOwO1Mn1RhzYKKEmAvxn7ga1ddkgGdAf2R0xLzDO/Swq/GgHKnp69
t5Cs6ynalzHe0atGL49icpSIwxw7gmbSnaO+Juddg9TJuUk7aKt7b91vQkhxZehvXqJ/7WNXdDQj
VrK1kZQnueycKVelmrwwXpwTU8xng+zp1iKSHHUItTiYFW43OkZdSXhAyNPxs9KyKC5gUbwrotGg
z2bC6bGY3/Fx7xlDSTvdfkacKiMgVW2AeM4uS0gqTbMTArvSEPJZfOodyr6BHNdjYyMkHbyFj60n
+KijRHpuAPZBZ0O2kLQP16gK8315J/+VQUZsgi/8/vaTFf1baF9W3x/2ipSImwlrBPkB0Y+3XyHC
pN+zjsIncAS6/dn+eAkN3MekpCtJUuzNghEldsEj3yLVMNjG9U3NiiWKxMkpoWu7VC/5ahyVPxmu
yMMC7uN9oVz6FTbtOxfkM6Ap20B065DKhydHkQJQ2B+g37gaDNQLx3s8b3Py7AEImRzHcghfHTWy
W3nsHAdy9jvFUisyZx5DY4wHQKNptTYKdYfg/gmsRixucoIWCpugLEzUqGHIOsVWd1uKUDvQYVVg
a20i6YoEq35ORLYh3YT+qAC4t1gCGvOr50b5HqS7qAqgH97KDKP/04a3BUsHmKHIQIIwYRg3MtN2
M6PpVxSpMSMo7k6kdhUhQHGZgMOqGrYUl7IAy42zOlbPl6IwGBdhjV9myG1vKdcWhTIcgUyAoBTq
4hddB3cCkbAy6MFki0MW/As5pUtiWRX08qlvX/wd0uPgUusyXMeSjPLDnV7BclVvFPlhNo0CEh0K
o/HMM/W5taOOV9Es+X9+MX5f4b9OPs5XDBtnGQJCJQQh1gq/qV+T90V9eR53o8pdnqM+xAdWb7yf
Ngg7FRfJFrgMx8/CvTibDqiVdSPDeO502VvGA3uGXhF532qmAKxEBVDt6EDYI3Yjrkr0DFhv/hBV
MBZnDVpyCZ9eY+ePCDyppQL+I45Z7ve6QwZiydGYdaMf9pc/owM+E0253UVwclnpwJMEjgJFbXW0
xrFFoi7blNyPt8W0Csy2ILgESHQrQ8dWY9BaieFm1ThoHuziWYMK8XyXpKruv2j9S3hnN0di0akm
qFRoO+/HXoDL5Mb/0Vy3ligAXb51P8TRRQeyYQbBLTb7VISQ0bYiSR6tjnO4DIaIXo41xw8fURTB
AeRBGeLsAJYRl2IiLzr42POSD/ygF/MoKVCXDW4d1dPur1r1/3pPnxbnuWa1o51yPcHODUQn7nYv
GhT3kmC75VdxtTb2I0nHwjBwfqG5oVNslRF/3eFnYKmtqxgx3tMz/QSezyilW/UKMdDeymB300pa
9ed65ue5GbDLW5IxQ7v1ojDhnhB6QDMj/lzmR0zNLIhQPkVdOKsGI0DzyBRtYY9JbZijrCoMHY3M
0WKuAFEMrywKhp2BON41xrJ0VoQDzyRSOKM51ssDfy96d3gA0yeBDkzS0s+ROhF2steeyS4dDTQa
dNuL9dauO49yykojHSUuziI/IVfpWdOL132pDQNlD++uqLjUb5Q83gUzYAxocqV4zDIgtSQpixdz
KbzsKTix9iT779/RCeoG7Pce193krHPb/YZKMOvwLam0/gDAqVFe+c7ewU7+9doGwKmnk26sZ4cK
vy1sbdIwZRr0WDpc7hmsxGuf9s5/qNmYWi49MgxJLWsJ5txS8jg+F+jz1qr1HHDlgTJwBMkvqcXR
igF6q8c0Oih40fKSuyCbOMNY6DkZC1tfTGC6fVB0cGk582xe34GjtEC+yiC3HG6fgwCkWzz5XzIk
2G7VPOnc0Va6RVmNqlsmSgiISImLUy9mDZT1i0dlOOJ4JSR3dUY0ReYy+ABOD+G0yFWjXbyyJ4oo
u2qSwVKJqorwo07428KcVO6YFSaRyKjU7dp2/jUBdwtoAilCgdMvQtRT4jMKy/PpqKomlu7Qs9zF
UOeB4ZntMsfOVKyINC9DCXoQ39xKg9Mzpmp77zOyjxP5zejX3PyIFy/iXbpaV75UJa2LwVv0WAYd
XYqr/UCciXMgx7GZfvr5bXpt7e/RWEjxE23uHs3G7IoDiThszqaXWjxRyv0wCVAV8NSUnwQURFBu
px6ae8DpVEkHdsVzlYOJuODnUcXV07FAW2jiZT6JeSjF/ESApaWzVeV6/yLKPlS4i2U8vmDIpPan
5ll0RiQd3iHCDLurOakktltkyeB6yEQYuYhoMKDOloQydIOaB3baE86LFlQ+UaTbLLU1VwL5xboC
HvUaMGVvuQJekYriWPAyN6giKQqie9i2ZwRJg0ERE3pYG9rBy1DNlb9IU0UIvCz6ULhxIT9OCVpb
cUt3sVmwwo5HfIh77wayihKntJumavC1jj2ilYgJqMlPDgHy0mlWGIMgCPalgdpfzEUNRAPtlveR
vDpqdcDPRBIcdU9p22Xn6iympWoh3to/MpBxc3vba/RWvq8lfUlLJgmw5w8BZL3yfyptQWovBqF+
XD+t1PVBrAxE5ASxGNGaLrEOxlHaqpY5j9Po44xyq5q4VjrPBS4kKw5cEny2QbZz7xXgEcBbuF8S
6rfUUKEbikCe4vpmPhTr9NYrW9ZpBf3IsPdXLo3lExE+cpLm7umpsihbIPLIg7d64IJl9nWzJ6z3
ykQKPt2/23HiH2x5GnBgxqeKRuE5u0nBmPjCg80WQyCcT+Zhoqhozs71KAUWHkbDYGDuU8cS48Tf
0pArZjCPkbUzTZqo/swPPJZsv9NHpX16DVLGnfgrvHZRVks+opa71iK2HiCLAICnmC+CQeZEMLdA
jDCxVMc+8GRFrnKlLoEmxKowE+DpA8J6H3DabKvs6lFC/lQJipPkUrQEOp5Tl5pzO1hNGhAvp+vL
N2hIFftXYIr0eyZvUyeS1SCfTD7eNUB5gqmn7fmIwkBNwv0eFyLw8BVtcjJS5XCBZPNKh6rm1r9F
8Zpr0Vj10pJlX4UAuwUWGdgmPy9sUpdeceDfNSXKwSZEMdNIeZ4CnMkDENz1W/5xf2Q3dz0Hni6o
m2m2uuqb9OBCyssd8d8kOW8Wl+aTOCsLNzvK9dYdptxnCvlYVr9LmBVxzTQFKz73GLqdaHDxEYDC
XVt5VT6jJsQkk+VsG7oOcL0wlsEnqynmmL5uUDIN5QFaCJERrZGGIY/R2RtWWxMIQOSZfEitM5JH
bbB/I4hKK8/D31WbchyMD6sm/Rk9VNywJ6VXHGSbi/1HEUGqVYmajaSgtMcotPbLIATLy6ANNNHi
EQtPDuOJz0A7dTJ0RCKftrtxMYul9ul4W6i8a5MGGX3fLJWtRnSFFDEk5vECVp/vbLewtGplpKuY
j6yCTNj3JMcHkX+EAx+fGlrlACIt93rJWEjBpNgVgDe6uhnfkNlhhIN93IMhm155D5sTuj3CLoQB
wgOlYRqAyo61/T+HA7KheNEXAIczBZ3En6ueITZQKnqxc2GSoTG42VhkBTxwQsZSgICzFKoADcH/
kzvn0s8ku+aJdMXTcd8L0eZw7OLEGVmoS80k9ZZlB+ouNO7EEjluBz+re8uIoZ0DiXJ0j6Aswg3r
1Fz3ENeBsI0Ny77fgaPU9/C/mCk98GTosZQAIqUiuAGmb6Oytr9pVIYqGNyzr8Gk30nzCI+1TWxB
h3pGN61bmTn8KFtXLBHJmv5DKVvfmDrX/X/sqHfiApjRD6ah5YQSTtmBXbOiw48j3XvnusxF6yqz
uTmhqymjVA9uqMZ76RMlWVCq4wO7qjRdLKIWneEpCVScr+dz+dk+rFS9dd/sxOr/asfaNkciXHnX
NvT9YtRyEAfZfQDIs1rpdx6Yg2utskrWm6gQ1x8dov7vWBjhVOLs6+OnF2/OBHyKyT6YIB1qkT9+
4mH+iBHVmIWf5n83DU1JemANOwEc9wMzEI5k8jaM8vuSQGvSggR8WYVAZ0eEXZA3Sgw0lyXB7rga
3aChR1hxw0/J4DaG2KKPbx3Z8GmN+KwN5MM9nBQ+7tubqIy6uBormCDBhY0wCn/2Q5WyTx0kmRs3
CTftnvO6LYC82qYGYCMD7LfVcBeSZtgVusHh55ShP8XVXNs96ofL9wmploKmZPPrRpyy/K1fWGWp
ZXY5A35tzADo5O6V2pwpCO+DgWumz+Jh/HQnIO5hWVq3b28Hu0rGZ/4iIzTBSnvcI1gEXp0jLyTh
zz6ikkgNh1R4ntcS+8RqzWXWSC1CQw7irqp9cMSVSzif+9nXkBrU3b8+mB9VIxPnTIAUk+4I4hFZ
fr4JgHwE39BRznciyf8PyErT9JfjoOXsWoj9XaKGSgz1dO2FBvROqHbaQTzBQCzRglGQfL0yhF7A
DnX/xfA1aE7YEJjpKlwfq2iPSo5FUuRWxjMMQMSII4if/L7x4LSj02XOI3K1fWCFXYCXVdw+Fb7r
qI7WKC4YRm0KODqJiG1Oqz4ROb9DoIzBsqPZlpcukFaU98DoWIYzEXsGtLwjSzb/nCHtiG+q851T
G5jU8/YIqWbyRMMKn9//WLUW7TmORBO8e5VH62WrpBgviyLmaGSBF4D2gILfIB1w89iMbzmzYLBM
dZyFY9uRblOgC/ZtdMnOrQI4Ml24hTvTv4KhLAjr+jJn4ldTkY1KKrKFmSBpGTcl2zKv4hNGuSbJ
MjzRDtViC8HEqpb4VscBbCxMbReGLIjHBG/h/gGCXQ+maTHlTwb6clzPb8BuAa9ts6L1WwStyGT7
GxWkltn5OP7mrhGmWXNAa7sSg10o8eL+Q9WtgrCUg7c/7D4sAwbewePlCoDYwbChIkKmIdIIWxmn
6JiULQQJIVSsiYiFaApZ4EkPoMuiLtu2vbx67y8CXLfFjnbDmwCOcE5SL7XIRRYHVlfqu9mh7lfu
AoTdQXmFJYjnAi7WR5x0BOb+w2R1BiXYBvuw3mcJ1Ekt01LXXiWM5aUR6hdUqgauH8UoJPLD050I
PW0bXPHTzxAbYUULApZvgXevaP6A0Fv/CeK8SDf/c3qy1L6Uj1/wxFpSnfYAmM0xmBWySjgErLVq
epMr9impTCWkjC9+3pg8UwAzjkmcK+G8P+AmjcsKF8IJl+UBfHgBQMpJQw75x4b+HweErcrk0HC1
+jhDx0I+tMo7fyvFqMUyr/mF4eqn5M/YIjNZRZ0r+6osmcTxZw7rMdRQYRP1j4400Uu69U5DHlcc
VVxZtlSaBIJVTeavh+v5R6ScKQL3lrSfOiN+Wr17+QqmfvuHJy+v7/3YJ5Cgq1KJuEXonjpFDKqs
YuTwO6sDBsgQ/bER9srVHVlbOUQ33TotD79kEbQwQAc+RmoUvbS4MS07PUhlB67iYd1VbnpKRDcp
KFvfIAZiY+JJst/7TsachEvdsKMgmkILhDviV7MGpBi+aWEIJZLjrTFOKh66MBLRefujNWe6Q06N
1TQwbIRZlzmwez9r+QBiy9XQe5SVbxW1UwCwWhM5uyYtKTZbu7Q1Lvh2Rar/6tIBOrARGKlGGrOH
OVmg8c1ueDQZcrV4iLtjfETK0qaKOCsQ9O7g9tFJx4DABaIwRLLD4kRgh99vkVwmbg5GL22aPXb/
YaehKHn+opS2sV0eA0C+AowJMAqq5jBHRHikvVhDWvWO0m9Vvd7UtrpjUBdwm8N0tu+J9RWYUYFj
YysGrz9ZaA1Ui5D5MIu+yXtdmGwW6O0fp2AoFrLPtiG67Sjf0AsmOI8jdyHvqvegOxJ2UotxBi2F
HGsyQbsCMUTgastE5X4P1+zYy9g59T3XsZgQjRA9/KW/7O+MNNJyKIsCzbgzJNhfEK0H7CyzsXpU
/rk0burPLNysUry90pwAadNdi1S4sbCXSsbFWHF5UelEg2++NTfc0n1H1hvVjT//qSBWlOPXYu/T
d23WD1bnhRFNMBZv9ON4RPSB5CZVDJmYK9INGG3hh2C7541JO9FVZLnfUsxXEyDuRfckfrUHOSr7
vw6c/kLaIeaXO6pAgOVsvZqAGuVti7YSKYs/RqYIlG7lGplymp0JaPTVySOaBLa/aNRpfCqg3nsf
Hg1al0svQ8EAOwyzJ5mYH0hcC1srKd7CwfdCLkyFiK9nN6kcKssu7jJIztSLfQLLzoBdysqjV5zi
1nbt5sSoOpTQv0JVxaW7ni/3s5F3MuEDSotUWll8jT+RJzj+CFpfxoRsAsyNWuFBe+67ICh+GJ37
e+XAnbtXwo0C/m4NFEZ9dnbpvOdFnQOweb8Zes34Nt6aV9akP8JHRqr5FqBHeFIOiIMjTAdE2Wyi
rfGSwyXP/KIJoJEP8cYnRwNn8iLf8NLfD8KXA1P+S7ASy22zMAZNSt+lWCAirV6WePUv5LDof41x
4ZwwlkDZGHh/kVo5ZjDtwmXAPPrqoEw6kdQoOZgVMd0RgPiqgo6EkjIOFxwNe2rUC87MrAcXaEXG
hTyNm5OQw4zemBGA/dtYMmuBPmTMbIGTjM7EgmmtZesz0Y62laLgGq+ZJWhfF+m40pUnXv66gNBC
YH5yL+DprLVxkmoIa0O1bc+pOotwuc184Pq22sOvAdAi+zKo/z3s1aQFDXPzJlLnVni24oGB5Ov3
QvCOGKkOOXzJbw7U7BzHtvzGvMhpOusfAZU5kTz/PkQB7P07LYlm9usx1QyvLHjNXcsQb3naufwf
Jh3UHqc4mMeX+mmvRRcdmX+boSDj32UVFMlQRiIxCh8M/nSJ9eXV9GkAAiXLB/Zat0PofvQIryN8
rHuPUa9dxfeJJZ2YpWdiR/5xXSE8F3PuLbBPYepVywL7jeITVmkh0rB6KMr8L6ztPTFe9wf7b+aY
O1yC6WAIpILxFpUO01eKNumtSrfv8+8vHf1QQ9TbwDEAIUchW7xxcwwVD4FCK+kAt9hClOcjCkWg
4UQiItr1A5jcQVqOMAUcajS4ILVQ/b8Jj0rrAIIQy/PU/Knpt0P5EiawsumJckkxnxEqv4wcoLj4
UdpsHrWQvasqePFLc86zC8kMuOsP3zIBZrbWazJe/a2A0rFBgZAm8tco5Ub92wpQwZ37I6iKAFqR
8sDaaIgD2htkmrUlhOOpWDvTK2xowwFns0N2lVHRBnGzLs2siiW/YBuvFU9HWLVpo7plPNAmgzqf
yo+DF80+zlXdQrjBgjT0XbZtkXwa0a1wlQlZNLQrfY/7bggSl3SHTU0piRMRN0OOWfPXnO4mw34f
pLxG/E/1R9/WSzJGZoZ8sAu7ffP73MP9soutTgB/nHFku8U1FgweygJbW9whC6ensTbBAouz8Wne
6k1DEx4MYEx7NPNBXmDuUi88P2ExPLdCrdfhMOV6vo4Bbc0+EnX8Hbmq7gyCi8wXFoaN9zYC5E2/
10vm2CzCOYR/SeArF0KzZ154UKaN0wwoi36l6+MNec/etkvl3tNrHeveAFmnnzF8v46MQfL8LV7b
UNuRatDvCzCLDvvFFqbAmLpvk5nSxrGRXrA1IKY4jDkW77kp9pqZv1/e/WeTZR94fB5Eq3AnwpZ8
N8K6x9fqz7mdHtJCAH2AtUtNyUu9/d2IMcxLKvphzc5o2VoMpTHC0me7G6Ws+HO53QuoWpig/NmF
jdi05cDc6DYYhqfMVxA3GmhOx8BdC2OHd4d5gVm6vaKGiZBX57fhF8/ekJSPVB2e6HHmAU8OBSkJ
XkI5eEwql5Vk0VTz38zShc4duMYvdeQkQgZVSKU69AVUCpEM5VFc8HvE2uTkD02RYCDl76wN4qsS
uvP/uP69rknJQxVzs7XQjduECVLy7DqvHtwOJ4TGf5hiUlh5SKODCyus5NzXTjU1+04Ls1Xw0HvU
oe0RRnH/K8yKFPB0wgqN6gXqMLJnK8mW1KknAlh8leFCSrCBhhfn4H/oqnV6tL/LDHnhIOBBUx57
dwVIyEBKiedl3S5xGfX7Nux0+wA8sa9B4F3KXl0+qwS3PDU+XyRHAG4BSGTh2jbLHvPHT2TzO0En
D5PKIBQjt752p+j1qd0DroTkrjuUp23hLhYiHW/A5mhsP16k7OwLOSdTXVyknydP5ZzHqW0/1RTG
G6deM2rYRdvYcDVIB/lHem1hpKi05zcvRZhfeKGAGwyEByKZ1KoBLPsxdykqRZDc7VkO+sbJX23d
jFhZlXdgP3Ue0Ih89zPsoFctkjMxApa2SNTzxsEubv/4PU9jK14LDYpv4mvizzwN/Bec0IhXgHU/
Gr9jZrOtSN44PtbKlP2r2e4nAfPDALxpLvcTKpc7x8Z8PnqMIrEjRDHPXbiAmggGFPZNeQ77vnU0
9ny/pUV+yXdfCVCqDEexs4SFFjtDEaL1mIZ1J1Szfec+qAF03TDz1/bTYf7ICjss38BIeDvN3IJq
7icTNU2t5zig2TnHdu5Pyt1hf9bg3pcOX2oDFvoJzl1ou4UGY7OTaPuYAjBmFvFW+Qn+e9HOKF/+
Ofwbe6T4NIMnEuUniTY0ta+3DFQ2bWwdTaI+1MlxTYgRs4pyovdBPCzVCxsE/efi7px6W2YvX3hy
4rfKZ0OdhOZtCyx0+zcSo8bU+mbH/OBtfgOOJu8gVC0ctrg4o22QWECjmXGT7Ipk06XnzchKFD+4
ISnWjghgk2JgY8CatiB4sRks6I+CCv5J5UYt1GgZGpFot9tssbHPSPcSe7ebBzWUa/hBPipW4NgC
xnXzIRl8BLhFYnC9dU5b0zhsP37ittP0+0apB9IMIaBcOvoZ+1QxzGpFahF8dutYuy4FizS3FjeV
uCQDg/kQG34zLv4efwmkJbfDbAYMbEDMlCnV+wVarD61Tda3n8zKaJVnPfvYZMZ/1qX9lYjFB6ZD
5gCLk5J42bXPs3vGJpg/NTdKb+OfQzsTITjM48vfyjJdjraA2tiKkyPhhQn6uxuJWE12yX4xQvNH
+M32VXRA8Js9ci4h6x5x7lneeJYcTnttVns1S1n3UX3k6O/x4hKOsW77RIUgSkzwvZEdGaDxV+ad
YAUK0NsBEMXsy6S06v8WACTKlc10WtlHzaIs3c/Do/DkRrGXquYpzRt2fWXbJAotwjL0aM44Ii7T
XHPGPFcyDUv69GiMe1+lohvEG7EkBi28KbnCiPWjfKPkN4Fycleixy5et4SRr8041p78xK6OJK5T
3JrW5yj4Z6lNATPo89BEf1/F0XXUl68LQ1Gjj3OmD+1Ndk1LUMC7QvQPF3SEyZliU/8m6xXgGjHs
dQe7ImJJjrSWmObxCuFbG/i5JSmo1rQo2uKxlVKNg91SZiMwT06SwAbWA6clh8AIs1W91+6B15gv
NiWl0ukC3z+ventvQhXvXjV9HOFpkByH/lZUgZqL8atSSOOihkEjRJZCqT39N+BWExohWdUljI3T
OLYP9bIQi7OHQWOIBjMXo8H31MLE2z6XBlWcC6yFTGx2Cjs8DJVYa15OiAhSXkhj6+ZNeEpENy5o
En1u3NIsF0/cw1yLqSXv5i302zPwmPAax5vgF5Z+h0+DeSKTKp/aCMOM6DZBFB6/mV0FLwAcxnvf
tMHGfHssiK/AKYZHE+pDXthogCN/kdU1cAViEaelk49tfEj1E4G1H2f45cmk6UVXWYc8IA9uv8Y8
zisbeh5l/XA3nxSiupJ5SW0DE6X2rM0UdhG3RiaM+m+OyCPT+ClFDFZV1uQiiIrRiZWn2v85QNfi
jZmI2kmsmoYbia58ZcNA6Z8sipPensIs5KoPMaZl5H+d+7EbnEEiQhgCrPfvPrfbElbvBCRY8PbZ
3uhZYYPZ7Z2yU37J58YaYNGsmOnibi5rA3B1G0gdDjXvWT4tRAzgrF7GNHzqfM1b5M4+Y8oBNS7Q
qVueCXNDugHcaKJFXskJLMPJGp9Zd+l6zbO6y2F+b73NFUdWcJfQlu9B2uqxeQbgbcbkuZIiAS3a
cy8X5LYdQRNMhftIisWYKwIMiw7ghXjJ+95VCvnHKcSQDUh65b6RPzlCqrplLAzei5CXHkl6xJHE
WX7bQ7Umt9YQXfOP589a5jxmCNJm9vDmXKdirWf0Goz4PZa+oATQuXb7RM4BVHL3KWWY1BjW8/s2
PfVDY2XYSsL8GTZYOjm+Jh8ydCEUpXjyff9p37pij81v4mTzl95azcrPw0wPoEwekkSIf6enz0nM
sGHVOZuUHhoiY7zS/hYoMFY9JiiPpUw5hsjnNLbqnaa7pXHgONGv3mML7bRWdagvkwwuMZH4elxq
k3Qs7fn0OYzEv87XxBVXBbZy/0fOZbphtFroQlqXlfVEViaA5+SewS/bylcfMEMEAfpClFPzjcB/
XAmO6ic3XZJcSvCH4zd+ZvwprmcHneBpEW4yUXO+6km738Xv5V3eTxlzy8DADGEdKXFFXxCXqkaw
9McnIC6YrNPHAm53BucSiqjPCNjw0NO6zOeQF6FVrHBFDZXZfDBuztzXAWXchA4iipMjtPz0uBhU
OrUmm+i7ndrs0C+pgQOjPjEj9svMcXIdZYEo70cqdCC+cg05RXMAzEcGXag7lHvkhKEqBO9VvVIx
WJ93P3aK3DbzwSNpXgamqyuwWl8kdbwKCyYmqLy7B4kd+FmUdXzwvdeIMbhFttCUhZOzp9LiVf3W
FMP/CgXmR2zHalrBhbXFRdtV1bhC9knoClTasZskZYZ9GeJPi4lyf74SZDT9l8e5yJ2R+eZt/PWd
KRYVkikEmwFLC8sWR1uJfA5dnIsPc0uyzhICwRaEg076G7I0T7OVegm1ToiyAhQ3f4afEmQuEOxX
BQTzbfO13AeFfvEpvOVwOKrvGs1+gNn6P5mE3VScS9BNuAlT07/Rj0Qv2tjDOjMqBOOOvEyUm9BC
jNXB19wTzEhdIoFfqG9I2yAodVBtaV1K2+C6YwYj8qqmhhQpzMxIIi0gRi/8AYpIu6QVcfiGq9VB
+CTq+07yJ4C5N2IIwvRTlAIc0rLCMOxEJp6txocZx2eoTY1rZLGUDMpD4CgQPN8yre+p+RUmsbJP
QlGeYqamDCdEnrCZ3D8x3RDnoBkPgbnIYmU1qztXtJuO9eOMANDokeTltKbL8wDzx0qmrCT6Z0vC
cE7dbJgY9B0+MHlo6SwN4W80RYeX5bVbi+isPlgvAA74dSlIdXtN9Nvx0t9minYf9DMNu7p+350V
X/4uh6DGlTUGIJ9bSbvV9BAL5wi53ndSzwv0iNDAC9rZQuok+8uJmTRLSdOB+eM8kgu4jFR09j84
RhkABbdMRoeMlhWZy5VpxhcP0LySxAZzOGFm5yYxDIEzrZHGgQk6BBc0IL8/AvCLTebgb4qo89dA
Okhb75bT0GXDSpGD5x6BA96EASuf4t90kwoA++SKzyKILSfMMnIZiUQupIldbizJWIWcDunsE357
anLztPg1Y2EOjsTSaL0i120IZusuIqU+/k4GldVg0aUJU4vzO+ZNCeiF8qJIeY8otPdKeIOt0Wkx
QQjn+w9gVJb+1cEUNGZGYwsHn/JZvLVwtzTWQzoqY+YcIOcCD3x9WbtpJSnc6P05k277nwMax6E9
WEFnEI5/y9uASGzWqv1PIHM/GiigcQ9BrAhZjsuik3sl/tjO+eLB6kL5xDgM4jUDJPjlEHYKWOx0
hVvMq+wKBf5HZ6yBHbucSkI4yVKMF6xRlEEe5uzRSukHmGFitJ14s6mxxQdXuD9reCzX0RQbb8ja
bwFdGxTI3fGsFgLWnbrz8FC6DulmJbSM2HEFsc5snEowLpWwBttxKbZ86u/hLJienYmUDffYtMyp
5tBuYEXVmP+X7Xi8GOOQJZYWsadVtQpgVxlQcYQPjYFnDmIaLJXaJg6JA5zqZmISGkdJ+hs+GEpT
L+/aqTmDJabsbeH4ml718FA8XaKcVZ6cSm1QZTbea0vqA6y7dvQ6XhpKvvK6Yh0qZcMM9RUVKKw/
Q1AZbvUYbDA/qIB3li8q/Ytcwo6EoeoU7Udohw4lnBfT/rh/5bYFnOFL6wEfzn4cSUvxTC/zWydm
NsNsVNM5BI5D/sCjweKQ7i85eFYsMTQ/+LvLomBUaOBQ81kfWA2HX6+WI8ymkEBux237XDZCGMzH
Cx67S2PZi3HhalN0nOur7KlWaLf3RxnSWwQXeLN8C79ZmWCJxY1+yGeiSpnUm/nDsVR+SwLPOhhg
LVhUjajA38W9Tzxk7lreDB0jsHSjMTwsEKuXv7KvxMGJOns0AmdJ95pWVw+zJQy8YP8tKWWQOq8n
6FApl0F2AtiL0W20DjoqJSKvIPpp81ddvjoL0IiQ80HvT520/mG9qaHG5T1rBHUyhdGK+UMfbHFv
zor4ipT+fjpZOJ6ncJnf058m4/p9q2GFHZ37pfYFFEOcP7Xl7Rv7lqiRVZ2p6a+FxMVQvB0KxlDN
AqLia1r+rnKbZXo6TTRRgi24evzmL5A3RYMxzXywvAZJ1EfWQAA8KCUOQwIeLQuAatY7lAVMU0fx
rxIWUnpfUyxZPXyXXQxiy+KXTroHhmhqT7oC3kljStxV2ZZ2jInn/e40mi5E4rCT26GPwQGC4QOg
Iy4QCGuvza1xF6BmUJf7MIHFMYVbt4YhKf9U7/wqW9zn6EeCQ/N6wUWFkmJaBR7JSNjgxdT14rEE
+4SjDGywBJJtA82tRw6CNPG7bYzBrO82Hcom9CrLkluqtxO5hoz+WCd1aCXePAE5nT5WzjXkLREK
0qO6J8J2twOzo6f6mk294dBx3NSWcvsoBHDDdvmRQdSgHbQ8AtOP6/zC78rpmoX5Tz5hjkwVvQmC
O+1fib9MF9KKOeD7ca9Ok8eGVKFR5b5x43z93lCoZCAYdTBF5reANPYTJ6NfW6QZ6GDVW/tkHtiJ
Rlembw2i+VxGoCaqVoLwTbYUoSFdmi1d6118eY4SfSlwmXPMbs5pVQcFq9vD3wxPln76i/dWI9sE
30ydXOsQ6piEyjIlV3swOQ3J9gb2V7GYkx7HaEBqGllVlOD98JboxnvW3AGQHd4LT//jBP8aV0c/
EpwUavy2i/ioQmFf5p3a9ykiPdgAw+Lo5BVfum6QKmB+hcj7+v5GGlELJnedZLyoycNk3nvwdjLK
/j2tzWK+3RXMcdTRdIPgZmUPAnbmh+P8QoHcOkUYycR2IYgsU2y34/o6mH+Qct2gD7wKKy4jew5s
nneyIs1RL9ARGGex6lbKWcDXy5RLHBOuuTcXjfs2xyj9j/NaLtkN3meC7MOO9yGd0GCT7/m/YE0e
hGl1XkItbdotRoBfaTLVug1IfTXSFXELd9T5LrTLptJu0nl1k2ML5m16jLaKXaN3rhOep4rPskMd
b0b+EdFxlJBdsXQCPensEXMbdVXKun0D56b2vtrnIMw/qMrkXdWqGo0fjCW24q6zCMgoIfDV4c/z
SLK1N652pQ2OAQNIj1nTSZQM7zPEJzAjuEF38CCgjZCw/rqO5DGpGIsvUs29WciQrp72mNDIAp/T
9DINaIiOmeKQp42JkzCUNy/PXOTC4BTIAGmsjhFJNlGVuej2QX2U+ZC1CKluBNv/9Og2z3NC9hD0
eV5+aAKtYc6r3apV/YaN5La1yr87P2TL24x6zTKEqsMW6l09EiHVc3QUwkPfv8FVdHBN+VnB+3GT
M7jwLusLLsVUH+LK5GjmHLEsU3VuYijmDSI44j9wPZzRRCXXkqKwhA4sqwxrj0K5st/2ydMOq4P1
aXodAvi93O+aZK6/lOnhLtZtmBtFlg0kJu/myHk2aio3mJnZgung50HDtnYFKFkNtxje3QSNy4GR
2x65g0h4JcFrruLyX1F23lIDFbsrMTvQZkiKmQxBqwIh0yUXinFzlbC8Jy/rhasAdnpE5CJFg5Yb
4Fv/rVPY54mBAJwtE3kCZJLUTSpdtAAEbKzGZNRH6j8+Rhk95ZOGqDE5T4gOylLjJX1IbtQRtEvt
fIinql8dZ+epg6Ys+lIn2EpYHaweB9NeZ0Bqd55MnBUtugt1LjmCdpZP/0zb2Z0eLbWggGVZNIOz
7Q3LEjB0bKAm+tuS+ewCuTyqnleWlp6eCGwledBPzCIgpl6TZA8xfvE8RTzXx3Dt4rnh837uwaIj
50jOdnjAa4go9Uiz314mH34yTKsQoDrw9WEirs+dEuW6QF9Jv4Ku/edvPkJpcVHOiUQmSdEmYkfT
86KAyhj2Y3q3keELH3ldWUHbaxYeFS5Ik/yGSNQ78H+4cjQTDokf7EaG/ffH+Tklzbq/0lsOE6ef
tfKQF8KJMErE2H1A0oROUhJYGuy6MUfOay6Sjr59xBUfunRPfQgys5PnuKsq/jsFM1K/BiI7N1ZP
86wTrsCudu5UyZ0fBZDRMp2BsJfEwLw35Rzid3sktNlcN6h8ppwfSJCaOr1bsjybbN6icWci9FV9
r4JYC/Qu4+RDrrqat4e1s0gp+XWHH6kY7MWPa8Pa2JKbROf9iBpJ9vDxaMFZZ/A+XGqcXNthRTav
HPWXPbp7cgziG3/zmfYjO8cF5twC1OkBmSroLEDPW0bSyKxdywbqH+4nKKzgp2o9NHHddxADXyHh
D+A83LCdVU/1ih9buaSCtR5c/s4RxkG6d6lnzB0+7AoeVmeNu6oZbc+34mQ1JqIJAk0vQIVA8nAJ
aYNT6Ngbw1IE6hdKzZ/HH97dFVCN5NPdnUH+JgHJ0a+J9cJPhooliqhxxSjRd44jQOk6kj5ajHGf
qbr3qTISLz5H+tZBcuIoFAfOF7eYAFKbJYSTYM6UE4syszaMxQ7U/QjVA4p05LyaPNVjsQdAQ3z6
q+g8h7BsUepJZigKENUr5zhEicUXHDVyPitdwVABNkIHlVQmIBMBeKh5uGrzSkR5VYaLC/f0SVp7
E1o18kY7lTcOSravmK8OItCXhW1OKeJh1+yV289i0K3NFVrS+y//AKnvcGPmSLOAojE8V9yIBcea
46GaC3JiDjedEW7IBMgerFUmXks/alv3WVntNsFEDj2xqpVEP+7xRBwP6ZWkbLtbiHlBXBPBgzC9
NQ/SdEmzbHid/RumIHniHsnUr9qEKMO1hShgdIp8mGdAgYL9oNuJQ7Bgcy6P/03LAWO7ve9m4UsE
KXaFZvpO4iqUimbOPZEikFELM9Yj4It3OCo1YomMEEKkMpMI3di861/zA11ToMMWXPlNU7FTJD/Q
jTOaNxBBeQjhRDfz1Ie0lq95fZyM7MZHp+TXaq2T1ZCttfRiSP1bQSuSjiWUbeLCS+JWJAaFOLDO
s7a/ifBSXI9uSWzO73lLlcb0oEvwKdwPqpQ35VtavzSDRjMWI358SRc1A+iSdp5ZV8D3QxhKEoN0
F56Nne50JXlVpzsTpewHiwrec7phelv2wuvPEjkXs/+LcyySMX4bZLrYlEWSUg8WBBIFXJVPvWal
Dg23idUeekEy1Bj0PhTC6th23AxQDVd1jntDW6aAq3QSrWzdXPy5kouwjPW5kkuAfczVFFsApFdZ
hJsT6hjwMr2WZF7EZtnQK9QHDpFmIn8SFluhOsRu1d2yUJ65oHh9koJBvtOHQo8yrb4j6j7uVCfl
0SHpVyKZJxH6rxV8Kzk8t2LKTIZVjJwvSbfylAejWjL+VQva+VF6M5a+zg4J1zaoOc3ShDcIj3te
W87olf9tWUoCPOgVDlxJiuQaqfO19sVq/KkJKFRDkarqVRw7zA7nRtEoT+3cTTOVxaRRCm1dJLcs
DWGRIXCGE0XPJe2Jhjd3rwj09UIS84soXDuO98L0GqO73jtWjiZnRwsR5/IN8GdNXvp+Ff0EAG0w
ir1zSeA7w+7KT1TxXk9o+Fq8HhVypTJ3GRUcVpsLbqyTUVxGsjIo/LuaMEVo8kUvRn0W+OpNozlL
BZOS7o5lxdrS6LaeLGr5FcgRzLQuCjTcz5RDDRFIPkwzazpO9tIO0qCZxkCtzm1W9Lr3qX3UTpCf
dJQke8I2NyPbX2PVh2ulo0Xs1RvPjlrAA7pvuFLBtf4zxZ08wD3o1tR7cATagaSNa2aiuPiJyeEq
3qHd4I9bp1GyHWcl1ybIqcoKmn6q7/0Beum3FRJdNcZbpbFP6X9OSclMyWnaVYoTycoEzFZXjwcF
pHFcRgIVBhIzy9NNr69t66Loccj4QeQuqe24ZExHNBjn0Oaj7fOI2OjkV2fKy8sfvLd+8xAxhEu/
4m9gfdBhxZifiepSn3O97hYlvQ8dWP1GaAdaouJDN1e5wt1UWRA7vWiUv3rdj+PBKox54M8ndCOZ
shZ5UbBYMXRkPmTNUBpx9taTLaw8SYrsDfmeH4hiyNCniHq4FNXNXUSyj6Ehrq2fHdjri6HdS07U
f9cSOv37VMb1BKWz1T1kHUKi46Z+riGF+6VKWdkjtstdbuHXGpk7lds9azoWkKdmr0X01Q9QauDZ
f0EMgMwRKyzwAdfvSO9oeh+K1pzOMUCR9M30vb7lyejcK1X9MNkIgk+BRUYQC36piPhJwpmeIwI/
+9yynzJOSAj0dqhIF759Oik5cnYtldFvbehW9pQof2fCprSozDcbI8cIAeWp8KRHkHPS7C9wOenG
ImSw8JR0Py2emOK6cza5D+cPWtoQY1atx3O2e9BDc7BGh0v4VGjLBeTts6uE4CBdot9aY4dih/3g
HUjikgPVnJhIWSwbJ94KQd2gfcja40y/CQMieZGVrVb05jsy4FQEq6bxN23tTi48m14n6GExGyrv
w3EMxvxUE8Somt3dc721Yy04V2uUdKjKtTwmoGnUs4ocsCF8ouPYGNADirtWlwGbm+qbCvxJ20oo
LUNPJrD5MubSghIll0tBF6fVmmMK/UowVwBajnpumU/UgsOPpgNlEDavODmFiiKbI+sYID1qsRVs
vGGu4mqJmyHazIjZY6uk+EyHCU20jiUu2Cowspox6KmVsMbLnPbTpefbdp/yj2GpomM+Si/BKsNX
W/LdfP/TG8KWCtrrL4TURyFG4wRd+h6vL5E+zBY+2UZy1hjqZce+m77pU6IoZ3PdSVOHVY5X0oen
qdUYVt32EGqwoirzIqrGyTLvkaitHNl28CGX0wT5lN5WZc6+Fr7SozG9G5lbBuewEBN37kqbxGTN
BBp8Qim9kxMdPCiw42JXe13mkaa4A46ae/fAhw962uUEwyixF1djboeK6FwkzqetdoFd9R9wrthK
T8siNlH8SQXY3ipd4Nd86HrXXUKDFXxAdYc+nGgdfL41rdwV6YPgqEJssfE5Al10/9JhzT7pnf9j
z8+qun0We/CT9HBZ/eAGpTlqUFBDc06AOtCopZovXIs4HAKFYg2vJQyYGChEts2IsAAyZL6PRUAj
MnRY43xSGPulT9pJImbGN4WFZizfmF6vEpoxnwX9crpFQf1k9PaIt7sDP6+kWfcoAIt2HdouxLZx
8OnBlQj/CWD4Q/5s5CLGm6rRvhZrQRHcXWEYPrgQzztO/iqX2V/DzdL+kKHesrWMH3gn4oORgB1Z
Mdroj0FQ60oKwdpOHjEQ4go3DYI4DdmfJNFPGlJ1pnwIQsYyvXZGi6mH7BjoPmNRgbn/HrADaTQg
UCEeQ8543NZCUtkp//IAiCuacvZwqatIYGqQ0a6B79nyZJLoh0pQzmf0QJ4iU8CO8ijmdgLkNz2x
6q+xgKK1U8a/XdsmRCzlXWtZl/EkRMYLRSk7RB3kpiDCwg8Iyzlx9uMC0P78LB1Bxn4EVOJocX7b
cRXAm+BFqJi+97+erWy9Hwug6l/IGrf5bHtOw03D42MJUcXUOEo3AeFlP0TD/rSNbL4xnYXEOtex
IvQ/H88p4bT91SONGBkKlY5WkKyYOA6VMR+ljGzDiNW7WdIDdVkhvhln3WjX57nVEXTC/PIh30Pw
0CHuMtmBzSutMJlOcCU2xBDhQgQBwaPdGYoV8lo8muf2gcZxsjhPEu5GutwRgOW20XXgvaAjaHXz
fy4Syzcmlm/YrO5pcEhsQWu3fGScsHAv3sAhRRzM6SRNHCA2ZjJfy6/m6y9MQEaQwyx5A0RPRRLH
xvNUyOYfp6vYFndYBVqi+z0kUKtjBLOkxbGVmawEVdNXeRl76/8Fd4fehD1nmMCTJQMO4S3Blg3Z
pzJ4Y7Y+ezZNzIdD+dPCHiCcy0uTUDHGZ7rxhFXcQpXnnpr6xLRHaJaHXYY0cZcArLGYjWyUGcYs
zoPrngEhpPT0Z4VR/p3xP173HTk/KVhGdzZ+rOWk8lU/1s5q10eDVQxMKQEneMKxzJiejsROFf3T
8hjJZxTwXMPWR4PBX9KIk41c9/GM7ep6YJNAyMZjQOLY6DWzq6Xuv1GL1H8idJmTw2q9H22aSvAW
kbx3z7NGQ6dSCKGjWZf/eI0o+FGAqejMWyR0qH5Pa6nxuPCXxzR59KHnMDDLOZSG+IAcc8jL6mAI
6skfumy6rXgMDmjFhzN9Xpn7TxhRgbw0AT80/m1HIB44OcSPryxpiPBRw4LJpD6FHRlhWj7WWi8g
ivpkB6nSCPJwLQizWuLYRTsp2MQoMmHZPltfink4otRRHG4wbd3oUP3RyjtChkFNUJ3H2u/j2OoY
MGbkuZKPQgWRxbXY9OXPicAdAb//Ua1TTLt0YbI9Wa9yPzAEirD6O6Xpkqa304GIfBJkcibBXxiZ
sbwOi6eNWpA8ZcUV5IRIBNcu4YbFL9EX4wcksjw3lyJgBYgHq2gwPYh3j60LbSbHxcjUD3Lo6WUi
cuY89YX6+Hx9E6YWb4+Uj9G68dpOqbumJrs7cu7TMPjyrIQUlJbezP/f67dijxsOmhls0uDEkYNT
W48Y3s7nmrbHTScbBCGrb/bP/lq4pvGmdK0vzCnusHBbhB0Ayz99FRDmQ7rgg1SF3gv3AsEfyio/
fNo5uhQyHI+1TuKm4X70gxLuS2X1tf+fsVJqsG2gmnEjvfGjpyptomnvVaScedIA3bqVe19HPTB1
wE2gt2XAhRvZWbwwaEwDT45S/lHEueaPYqi/GgyqWOsLVlyOYxYcCelon+ykFPzVcoaL+NozqzLV
d92KyZBkl3Go1f/XBut/ZXdGlNfw1tDfEWcCOc6aOXhGn46udQ9FFveuEtKUxThjtNlc6uJbvioZ
G8Xdl6IrPX363Xvy2LCIYK3umu05VizXpaiK/whG4xy60SDa9ZgzKbqeytDsxhsv+WTd2C73yMMF
p6rQDjYE4h72z2dK/PzRasDVlGXPzIbANkHjKtdl9RNpCW36jfDfF0MXrvmIufqxtNj4DcGHqhU7
gqJoBTM6EGDa1ZIxD6g3eNVGj3VVR5iXg2hnoHJTA3roSkvDwg2VFrjL+emvh5j7gzua78Mv9+Ia
azaYr2ClxyOEA/6ZbKsbzdR3S5UjgjgqvH9XKq0JhNEDaRr9mHK+fngTz8DdgigaRqPkgclYlvAo
MX1W84BPVH+ze200h+yFMIM95spRIs2CfWNRqgUOedn8IRCA9PL99MZz/eIQopxG0dMdeBKwF0yG
GWBk9i3c13AzSNuxE++MeosgX0tjSYfivYvdOnzqFgdtiA1AOfSX2vSTvyxU5zAQ+zUdOMr7fl1j
YsuhP2zMwWa8Hj+NTNLpAlKNuERZ97kFYGcPFQBFt5X9sFFbXrSwnLymrm0krGIQ4yrYMcJtaDUz
qfSDEf4Dl6ej/k+/+G8XQk6OAxDgsOwy6EaTc+rIZapoiCj7jH1soe6ndMgbby8zBXvZdSNPhlAJ
wYH9jag7g6M80igBbhtQV+H8EayAt8a8teVdt/gyDS8Q4iVok2sX8KRJN3KJn/dyiSm79wpRu1yp
3eVGo6/A4p9JDOlVmj02F7vvI+yknhAlDQUGGn/QcN5oNgZ7Vq5QjS5itMud1LBLp2Epkh1Wa1Yw
eER2cwDF/r8pvjYx6c5+X1uB6mOiZs7udSUona3JnhEdRp1oq+j3oIIYWyiqDWIWJkdaWhnAGU8p
/REv4A8Wj4IEBZyYZht2Ujhk4mvFvuEmJT6uf50SUeFEtpouh90t/8UQX70xeCvuZXSKaOcJ+FPn
a2aYM9J/PSZJGLfzsW3+W53K5mBAMVrqAcSbJPFH+21SPvGMqSPkzmfnIstW6QoNLUWEDKD2nUwF
tquoGfgDzlzTJQwe/Cic7aR2Tp3qCw5u4nWrkwLn/C8H16lmJiLCE2DNi6NITVuO8l5xhh+z4P9W
0ESJI2rSIfJX9WdQSbIH6nQ/6ncygLKS33xzQp0jP6xGWBNq3WicoLL3YuIqguNNsnIuxyzX7K1v
+Ik0hQ8+dm/kX3b87016zAXY3DAf3Was2ZYx8K3+y7Ie7PW00BHExSfbFSbjC3HEdXz9mUS+S2ge
3922qC3wyJIyc5Eos0X44DF8ll9PpW986/7QzHVEHheB3mRkXKY4UinNeIjyby/BNv2As55DZs1R
grlY5AWzpzK5dGDUzGIEP8P4KTnHZju+l5X/V+7Hf/7VQGVX83lLYeRy8y7qkH05ZG+vEdsKKpEF
oZI5/D+HVlPkx5tVpC6tVafzr7FKRFTzE4p4FT049XV11OicG4q13Cgs+03KPs+tWB4PpCz7I02N
l6fTTnsPCG4oMeW7C5oZuNsruibFTTOiVUtMLA5WZnQ83A+bApQL4TYk+CL/b53jjBcxS246uo56
67dVXbUph68OomeAsbND1ySU85eiOyagkVEQxRQwieVDnUEMwIPxSMbRFAaP3UmmAWC7+Dd2h6ml
xSeteIVJv2g/+bN/8VfZXvzI/ksgIVGCcAFSapuW3rpiU7ziejOeuLHNerV6QU16mVAy3PzDZ3qY
PNEPz5TMAc13EPRT1B/1MdBFMds1uIbPjj7cKsRSHiLRslcTX8KNXdJPj5v7OUNjq7iTpFeMHZC4
Y9dPv3NJgs8Ui1Iz3qpKRGqXIKBGG8XMBqoSn1KjgJWUdbk8OBvloE7vxMm4ujvYhwzqefJ7X/Hy
7v3Tk9yf6ct+Ig9L/H8sbOA6SRcwdPDNIlu1PXMlC2rNvdb8u8wC7PZZ4uTMMV+zMXLdJpDFOW4X
6Zk5V8knY90+KICkSOeFPCzcs+WxXbQYcAjS9+FU5VNz9xRKmgrbY/DSf0hIi0nPY3Kkz+H/PfJ0
8HVkHeeX5rq9XVnMpLdzWkFNEU2haSvDemLUe57OF36j6UUetiU1/DevxbIjGNv3UC0DUMAj4K9T
BzVFAgRpe+gGc9e3eOuktWseMvdMGGz/Yp/ezyHSx9zZdrvmexRlY+w9+VJ1yO6y7Z5yQ9wNDzAm
KssNe3gfcynT29S/+9FGOe2Mu5j006EK4r1BvFA5VxWuUZNkx/fcLPbyxHjI9hSOjo3bpf0InAxV
nzCGdcTN1T5wV13cjG/4RcHg0lkcIdvv4DFaSPNzw9L2fsN6Lw7Xdob8Mq2mZVFQb2GO9U1XE4TC
f6HGdXVENfZ+2st2IUR5t1JxrPLRg2NMVSASnpZYHUeKvmQbU1PSVbqMWKqVbYLORR+6cVz2IvEQ
xp/ylxu5IYuPgwlAZ4TMZ9o9UcMAn87bck5kNxFlt4CE21Ki5kQFEpYYZWCEwZLY2uCgNHAG5P8W
nKXopWxTaajL06scwpSb7famns69tWvhWZpGuiGifXGib3BvjI9ert6tIxk6mh9B1N+1ZkucGcrI
DaoT8QIKn00IJewZfmlbCOF5uu6vJcMDQl4xnntjZSlsPv2e6tX81+pXDLusrXn/sUWit1gguAoZ
IbAOblPqUJa7MknmXRwfgjLd+gkgqXgC7rd/qn0dh0Vzx4Qxx2jLH7HboULo+fJXO+S9skFyuQ+r
+/w3pfaPBIR4nEmqKeNUzx4aU9EdINC/mlRX1MFrcKX38yijKpqzvlnA7fPYRTgOYVdKbs9tJWB7
r890ne6jETcNRBN8K4xUdu7MIzmbMY4tLf8lvh4LBtKC/gsGFILO/Mnj0PjmCMYyH6eEcDr/b97/
nfIwL7VamLPKAtflhaCCvBYpPxEhfX+UXttkGC8YwF8jGIFpaVPLnEGdMbsMLqml3tbiA30duvjk
CTAUy73Y7wptBrl3pSqLm/QOr2A6yXK+rfCuekrZtxg5GKDNR5XedNUUBQIEaY9irmDLzIAmbrel
JCgq2N4Qcd6XXFGTBVcJHpM6nBU/4E0UAm7V7IDtgkS+B1Etb+3inNcQMkBDX9Eo1WaMx6CBEMRD
/2tR84hJv1N14fmSrmMnK8ql6XPBUIDIkf6l1TaN938WHjYIjq0l72SCsHpr3o0wwPbpXbQ1OR9c
p+uvHAlPFZwX6I+ZEf6njIoazMebIXRqvv0Y1vMRc0GvCZN6NSMijEVKiJK6VjNGQ2nhxBSEY9vX
A39tu24YMtDBgTXAS8G8N3KnTOKybOoPs2GeVI79ELnT7HIcfDJVpskAMCr4aZraKTR+99CaN+Mh
1yKObN1/hS0wDnvm6qt4KjmW0SIRaTZj0VLjwFvsfl2Jj+OOLz4Zd0PmWK8qJAc/J3j1ClByXc0/
nIdY2KeSNO698ojMEQp2YWDn/+y8q6LsQpaWpgba0DM2NhSI7gPjNH5PY+ucZmvUCr5BTO71fY3L
JmJalCtgR62eguxywIsg88Dmm0E9yxGQ6ecUcDzkp/Z2QtjgRo0ce9cjulBZYRRW53sKTdG4iCW9
4i1NuY4GeSBgYaLMj40Jync9VuAjaLiV8Jki5lNjBd6T+gyBskV1qZPHBSKASTv/Z4jTnOXavsNQ
o8AHnx57WFsDc5Z9fDJPYYwh2QCEBw8zJVblJ918vrTOTBeaI8iIzZiMWpZlscffZ7mrLce0bXfe
RdooD+QLgNKt6tAXq+nfUiSzEJTfLDcpPS4PAQ7+GhqsNWz2KScW+yZSoCbEqSMhhdDBEQyPwyi/
UIEdE2oJW19tJrFXU12Q87EB3d828NPX4W5rAvo7JdNOPSByA0LOoSO8koT/lheKngHSBqkPQaxK
g8uozbNd80HDzvhQ9YehZSmWCPVtqce5VAOixORjwVyFjjjJQBuNvYbvMHBLgEdShyZ6fmZlw5DN
UZdhD8nsFuIfo/w85CNDqntkRvU9BDnPmv/aMv2nZ+yP2O7yrFc+h0er0BH5hYlfzSWxaKwQWqLd
xHJ2QNZ9bXuBtBbmB2F4PXyycxjlSfTXowJYCFEsT2GPLdYzknTbTSEEWKRETacFGLAbF0DEk0Fh
CZzxnQosQcjqPDuC7oq3UJHiryuDn993ozJbqSQ6/bEQYRvRK9Z+ASMoOOMwGWoIA1xye6pGG0Z8
010nGifG1PdH5sxbwLOcgRAPvkbImDW+k8vWYI6r08gRNm8zUp/vX6n0n1YeZX/Tw0ziiOHxG5xv
6AI8A3m0+BxBZSyALkEmGbSr2B8kOvIJy0g93Y5dfEQUosYqzbLEMsJvaJ9VI2hpYVAZKLfBjwuX
7awHhUF3r8367JMQlaWeOOkQxlCyf9AHZ1j1W9IsdPMT72A/dontd6e15frJ2WNLDLt16BNtbmd1
4RkMi1ykURfdo7jK+tsPG+ytxEWIkdVjQ3166bDXGPpoBTpnUY18dOMC1E8m2koRGxVM+uGBqGCF
K46cnvTT1nZphaFQf3tMSIaNUuXxCJDcLYkALNSkZLXSinDoR58howGnXtMK/Kslb6MzbY0lO7GD
OdyusckBhUnWyscUeJUz81XI1V98zeutjyZFI4d0TmW+zO12njf+VJOofXYIF1ab4uHGLXKz7tq1
EZtLeQix4xZpmt1954Z1y9RFQuflZCS+p9gB3BccRTHG0Rs9CK0xB68vXwKx7wyu2ThqmSkK++1F
h/pLs3iMqpEILFwdWiRBpmbbKfCWcvzcCb60v5+S+ySfoaxpg92wBLcgk+F6m02fQd5gW3B8hKHZ
YicMu+8dciK7064WGyAbFurBpDdQsLOVOasFR7kvj02sL9UF6mmmNpD5GG1wCaoR4jTR6j+SbFep
XRkVSAtwk5UVDzUogt+GEm22CR0IOap1UOjg1bBeWRpEMA2w0p4xWp+aquqArH49/kapmd+ByvbB
TUU7pNUiuxlp0Tdi6H08XepL0ftxHXGoVej7B9arfWnghmv9J2N/4KAZwbc67OWpf995HfinEfIv
FU79q6dd7lCSM9LMYiBQLFoEudMFn2ZlefcG53d8ux3TlnMH+UB9JQtPLPRYHaBbsVoCIDM3IR+X
p8tN4I0D+FLQvm/4ZXWZGXpx8Cnn5sWzp/6QLMDdj4M1v/7suPLxBsB6FaX1f3w9RjBl7AIVP/Kw
HP/bQfUut5FoKm3dVOlAI9oMIxnQG2+eXgW+E8sPF/6xxAIg06K+j9fs94ezF6S9O369tkxJOiVl
/dl9apujaa1ItOn50A3vNFYRBg3ocufJGDau97zXQf85jWy9DRHUllgGAfp1vI6Ov87ZF27w+6+p
WJRlqvZ0AlKb74iQ4PlqbOGi8d0ZeNPEsM3XDaVgnnHAZIogWRx4hodIOBP/MlxWvUx2Iz0SnU9d
2EMAd+EYDFmZTd0wI/8kjrBFmRsdeC7i+XhXQ4eMIocQCc4gQQBCGnwpI5LrwZB1lX5JNF0f4u/n
kmVU24Gy7+IyMhnKBZrF78tSbcnJw8drXmt1ZzhWRzXjAYI3avAqUt+phTEa5H80e3PA3IoM9WRY
yWb0EYyRxmE+7rwPraqJwNZ1gNL3jBzhCZhZQANZwfDVw9PbShn91EFFDbu4gQypCVO/Qf+WdCyr
5MCop91wn9C17Jz5YZAufcHjKiwoWfkDSS3QR1fwMxNHz8uEFAKAdcc224FqQ0Nh+Xw3oFqMJYG2
SJHcgrFP02J6+Dd68jOPhOa8jcLP4mweVOw7A6lEh5rX+6Cohx8z3M5xF0ILnAPLAkJnpazxUTT4
HlyYN4h1RIS1hGqt8EHq/BJBsH/0UByfFN8U2p3Vxo0nPgZLUXpDHIqP8CzNYiAT/kOTLzA/GGW6
hZWeJ8+2PXsm42E9kThcvnQmo/HRI2WYqByEIjt14p6adM4ehKCrmFMKW51Wa0LMcQFJSpf2wB9V
RpkZaoXSjh3eSmngsplHYowFfbvCeVBqjpav8vk+2flGipMLIrNGdDsAyVvR1ki5VjtVnXvEE7e7
NTEqWn3OgGHbvhHk/+EFUm1OyLGFr9QV+49GG7TXBReyvHZ5JbOa/2D5MLGP4FApRLdOx9z9Ctol
P2L+9R1rFlRLelPHX5nz/n5x/7TbV4ATNGsBn7E2UXRKy8xAKZz6codgf2wU/Mz2vPBhwy809lFv
ZL5DrLoWd3vbjPJEEJykFrkiVOgzKhxdEmDwlgZ7/wTAe5j6jo1QUCmOFuss/6eVDUy6WlPyiVG/
HIomLPZqA6Gy8KsbbAXRHUPmCXcAOHIIiWKiFKYwvXnJVftyx0cMzhzwFKYWSWEfIZueOYqOz4UL
J4JVtzfG/yUOYwvPBsznloQmOj8+nrtxAolzykxFS9rAhJD+bFxuN70YT7AasYHe+iE20VYb+qi0
SycgSh/5H1YbklfbEocujeQjqv8gSkJk9v/u4cszi9uZ6TsuRri9Ea8xMcUjjmCoh7kTeIvbkO5w
i4e9xGf/JhpuUc5d+5chAQrjedCSmOUiM1wS7uDNk8Ktn4VuLJD3PEZIYnChoIPSBMUgkianBrrQ
oQmZ9WFuByc9e3hVflWjCK9FyNu71/5nHB1LUhGs5F8rWW7yeW/QwKqy3wC/z5kUAUF1YcwjZHON
beVl5zU6yrik79W6bSqfo+VfIoU8yH/EYW9GE0c0CHJyirh96h/L1xftqoGPkizLPw1DNTVADfqD
JGJ/SINqF/mq5qK+ffi2R8NKLgpO1z2FvluW2q8pes6rKGzn8I3d7fbKjFvp9FySEj0mCaCkDGwi
M2aX4sXl77f/afxnvFcwietrNEkZo3bqtMoT2jEdnf5VaHWs/89wR76++PaPVkhZ1GGINBUUZA5e
/iet7iqFAyf74wF58XJUF1f1pVBIvYWilNJMofs/xd41u2epKlBkf2Fya2yTcJJSiNv6PTa0PSFJ
rKwc/RUyFZWNYQiM4N/iCfyVuku/wiai72M8VAbjChX978Phro0JKaSwgW1VR51P5ong6ijo7Xep
wTnx5IHTxY+us0nWEE6kirBBzTcndX3k7zxT3w8C6bOU2OJNqusjwDunn2eDb/7zrMji548sLn3V
HLk7osM1knvrZz6qgeOKSO5tG3PjdFQRE3b6nWYvR+oMwIwb6+BvQWyNINhzliB/qY6mqaqwPklS
8tQ/6yywTOGewigaxdWUFYgR6yIWs4h2PWOedzSYLFWnoouaJEXPLwEIc09g05FgpXVd0LwYlzda
VtUpEPfj/6it6/LKzq1AFnOMdLJjx1fc5qBfS+e1jb3slwVtqLXrOh+5cO5wqj5rhLHNwilRuiDv
BBsP2ejdpaghnf4yrVY6NBu4R71P41Gezn/mjDdI+WEliMc2123fHdpIi0z2tQW29Ksl0IFbIV37
7rovSG2sOCsf1b7nyZ80IUd9R1AVutx16CfBKVj/IuBvIzqAyOKm1y+kuDkBPaz8YJjvx2GoIeZl
AZYqcvzrh6vaDYSAf5Gowa64h3qXW07bomnMP2mG71xQOoHy7NQCR7miIUT3Q61Pntj6dCEoAI4c
mhjjoy1NVCUuws46bxHo0ADuLXmyGDsvWET3XJ56myGS8uOPNvHA2joOStIP+eutNaNL4mHQbLde
F1Hid+AyDR9SxEdL8nEFX767RwD/Ha3C4UgQ+o52hIsqCLGCp2wJ7qxxecLzI7Upsvf6+HKcYGlk
k/eHJFoNBpHEoS82YFp7RMxiIF6TcHEy2Hwvabd/yifPbQKgUqSoIO8YBzWOq6HOCXi1yfpWt60G
OHRYOQiqg+puFplzJrWJWRk+IoiUmCFuvbbf6NeAJeKdu7WImQ9sQevVNf5MyNJiChzGeP624Xix
nx2u9ycbkA4iVe6Scwa6jCKO3nSCIAeTB3Jos3hWa9OjsJyQcG4U70CnAF86+jkSaGdRemRqZP8T
UrYCGTEiOZJ0EF2tu2PvZkJmQLkV+6PTCkBoA3uXaVUs4sSvmpq1gFfU+nF7uvFqWMLkN0Vo4Owt
pr62MXaXjI3blYNJrZrJ7GP3H0uFBTEKpF4M66D3NfaiI13iKxCx27LsmHMoCD6nWeh+ux6Ilbkg
SbRhC0YGWQC/tWHx0L/G9xNVeTsrTKthySAwQpW/WdRnv81ZUuERVrdt01zh8ezvuKe6GPy/lmdY
PYZw2C3X6EohyG7BGZp0TYbllIwFv+uf+YnLCtV3i4MO1q49OTssrFbTgF4jH4e9WLQMajtS8Org
Ba+QhgWFjjKm3ZNHh1+S7CyDXSjQScFA0XMBinLy5qtJI0RN5lR+pHMkSHYf9buUUpxq+a3+BJP6
Mhnq27rQ9JouldC02eBq67fbdkS0wVo92xRhnUoEG2T/qQ3SJFQ68kGo8Ki8xhB3cnjVxmUgYDFo
AnzX6IP7vYv4DzQD9m4yBZjcty/KnIufmH6bR4LNncKlE/J0RrIzRzLa+PZaeANX8E9IMx6QNAm1
KnBx50rrHS/b/53U73dUkt/BlThSZa3Q8TXnisJPekIw79ODBQ/X7WwnR8vEP6vwaVteaeaI1btQ
ps1zWjBSYHT8eV37wzJzuDAW/FSBv21RCL5fW1HajZCEapch4g0n1QKIRRRFOt4FO4+faUrhd3eL
hII3Y7tSzfe+qw++Xrtw/M2GhxvUuP0/pLiC4k4yCnIjqbxfqPp1BNnZNxDrWq7QFCpTf8qCqXcz
bf7wUzzZ/NF4qRff1yrte/XI9x7CTfzVV7iALiYNKw3P+2PxoMK/LZ26sg3R7bxpf9JIFKtIxwo5
5cHgiWSvn9dT7h/x4UxpjRzm3lWy4y1s1c0iGtCJvuZIwpijMp7k+N5vp2Fj990MRrd0+6n3jZ++
MKdG8ifG4R1CSP2bSqLhNGyc2TfLCrPDDVcpsqcPiy40t8vp/XvQbJcKFO29zJ364JKcgrt6cJJ3
2yDD+J3JtFvWQGNqKNOol0VFgczTCZG6q1wZh7yPq4dgLuxpnTY+NZQ7CHl4W3ptKx+nrdt7VFDf
EXsh3ViYtnfVkRTCqXGhmt3QN0kdgVkJSHGpEFE3MgvsCrkQ0pF9eA/P786J2r/tGcYrFDjomUEx
Koei0eNsoQwQJ+NBXFjJOuej525cawsbm9+WHRgBhgtGGMpWVQ30Xk/PHpRU5l8tTRtF2qk1+UCr
/NCTUBom+d5fui/NOX2wNvEAqPlSRI0G72AsUR0yNrz2MjViRMUBLlO9Rnsqy1HkforjKFaxVVz8
8El1RetGQ2eXuFoKb7b9CeswS1UR9sGOlWfDFou7o9XvNV9HFCKg6zNvEV44NOXM5UjWDUUdq0Gm
uK5ZknOs7mw/c71kD7Vd1zeDwegwGo4wcW9cJe9ZB6shQA0xeVFAHsaPFp+olXRPpJSjFaa34ZN1
2TB/gRpz0wd49gM+KOfClB4NbKeGQCy2dR53zeUnHTEKaB735932/Y25+DvRLo+NW32QKPbGXHM5
P5YzkffmM0pJhIx3g1zNRLEmcdv+6TpZaSNLR0PBSYpWxnqQBY0upsNZmMae2Qrcf6TP2NbH/8zr
BsBOmUcW0g1FmQzIimG+2XqAMycrMQUqiHEJUIym5WsZhOPc5q+S77GRzCV1yXRGXGy9+pf4Rr4a
wf6I1aRoYCv1zaXtaglclGSKnEOx8LgFqPVma5PG3nHKDBs8BCGuNKMxRC7qnJ/HqBm7as2NtqTX
Dh9jKCzJr8I2lxFVLLOHwau9q2vzJzVV8+prRQmMe6nE6KFPFUV1KT6mMf2mnyLR4jleY2te7EFV
8Hp70ZfPxBbqJI3b+zTh8T1hZcvXrtPWRdtp+VKUiXQuHxnGLI1c9pRwBwmHN7ON7vqh1AV0iqLj
AYalkmzB1Q5zVZigx+tJUBLVxTqGimUhhjgyxLcQGa1/UnYnR5VB8QQ3EN7VtUez2RklDkOd6bHU
hFEyaRupVMgfCcdc8hNX8Wf0dCt+/oEgL57fHDajab6lcMxBwINROCGuwRyfGUpXiLYZAgvNIzR1
c24rFR3HsCDjUn709IVxiG1IgI4c8ZPJ/1a6kd85dlv62fDl3jhnwdQB2HAeuT1j1MYrOQEZsHtt
Yh1XUGcKdjkiGbrk6akSu1wknteYJ/DZjpd0ibdKYrsK6DQK7q3ACdogxiBazYy+BwZpx5vrdZXJ
JyI97DrixlRa/+py6oPaY63NDhwScriGyH5dQLMf4hVeUhlCkFi/rRZcLlMd5MjhDLHemx/pVeCw
9aeX0cqwj8BJLrMadz0/Yo6nVgIwxqWsAHBhfJP7WHcMQUXiG8qYMipuHPouJ9QeHHN8FzEv4yMI
Vwgx/oF41HQ23gnbJQKXR06tejbc3QvY3t3gDOVIWE4AUBfKoYEEO8kFMV7fGjGUoKFDFMmoKKO4
9IMqJRqnsgCYWjdg2Vzf3wAMBjXUr/adaMf7a0JalDzQ7XUNEcEDAOC3mx2ZqzCvGxqRbxNITkj2
FX8tKrnD/KhziQ+57CgVX/Us4/nBeyNbv5JEt0S1dAoDAbBDIQEXYpUdX7PKdt5ZRo6GmrCsOTfL
Eoddqr+VY9htmzYpcTnefmDGwCVW8+HRiQA7JK0QYQtYet6f7fkhOgLT9Zf/g2Cnl+pmY0aRwefU
JQojbEA0WiyILFT0KqSllS92/x3EP3ajqgRPWMy1/7ps9Ih8C8Rroonfz0jpLkfj5gWR8ftVSonN
Q1k8zyMMMVbFqK28puDwyOahivYEJlHm4r7QRIwd72h96sl6Yl+rUE2wrMv97zz6vYGLmeI9DvhS
KAZizFOD66dAwT0bYOxr03MXm+aK30vQ559ZoScK4stnKNvALrVeiKAMnWQO4KTyhHl4tzRXFYgf
k4X8Do0ZK3VQ9qS3syuzYD5IuVkYarCuCi3YK5gk75Q745cQUuoTDuDr50I+cGRfrL6Jr6GiS10X
VgOy/2iBxq4F0JX5ovs6SqwziCT6EgvZbQGcXCwlDNR7doTJHjwPvypao/LS+eqWNNeT/4TWQrhW
kG51NQ25TlC49vZpLoIRp9CjIH6c4wGviul5RtevuNatW9SCQ/sic/idwedPPQ57iNL8NPm+aiqQ
Sf+B0opfKGYxBRym3s4Ny8F1GzvGxEdFnHZ7hAWALetAZyCXD12snm3w1eSik1wX/CzhUeHsjlD4
wNwNvWw8Dc3ukcX536+AveD4sh9bJnJ7YnI+kvbEl3SDIbqGIDPkUTSNB2EYFHD5TeeiXFP8MMzA
YLQx5gjMMZS4KbfvfAsQXDJ2XSlCw/SAa9NZf+a+N8JdsRtRfpIy0M/IZU9uYXec37y/WdY5JD36
CqSp4TzANnu9WIVI5Wc5PowoN70QVRbQ5kRMq6IMTJ/+ecm/ZBDDIjJ3BeEJVl2O+aT7BpnvCIYH
SiXSx7n+6dzXAudyYA0CGTa9AJDnryUgLuO8r90azUM360/EBUnV6kZF+QR9HSSS0S5X6WYMDRel
AeMbmMnpTNHD4SNcwYfbR43xWHv1E5PlwEYSddhrgZyrMyCOTJVepOMBzIxCVgzAao4RstSmbE+p
Q3c5RJbkHHQ5pvq8FpYCTxDzhJE1w4dkab4H+DpqCDof93aGW0fnIWQaD+548MBxGNA5HftQGsI7
W45H1ejd+7TyMrajV+aKyLW3PDOiMRDbL2fP6aAk5Ad3KBZ/w6e9gxHGyJrRs+Kb77pWrxOjgJi3
c4dA9GJWRD5FUgkEuRjSoA/wtpyjUBUScmYbGF53Ddi/C3FZKxJBTiu7fkKgpQhb80NoibYec6yH
eoxrtj/f4iDgWhIb1ZZRzIPkPpjnWuPnG3Ly+jWQfHX4gkYEby9iRTAQCp6ru46Pb0ODDAvLcfw3
XA0Pnw0+K+/TEzaTpYnjKlyVEgDmE5o937gn3f/1BmefvmNFeimmyRpnklkTdqnffhajsFXRNI1x
bWZVBad5eVTVXqj6qfgjtfr/dRGPnOc4vUMiMsxnQW5/uG8eFPaHiv6mudzPxz+zqY4olVCqcbPY
uISN8doaAl9aep1NU4So0LsxNS1kzff58vhLOpsjATzgMrORRlf8H2CxjKkPgxqG99p1fnvVCVRo
SM9QMu7E5gathwEIvrBIyJWfSpHah6F/V0+lKXM+rTsa30gmhgBteP13Nu2J8KpjM9nPBbHiqEBQ
Xc8vn3qTK/hXzxa6L/rNpcvjjv3STGfbn5JSqKaZ/ZEXdOIc/R2IWop/02wB0jivb9n5RYLvwGzh
IZyK52vM9L41wrm6fY4aKoTuMVtKEzogaB5rsUaKOvdNOVcQ6Eg5JTR50ViLBheSAc6JMEu0J+jH
LmD3cYtonfuvam/F93FLnnl8cm0B8JeCQcESl/ZPbXRZIGqgoAbRtcsmToIL4nVcvKnTqAAHOVi+
zJhGxQ5023kFAie6twME51cDHuunpbq5G73GeG9YSc1z1iOMbArRsGdSI1Ri7QlVQJPOprcTkUUK
B07mlATlEZZfXn7ScHjA6uMhb8iCr8Q4BDANTrSKxxYyKTog9Y+bBpjd8cUMTr/8pFf9Odk1F9hq
YzicHmPvsOzp/9iJDfhXbaLiwyJF1HotQEFLXRB+BHjGgMcXA0cwpAyECd/MnGLzRKwQ+T7bIIdO
De/wuKHyx2rwSZn5c3jhQLJSgdG7m3/M4ovw4+TvaPxKQ6C8YCNOa2RKrGDVNdw5iuk9RrP3vJOz
f3q0/Rme3/xWYnu8fIWCBVdoE+vod42ivIzWi/gLtfgrAPoXLaLgSa70OXOj1DGj3RC5D5XR2xPX
T5Y594el1DgIdiqft9kTOu+D/evnOpZRW6nGeKJHc6bLlSqJfcOmoT/YDPMPVESWAKucCVMIDuIF
YHcO78eZynkt9wJlVY2t1+8YQSqbKNplfcThrXkj9VlSsDz6l3FqoAj6ZcTHRlNQptPVGxdHCLrD
3+B1Y2i31bxbai5Ft2sOM4CtHLnDNIlr8sR4HIAUU0lsaQEicpR4tCSgdZNIS7Uw22eavj0f+eYF
RNhQAZxGcMgih8Iq70UYfwK+cepkowPxBvq/ti9z27ByKqeAKvBRd7OMALdtBy1jVi7xt+vrasYq
1IFXEawpLrfDIlh2FSfK5tsvA+USEIH7WdWMzclXWdKW7X1wa1rSaCaO7OzWxCkqnJCeBi0hOGxo
bTG7f/wUWwwCUKVeAKfIYJC0E2KGQ+juJuRrJSrpOhSQA1opcJFZu9BDWHoQDUt3e46A++mifuFd
ktcTwr05E7ccBOHAiwiiSjK6bo0Y3iOJIrNcYxnMS4F/YYe2B1gY6VC17qkvByhmVmkCpIQ8sSCB
FEqS/zF98gbf/UNsd4hHasbt8e3jKOHQjAAq6eVJd9RKsGz1TvcSmEbwiVLxW3btkPJGTeki2cHZ
YEEBT9h8e1dN7DDN8S0u7JDUYjju1peCKx5wrjz/0PZz/nO1Kou9bFI6Zcv9/XLLP0mlm8PWBj8C
p5MqOc6BwOLpvLMZkAMZQhz8MK4U1HSwqd7zAkKuA8CGtSxavopwDlOlnYeKCiSO12vVpRE39YBJ
ral4KgvV16lLaIOyhgsCMdQHjadAamOuZglFbLXkiUFzcsKzwIlav7ukCp2lcSmU+gQduv/yzFvW
+2bLBrPp2U9zdOHcmz0w5X2x6Qf1djw1P52tj7uKEoxvKaQA44LhhSzCEbmwwcyIz9TYrvaS/2uz
iz2jUm9z3cqlX28yL3gyrm1LsT15OgAJ4hyMqHnqmW29JQWW6qprHSL5WnlBURhiKb6glIErOG8P
ZNuU6t7ijUb2WigDRXvezBF1f+3ZnZ4beFQecfTy1taLWMmuC4/+tx13CprkfHQfo8P/1jrJ9nfU
LlSgiCgvK5Tv+0MFFcX1pL0WWNzHWs9t35RryWbYbMzb7Hny5VVIaYO5pGnVAoM+HtJ0HmGFBkvB
2W52NpkAr+9lWZt88Nne/SBJQ9BA5jAVAGCedVU6LNi0/tSAkT6WcRCzTQMBewAs7zIkqJpovwOJ
2KHGnQKUUjkMzytkkbtIzafPAhDZ9Hfv35ap1vRjIoR/3XtuQ0L5FXAng+w3++30SWlbLjxxbNM2
CokGpSTEkFazUuowTt0beyUmrbfvCuvYCuAkssSws8yESR7sjyI+/kuD1X9hOGpZqDeDLjAFO2xj
1BHiQZhWk/Twumw/sEvIZp7LeekUZOpv/ZVzfLqEYn/OdbSzWzpcPp+EJU/FmFBHC77l5tjpYS5C
rWStGNh7AHLFGMTKC5m6KZGjEagHrZmvR62fdqtMyu+dPSqvffNXKI1BD266A0UPtKM70FzT6RWv
s5UQHLx/KhnNemqVpVvoI1wi82mNX3M/SRFNGP8jfOxoOIEpWuXJwGie8YucwwPmbx1PLIveH0ES
vjVhx+Y2TV943t6iPmmk0Q/ze/t5RVDHpuvvG90T+cg9DbfEjlfkYNunO7KXg2U8NBEVZoSmHWLv
GnqS0vdx6c/jX+AHPABCyajZCWLadcRVLF/sajBiNsOhXyXMwq4mwwe9aSUosV9+YUop8GxSa1W7
7NbGsYh5JPl8aky3Bekfq8iT9o5x5Ivc/xRfY5yp/7xqXKXXgB197z3+jWmauicrFrkoSA9eGaRu
S5Njq4q0Fw/khYpcIvJci2jMxTigfVkXdYdtVqg+fSwbOIwewnXBvBJVj0ayPFNwOnsdnTDa7ez/
fB/Sw8z+VKkXi4oYvMvaabdx+GJtHTpGMqpmJ/6QKoTQlOR1kWrU0i9sbX06TkRmPIZDyjn9Gc4C
DK919hVJ7gKC7Upv0ofvVQoPXFn3elO/xyj1yHLPQPFfh3+AEtg6iBMP5DFd9Z2snhd4HF40XpsQ
g+qBr1Q31PNfmE4nO29FZT9d/wjSnrGML7oUfhmaN2CPzGNMJfr9KioPeE8iUyqM+aQLZRVmBfiq
braPYlOzKqg5+xPOYKyCIqliGoqI6Xvk0e9zX3r/thWwbkejnuhuBWKPPCbFksa89Tnu0ErvpUKv
mQP/FEs/zNVmP/1jToUehPMKi0hQNTFAOx6fpl9hkbaMB5we28+76MOGJ7vpOboxVb4baugshOPf
v3/Q+nLkagJCh50jdACZS+JyjE3JxQOY5C+MQSw3oIbRDuNkkvZMa7sm167YCIyyT06GEEfK9gtJ
KC8wp2ETBYx2sJF1rc+haVXe+imCylykZgA0EJPllfzM29EoRgWcMrlibP68V6f+03/5wXtJ819u
Jv35VfO9iykjZ//RNn72HKd/cVVTlU/XRLU0faOBgENcOP/YLfKnqJNLu9A8YWsxR9FTDaPYj0Rj
KyjHPAZGl3dkXNruJLVSaov82Jbm1ypsS9QEdO87KHg39p4vg65lOYi1ms/Ko+x1z44hLXOYbEh7
xVo7qWNwCyVlmmLmHazeZ1YD2bi6owA9hbKJWNcy4LhuJtBKYMli/9lKY2wVPQDZeIUG30We016Y
Ipp78pyPRKjE5dhpK23/K9mFBDyq+WEdkEfIhiKOgVOq+grS5HI8/R1edhhLIQ8q2PxNYC382jSo
DzbARqWedsQojLhLrQ7h1I4xi9QomH0hUo6qYP03Np/331sRsrEQTXg/fha3ZDQ1wjKOfDQ/p5BN
nuuXEblmzC9EVAGoA9kuULkH2rMs39VCOxRorDP/DhdC8BhaYyiszC+sppvbZTZJJAWIXU47BThF
V8XgguGVxpCASvLX+IetSrezNpP/FDIP4CWgjv+Xinex9Z8y/V0FlOTQfbly96nKPAbnzMksq5D8
J0pj5UYxm3Y9Th90oS4Luyudk2xrBs/MXUXELFfqHQ00GLnODPPGflrmhGByzat/6dGi21ow+RNC
P4VNMt/kMwBvvKQkfJhuVpWHAKEANUSPNT63U68o+zKx4o7cUf/niO/Zq8s53E51IHILPhHE8RvJ
AqcD7aT4xh1/ZHS13O9S+UJurKLRj6q/BNCnYyBn8/7K+pgZmR2x8ResdwnuDEgZZnUAIaqtaeT2
ZSEACniv69o6hdX487K8jekY0hoV42Pn3me1YIxoRZrzEHsfUQYHk9DMOEA7hIRXxykS4z8zC0nt
BibNGS69PrA4aI9k9prKABC2jWWgM6W55ggarVsKR8v92dm48NqvW4o6+CyIhizq/Jteod9AAkTD
6o7YoT+SC8Kpq77CloYU8P1D5lX9zBarZa6ctzwDC9qmHjvOl3/Fn45LhWfVPJOWTdDqRONuIPBO
N3kJGwh4TEauNgHibS50hYNo3G8EofNs5pyF7rA0UQjcNV0Dlv8mQOqQ+2vsGS3D1qvEKWJPlSC5
X0Z5zIVbaEcJUMnDjoivWQsFmwhw7X2erMrKm/wUtnhuhBuXJEskXM4fzOC6b+T23G8ZPQrgEkRS
3wt1ULND7N6HxUFyxHb3ZqBhK9bmdTKL9WJCwELjh3V89459xEc25Ocoy0z7C1o+WB1Wihm5m4NX
AzZrA56bvKtMqC5i32d9M15tgDfUhO30YRTEWeW7YlYQ2y0VkojEfQ9m95BC8Mz3Eg71ELzckdDa
YfrkfCDGeSbb01zfTJe8PP6UQtvw38snfUb6mmisj5ZtbXrKAbd5u4wx0tY8mD9HsbjCE08Mo/xp
A1nfO03dZDbrCFyTDwqs5UkcqghtWhGJNvsLKD8sapfhZO+z6/VIGOAQAkXl+1IYYJlC2eeIBFpJ
cfn2l0tuFNKIM4OT84M+SEKdRSR128l9kFNbaLHOarKcLYCE4p6UaG8JHt2ZufBLO5eoOAsggf6L
yXKHzIBze3cQ2ALrQnQ8lRrkzSlDR7DYcwvEeL+8H5t+cWGszOQxVx2ObwtSG2JhDgeAL37cXLbP
Y6asLrTpnCt1IeZcJnbYpE+5gisumgY2ZOdfwf2W+zthozeEJizMI5swVGWhu2spgtal2g/l44Ny
yNd1c4Yo1x6nVELs/QZI245coVki4FhnARNpjEF+kqyVf7U2aAs7Q2DZ6gYxKUiysNDqvYdn7nsp
5Tfh+bLjANIDoaUBBwdDIZ5p2IbfNqIRGZd6ANcm0ECMc+/CLohWpvQZ8oYO/MYuXmT2sSIxYoYh
doF5io+fW0DofcgiN9gP5djVl+TiseLhxr94NBjFLQlJmZNT9rKoUuYXWJgaPD6wbAiVBFzF3ICx
zg2Hcez9e5OAZnjdCIYAWGJgXUW6y+CSf8HFj0WQsA63r7jCzTotn3ii+3CUHKgRBN6GrHTbeIS8
fHp8dXpN6QPvSQ/M/lN9ktTCORleghgDWa4JyVsEELNYC8skl81aDMQAZToj/iVTNw6OfaEnPtg0
cuQNedxTdAZmga4zqHyY9fatmVVAds0N3EZOsAiExB464HkwdoQakGbdh/9EdSrvhC6cvYjT1UYy
STN/Tj3UpNDvsCdzJWGRSyiu5vyxJTlH+NWUPUq+KktU5p+2tMXQFo1AyIrrD+tFCWGG0RoVcbvs
uCuQzWh2iPKIg40ZEh/QWW7S5bvSrw5MwxdEEwac+7Aam4aoN4/5ba7OEeo1/1aTH1p6WskGDySF
G0zsNrNfIM1hG12R7M7zsER6J5IpMx7hOp4ntmsHuYBCdGB8isWXyblaY7FwSg4TKN6jPLNgyu9d
VB+Lrpjlo2HkTT3dL/Np5j1SaEvGoN3oPzp9MgzFqh2WA3qy5TfQD4NzeosZu8e+7UEtT0uPMjEa
0aCPpBGrSEwesMItQA591brv3ZOUFHY+8+U9vjICfPc6KYt9lejRhxxZ5bvi8XtPEp6pI7wO/asW
YsoiYvxeWsqLcdhSsUaufhX6opj+kVwBIYzV94ZQbqjOj6DrvWJ2lWTGW9J8Mrgp+YEZj8tsjLJC
jhDzX9sNDIKqsABCERmmgE496Q8uRu7oS5TS/Wdw1upEVCMZOKh0NYm0b1xNtVkfGwNB6YSVwr+h
wWFox2a6HN9nLSYB36cV0xAEE22W9OUal7W4bIgvI1QmIDW6O38/tBJljD7uDbscUl985/kr5Ihw
ZLUUHxfdpYJT8EDojJ52zgYsEjCKBcKpzflxPJNHD7UHuses/f1Uewqhi4ca42pPIaQvCQ8rFAFr
PhaS7W7sYI1hIC4F6pRz+2T2Owb/4vGhOuji55mCQ416HiLtywN8yrxh+usVRtA4Pr+weGEB7CUk
fu1UmysV2RjeLjdT1wxuS6scpZZGZEXTTQAG583Ho4TFjB+VUPQ+381dOPSqyue1lMS4e1qBLcW7
GL/7nF0EpcgEsH2urRxhH1zJ2W59rG/IqTDZEmB89c98nIiPuJpLinaQLvcTMTwEICScE175sHFS
FdIOSgMYDz+Fou+hjAgKL2zw8qJbM6VMtu3dgbOwsLbr8ZkOAa8qURX7cWYSizhUAM0cZq6067OQ
KQWbker145xx1ovjiK9lmNCAxHd7GE3PdzPCMXtzdtzkB0nQ3MgCvlsjRiU5xuqFZZsj7vIxYxcZ
GJTvTAQB7oxiI+jNecoPeIfFU4o+uQZxPOPGWan9QeHzhbctN1ZOKzjsdHAiklGbyox6rNxQEK4J
UE5WwwoeIy3rPa/KpOhkVrFAuGfNEwmBY9iCaCywaJYw1EKhYFCTBUNRKAPl3i6nohIjiNqagQTg
gHj53GUwDcrDlvov2BxWYFsKdWFLdOPq3Z0YmNEy+UoSikFqCTBLyta+Af0d9oUl5nZWF8HtCsMR
X023g8sTF/CMpakK7F0I0xSVwVcQ/bjpEceLxQfHSu5e+Z2VJgraxZCllDytjTrrDXQJIEOs1Bvh
DMn0FR/OIYprKLAbTyU1/LQ+D4xvGpp+CDzjY3TJQAb8dc91jR6aQjqmtfyOe+Aj/qmWnO0yrcbd
TC8wTQNsihAhK0HhDFa+o2tJ06c/haQHsTF/zehII4fT/OUdSP2xkTTLwikMpn84AxcNkVxegelM
rWGvpQcka5HwT6JU+KWwiH7661OBXGf8JL3oApn+78TgIbDikOxbGV8S9C5SHautdXRrEob3iE4P
LwlfQm43jVdf110ai8aXaXh8CTa9jcv3NmWuC5z528ECz4XqCyzitMafA8MI1b62LEIVR6KlNyEV
MsMW+i7YtOLQt04tDakHl/onsbAZaWcckGILwBpA62tqckOTdEvvcg/ycp8ickDy1Lx/xoAd4IRp
tAeozG/Be6AxZkRCQ99FP2vbsbezWOSCdn8K+6FsJOaQ1BlJldnDnS7PaLJExm7HLDC65EAtA+Vb
KyTHarc3KF3qbAVSdemRLBC0QT3H5jHY9q3V5nMuurrRrALtRMGxvfTn1WqzklgqnOg//xzujnll
lpmqiKhIsjkzUaEyMTAPmY0XWIff0xLEZMB+aO6iYp7jNed60hr661hn+ioE3qP9QxVnj0Jn4aEe
J8jaxiA9FbG8zfZ1ow11XaBKb9CEZltFiF5+qlaeTg69tec/3RhOnvxr5nc6QBxxyiXX7uXOJ/HQ
JxfNHJJezCUzmD/anBv7j02ez6bUOML+AiI84ZNiEBvjYbRMPMFaMvXNTV4KDcVKsh81tWqITdUi
z/vrvT/EYHuKRII17DbRvD6MUpPTDu0NTERTXDS4LjS+BiQqBaWIKZTj7AzFGSjuXgW1u0Hn1/f9
L6ANLG4qADdeGFruym1AkDlNoxKTQtI70tvG1hdVlbqyXtry+kuK5WPkJ8NMR8jKgL0SCeZlnKlM
gQwgvBPOz7AHBpfJIBbwhLs23zexhc/ULTvPPJJ7KZ+rmFuHn2wosNMnpLlHl27VOUpohsZYhMDz
KO+qxPns+qtCKp8A7ugl7vuA4fr58MbHpUxMgCwKouXCHOTfs+/SipOYqN73QvP3C0xPC3Ju5liu
xoLWyrVhA+CX27lsYkG+VYEyICe5SHriJ2Lj4+s0Urrx3lxppuO4fFx/ZvZRJwd5JSeyrU34rmdQ
2zir3bXESaWDdEKDTvg/PdbWAN9ySmm5GtfqALjLiskgxe5HMC17cfDK0W+sq2pIylnlrfVy/EiV
p/VuyzFRoaQKFiizRwx7hJ3Yehld/oxOaeOA9uq8gb+j8whQuOYaa5URzrlxE3mxdFhbcPsrniqK
TEhiLA7kDOafJZNhii539v29pKK+2oZvARtMP3e+hN/zYtTTh+SKXUPYTR98EL2xlF4BSMHPPedO
5Oe5ZUUVO3tNKQBmiWR6LRffTNvy+cTKJOf9fpx7igQj32fbdsUC81R/pjw/75NmM1UHZCUg8eW0
/fO96msL8GWjeZPRF3P8CApEXl9ttRA33oLyLe6kH89MWx7XM3jYJaABYS4KKgAV9bAcLVB1GWvE
2EK3xCQ3j7/PNaxurLKkWO7B8E9HN2wsK874WpLCHzgcFE1qzljM+UdJdQm7z0T+JhMOXQmdkv2O
UG7iWbuWc0YMW7iQnbrTuEC1OQw7mIjW6a09yJtdPr6R2pmljFEk2meqsB2TqLfjKMrI5KeFqOOD
kljEIja5iJPTkid4B5TestPfdetGUDfmQl2cBSRjZLiYbeb6JHNfoBgWrYHkS3RUN0Cbj7sQa5iD
FFGsjdj/dlfdMEbwIdmEHuyXV61ZifQ124UsLGf1gNAr8F9WrF0KTQ0vKZQDZ0cAP1PUCI2eZSaC
5TdxAD40GULKl9AlUdVhD+UaLFAy12NbYFu8iKcpanABPv3kzGZuOPBBPZUou8tJf66Gphqz1nuL
aH3e0lKNca8aFhPBwfImnAQqSImMcFD3anOlVgutJwQDh7N4LqoZMC/TFgYo8LRYylZS/kt/+Jnw
nrTOItj0YF6XN6ahqw/MEj4opFzCHLC6tkS+Mf5wRqrVzPCC3IpLVzVevbaT2y8eBCoZ6z0q7ENI
C7TH+AGLpwiANLdlr0EcDNP5W4ZTtRY3l1tsCwg80a3h6ICsa1ejWDAlSEJNYYnf7GLj12zfTVQS
hYkg6LIVOSSkUCI53MjBk2JGkaEaB8uIi5qw0fiYWepyaOkQqm+npZ38ZgW/iPZ6rICwj6om0htO
9pTepliF8kmM0UqVv1XnCjGVc3zTAbmk8qmC5PLtiaB+lFbPdkn3V6sZdbwDMe6ZqzEKWHjlv4YH
BbK00Gu2mXX+rRv516aC0ZjAuuObjRjXRaZ93NAXz2WRZbiq+UpOd+W9e2rSyz4kvJ7rPCDlQ2OZ
wy9H8rb8wvJ2lzO6DhA5p2QPl/ARzo6Mwz4wUuNW24tOgKb+IGTsyb20CGiW84UNq1l3RLWzra9b
7C3zBazP49vxhgjK1IO2wijbdkSVyS8VCcY7eF7upU+AgSlGRtYEIEahuulRGe8KddoFe1d08kfk
R6GZ44xub5oo6olwXqHSNGJVLgIYmz9rlu76mQXNaOMK4+bmuCB7VDYwU2GD/VGARawil0FV3lQi
NW1dsVnz7KYoAX87pA+6pbt3ADJWJMxhcD4HYTIqAZHYQH4I3QhfiK8zQJRj5JTLCu8/TtC/2oM4
kM+KI5PiDfBax+CKxYgej2K/S+ve6T2tiHVH/4b02YHz4+e5tx5SQUnO5zsjnwS3TxONTc/Dnlma
cplLQKbNj1at6RwC+N7zFTEwTy3kWm6sEaQ/o9IKjGuRr9bJRe/cf36F4YAq7uJqI2djceAUNwTq
j6SE0zt+JIWPpHkexVyYSpXVQqE94E60HwfzIGb5b4kS3hIBJlyyk7l3TyaRiAq36glRVBeS2P/6
py8sh0EEEtv4+LkCwsOIlPjEMbgGej+CBBQD64chTBmsqRD3OWN/d7mx9XerfpeNP2YIu1a5ZfxB
FuZ0ZbF8emLEAKBKPdeWEO1k4plfDkkc3uz+OPBCTBuHRWs48PFHbixh0WsA4TPbrd7cq0Q8hg16
hoiL6n3kcBObdvOJRxWNZDTgp82CJ4uyhYIlB9ZERwYrpzjYKqsfsR3a/fmO1waoiJ3lTAb6VKl9
ttNOdSN+gsBVNk30wtlkbCoD5fimMM799D6qRqC3Vz97u6ZWb7e/9pzkYtkfE5Dk4CDYMk2NT0V7
LH8Ie3mMev1eE1ODW4FWQSXSnPjmDV9uyPeqbiuYervi8435zbes0TSrVZgUSVarDd2aUfY6AKpQ
OQbWJ7IAgaa3kJwoL3zKykYhD6U/mKTAbopq+TdhHtRmEkUE1suXEI/s2z7fDmVTIoCdh2J62xHJ
WmqU6MnQV7+3ISM5Mlw4iaXj+/UNFWXfoIO9pExlK8lajtza2jGErUuF+mXvYGUoDUmF3BgOppqW
uJfkNK3/O55NVIxgny6ytmPw5OuZrhSEfa6UmvBMRHZcYsGNlJNGESFhG2MCPLUiwULKO4VwCmyj
nz73TCuLhQ/3i8VQ0B+v6NcK2iRX6Bkl6RYcv549jay7UOOnm57Sni/bVjUI64blFE2V5To+caJt
wnMinSgaQ9vEfbOIt3+zfYHU6tAQnuvsYvCA/R2+b8Fmu36VzRnmACoRJHqvUIgxmF5JqGox9WXo
G7NrkGYImm7gpY0IR0vgMqGf3qMQuAk/WysN1mQVz1i7JPZ5g2zG+HwztLjhAY+gq9sLMcn7aIEP
FnOkPFmuBQ4d8NArctxGyfnmBb9+FPEEFm/kh00zxEWrd/1rimYD958bJe6yCq3BvNY1xB+W+yLY
AMPdDPKvT3yHs/2b0j5V+6MdsEta25MDxWhn5R4kNuVqWz8iWICm8c7jWSehDwtCEezxt5ldtaOH
Y+9zRSygKcjmeT6BACUyHjo0bU7ZH2EiELSj/JKrMW9C4evF2Yu7uPJ9GB2KbjJEU4xn9GyX8J7p
yN5QxxT+f48oBsb6pmJS4NUgM0alP9xKUd6UxN5qp9KrlOHOG5eVzxmb3q17XHhhi4PnpfCd8GP3
MJsnfEWe1ZwHuw4VKyJL/YVfUNDDKk8WpkxSmHi5+n/t40Kj5QrEwygBOal19hNqtmJMN0blNHey
0Xvasgu6GIjTl4hsFrM8Neye3dGi0Bfow+KI4E3hyi6RcvAnOD2UKg/+2eqtCV+jcOQdMwI3SrUa
cv5NUmnquYSNGiYkC5dZYBw4oDGvucIbHhgMu7wFMRAVvvM3rbO2/35rtbr5GHsqp6AC2BK9JZwM
gF6ydy4H6am3GUGqvIYExNkHx2U985UPeZhJj/ISuGYM/EVc2eHPXwDIlbLNIieSxqYR8BZzNVL5
B37OrtNji9NHi1oIgLdb3DcLu/haznqcd4po59NgOKwE5WTfuEx83jxevQPCWTgoZ3OU2dbZ1Pew
dUH47xHsGPc9Mm37wKm8FztKlpIgt63Mxz4cDvBXo1IP5qYuePPn0qzEkHSWuJOoxhRIy2+EUGDE
gP2U0FDyZSJomTqM+eD/wTEiwzpWR3iHOSBq3vZ0vqmcO8XSTkG/SiYHhVm5+zJG4TQl99BQnhCM
Ptj5DWsRhkI2kL85xP9sxuHU7qWXamB6IGyv2x+x5eXKAoYna0l9uHKQjoozPbRWeYI32baZtJoG
TQxLdDzQFe/GJikUHDpOwRDXHcJqFhmi+YBAwWJEI/Fw+AxdmUYFmZpwLmrM2bTY8qEmKvpT4NY+
VijwQRmKSq/oc7cxKbCHCwWRq5jQza8rQrEGr/74QLWB35NCM3Q/W2Di8cmzOLTN4BFRZ8GIMWUO
JIGgIKyWBRxuLqbgCdaAgNKBFc05Jjs501ir+ZMe4VDFFzCJzRX1Mwi/MGm/mHnJQRVjCnyjm2Ji
Bo+MWbQHtIZVtQY9hNlJeUnp13zDw5gzeyJ2310aV1t4jdAMUhxBhH4xpAyN03RVrS4PzuiYfyWj
QQ/3ziK/yLO+XbcbMAA8rsCfCRb4UxUHhVHC5le0b2MKhQy3c5sl13PgdrWfBHOZJUVNH7XLix/p
Km8+kzvsS8MUvKhP53lKiCNhv8LXnNGqP+MnPe6D5KlQc7M3rFL5qlimxgD1DADNru0pEBZFyLFP
ExupAoSyARkICLh7eIzbU7cZ01zExOY13aoSXRp8tYKKifc1Hz+VpddrZWAosKv6YVu8f6CdxWnL
VG6ncYqR8uJPdmQQyYa+R0dy9TACJ+cSmVkC2GnRwY6bux+Nc1mpwNcNVfuIeexEEs/YnITUawCh
M4X7vMN8HZ1BUoa1+gMT0Qq+EA2qs6f3wZD17d4EayEY86WLFdy3Gxb/tstpixHKZp+cw6wSiY6k
D6IFqA/tPBPMSGnfWT0Loo+vZulsnWNeZbmJ0W0FwM4oRoYG76iZQdd+Yeq+JBNhMEmtZcPxkO9t
R8KaaXi82NuU1oq+rp3ADgrPcp2lagQyal+MyFL3xL/7Y9BjBVQIVipK7tJfBRlkdSfv9d4OHL/I
WXuHJnAKwMvXQS1Z6wy0cXlAl/yoU3dsIQI24sd1VcoRdSSc/DN0mCKE49M0G/2axXVT/QZOJNub
8Kr6YLrwPY9l8G+PAMgES9fE05Cgy7rnMnlJ1TmVBdpdvQ8loMxz61xx3eaOuv0rSm/zK0pJLYME
CFgeLSwuQIR2eMgs1W+2d5e6NLv3cDB5jfdOx46fH74womjbMO3Eu0pvB03Y4zk/BUAcu1b2it15
ll6SpDjlTjtc6L9BXsRg+wjfuhclAa6oHtZ1o4r8CaDbf27CnHh26zBi/iCn1BZkv4frm+W+2lw+
E1+IGh/Yc69Xv8rSDtXT7xXIS4ZQoQJJSZhXkCMYIEyDaseInEqRfC9/MnYZKt3NmNR7FpXmCRlu
dw+M4NX2dX9f+yj08QQcRcrBwdSmbo76v7ShA3vr6KPPmGB4aYNRPvjMXk3mJ7VNz4E/w1eoJZ2E
nEwJAKuYmHefpSrFtn2iSdfrNK71yDw0/onjhtCrfRmypViMHnNxCdBDuYsw+9fJuznZ0SDTZFlH
6Cy57DOijrVb/vB+SeqIJ9psfHMtttxPUB+1tf0BzAQ4jmzrkvE/xxfendYjXLEXrLxVeOXxAt+6
ie4CAcHgv3eVbbUcYg1L0qpniYov9qb6DvI4EApHf1IRkOvmxpg7mR0KKuWPQDCuQEAhu9bIL3En
Pud0QU+Uy+ybVYVEYvK2EIY+2mQ8obK877FKFvp2vHi4m2WrMrZLq5LPUnnr0lGB2t6YF9nsLGlI
5f/VZIzeyoAnpmPVw1PnfW4gAeic/sZD/h/C4Hz7S6ElW+M+Yts3KVGVABzhQzINdzcXzOzXY7oh
UKwv6zGxE4rsHBCNns3QbPLRJqKW/S8m+CUw5xdvqTGjrAb5x7mtStFjdk0qzgjuznPc/bgsTlkh
oWvH9r6EgYhrMfhIsF/8s0Basuhn6vNYfS2U8Mh7SYvwyPBaFB+qmN6peW01RctFM7oQsexhQN7y
0CjbWaKLR8UANGNzq3PacbLc5MTdVq1DPhGzpA+qK0ClhvIuvLTdqNk64SLEVs0B/QxMa4VYReAX
PXI95EvxdGHYUQ3VNW2kWzbY8xeIjB1m5APFF5HYTATJQFeHGf/ao3a2bVLSGgHFTegPs2LgKLV8
9jd6o6RxJSqjvaBGxcr5p6h7kBxVxAvo9D9P1GVE+vuLazZ4HH7+Yxvbh2vQLBzXHummIDcueklV
44jzpHsSPxG7a41h+XQRWkw5sEn6akqBz0966elf2XE/6zFRWfMSrkmSiq7j/oPL3Uj8fosVmRzM
q64mv3qmMhqM+m8CIa9KxOd4CxOKYkGhrHEjRT9qfRbO6BMOD40RoADkcjyJrdI31ULSMqsPZ1Ml
uXQaT5TlmontJIpzwUFIkGe6ZFkJVjhuPzrs3bqCR5aqhjOm2W4O+fK+lCWHZuqAbUX5oDfA7ZtJ
/uFKFYzOs4oF8RolUrSc+afvFjrW5BmPyTYlJyifhph8DUMsjjRlJN4U1QVg/noV/PbxPGI8Js9w
k60OCe9opZQr68N8PgjThrUxOy2yAaN9P7ImTKbcZL7PTXNWIPWsBBwlHYlmAFtxtEQWe9m43yWu
VopW4rOlWiw7yMqgpRrXETqTJXK/a50x4KUafJ14mr7sh6lUv/Ok4ZQCm20Jnc+t8hYqsVI2MWcb
YN5bIejteb2Gjf+IAXQdXG+PNWIXlKL0DMBq6zdnuM2MLiQi19cah8xHOJcyjdNrsMRUfgP5GgYb
G+yKqNFPwJ4vKLR9cO81q9r48PTxgrPRSkbcdZmpi7CE69FnY2f5LWOJjG9vCmaDiaN0F9DhZ4Mw
L4Ee5FbqXxO1bStHqZYgEXK0mMF22eHb+btDXDUvSgkKZAfgusneGdQswLAqCQt8gknPnQyVD6ln
oDeQ97+wLNXo3qSRlihJmhy9Jebp1D6rbEYQoK7mZa3a8hSGKu+sGeIK3oVwrurnE7RSykWq07C5
cY4F7OW/wX+yiJlpmESzW+uZOfyNvhEGjYpOJuSvqMcBghNAj+awC2D89P9ez8YnIdCP0vdkTfgz
XtodMWZq+ga6xvlDT0IY33wyZU3rXk9G6iUVb877Qz8wBYTw5Xhe0d6k8mXpd0n9iEKZAgeuXJwJ
XgdN4UnGkN0Gy+qBWccRIUUJ+XzY0Gqf0EKZ54tO70awr6HFEv0EwS6Ey2Re/a2z951N00nZSa7H
8hqPOJslF/pU01R8tWuSncBwWKmC73pY0rmfSMIqAyKd6P7kwuXsJdZforIVA77hUyQupY19213W
APrVap/0LT9nh8pWeFbMYPjmgGkI6qVVzy2yq4MoCTdOxRTUDb3aBAdnw87L22LJal8gvWMWnSDp
bKnPJJuekCalWTrd7rvR1IwrXx+XTsWXlQvqUOuWe9OkPu1M98tpY6o+TasNiWKUypaTUHAkl/bF
rVsJQQv/0+dYw+YwZA1rP4QQnG1Zn7zxOJe1ZdF4NBjOn3Frz0A2Jds71Q6fqSaKK1lN1FY7cTSC
VXNQyCeyPFgx81gpaclrWXvo6I3RuaHGA55ZgPVX/YZ4MmPShXKeBQt7tU67pScoGrtJ2JvGWokT
ZyviU1hVow82z7ngvqzSt5TZ77x+0FkhEHpSJIjIgNeKnU0VVCRP7MgdISBmvLN33JlZtiIlkkcl
Zg3wPHeyiHs+FZgRa/rPnHRq0CKfH3a/kVn3bJMqY4Ymt9yWHamDKCEmaKBuQlWls09QX3Mj7ck0
reOVQwbheCeH5QMaMDL0ICEwKx2uph83Uxi6y4mndZYIsDZ2vRqvgqCQz9QEMEi+N2zdTYJha1nx
idnDyx6x9Fc0Sd75ID99AK6uuKvGqCXIrqFceyVigJamYKkhMwS8i0Tlqr6swwF0kFHVANED99bu
w98o3XVl6+BnbT457LNWguU7igRfmz2ON99o/+9A4sqH68k8f4mTtOoL/5U3gwxxl9NwJSlEcje6
qcySBHSy0y4vHirlnbiwYUkkX7dFTCcbbiYnXi0fAOxwsKdzyE8e3n8crYlON0MwxeTFjSByN9ig
PGgF2ekSSPV624goiaD/xWOAdycOpfC8TkNqiElVQL8s15kur4mv+FiPwDWaAL+lcEnRxGvNSwJw
k/duwliSqlrxq5POwv54zvetepxwduio19dHPUJw67dm4ybMg7nGdcw4gKwnwGSJkIJB5qq6eqrZ
3xyVZxGH/kEF3O1KLYH45swjagURwPLzNK74Coy2uk66p6tftSPP45eTvDD6RrAdBOsS0JrrSoUl
uZliWVvUdBZLgN7adXA3soUVKFn6pUJggvU7L0PqT27UKnn1Pa40qlo/Rh8PdGXBlKbGOJZMKT9T
nL23n2q5CI0lGdFz4hl4cWbvYtg62CPpFJwTUJ0viXm08xAKkPdz/fJV33vkUGQUttU96+MPsSE0
nEslDJ9xW1UM8hcMGBqMrPNLxoaLj2FhNBVOJupWHTXP1giLR8zxWFeJ7pgzYuTZ3uRtwKTMxeK4
jtGzOcah8F7s/7emCcxqnQ0FCroikdKzlq/fnz3xiHvZrkHnraTO5cRBjeRggVMm2yxmVCrpUQxr
5Ju+oeu+5KZRX10iMQgsEQiLpgBtLf4cIIwRMKFb1NXuRd76aJwBSuWP9VjWfevLL30uIUDD1Q4Q
1eXIAI1mXmg6L5+fr0cbv7DafGnWkjcPTZISyXYeGd/CTNziTiwIh4OZ0dEQNF2GSMwMDlPFGxy3
VGqfVAexFhO0uMe59Q2bNHOPQkOq7ZVHh7xBgp2ubSMuCfsye5HQPBkeTgCNNBb4+yLVDWy4qnBH
/lq8MEeS/soff66Z6vYmvl/eTmsMwiAuO1U0T8/qrwxJF1aUQq5XguI/mCv9AzbKcl63IH8ieTKG
6G+HeMKmDZx5SwnwS1ELvPtNPAwhCHIiKhknRmVeMIQ13omBaazD0TknjYStmI4HiKh1oX4Q0I3c
0WhCAvGhzr4kW5zUj0QmW8DrDncwC1oO/G0egJqHZmZz4VDiDb+ozE27vKzFM7dY4cSAj9NN2GTW
0V+3wRE3HGYdwg2c2dk1fPWzfD+INdUgYAGhXfjtSTGWfPvDlQwoVtOrmTFQbWjcQe/E4acCMjuI
p35KIONP0JA7gVZ+wNAGzIwXJOc2Mz5vqEoVRVa4inCYu39M1a+sVwuwJqgNL2K/FZnU5wIA36bq
Un5IL7SqrfiZCFXVvSyzOAolTB0gJ6ZqH6/fEA8ZHcLMmvc24psUg4AdSnjso9xIyfPfQjA0MabO
uo4+Y+eee6PJ7JWCdjX4qY0lSGlzkRXIkr/bjxNWBJpF3VeAXcpJFsgY0+HTK8sZJ7Cm13o0cP2p
dzbW6puyTeLVaM0AxNGuB0me9eNtQU6fzyY01vcN/DaV040DVI+H7LLuRk9xUcazRME6ieqlu2xI
hMF3y1WxGX1XwYsiOtHASbbwggcLqdKEl7otlHhFwgxhOAac6p6S8WfZ/4X5i5sIo+I7YS7gY7ho
Ag6ltLOkGVJCwqDqHCcNaEV82dDLpA0cbJh+wwbRe0Z46qdLDowdmxt02LMSROtX6vM96L7A6e/E
b8o4RR5vQsKnw8XJIw+J8nkqQkFtLMwhAbq2HnOdMhEe0cAiQMcf0fUqtUqH4vFdC1PA8q19PNW0
4Lhzqpx9HrFcyD0xOSjifD29hqCGNLvEQiqt2qBdXi/J8/xA+VtOsZ2kPKzHzdQBdVmfcXikPVcm
UleZQJ4hWZ9iZ9HbQmaNyV1dm3JO7gb2nOsN7Kq9xBJeqsjUpQErhsXgXx276dTZvGq8Ev14P5Ec
Jp9lIfsyQLvrbMELZZPUIMT96ftrBr4B5o/q7NsvfubsHeQMGqAoR8WOlWjl8AOL5qwkPdsTRc8G
EyvCgEYRq1njbrLB874wR6fuNr4eLsIZ5XOJM8wiD62ia0YkmuEQrozh8ymIxX+/k1XxJZpC4Jtj
emOBVjtqG4PGfp/k1IdPedkQVEwDSag/+ODmqfaxYWMzFiPXVrv8daXJruOQwDC9Zyz1hPHgKYMe
Ey/s/y16QVjcn51YB8Y8gS8LtDDB9itcX5A4eh2ze+y+mqZCf3YhPv/uE34oGpj/yTHbOU1SVGel
wpvM+LxyOnMHWWmizu/ULUizAuv2tSvh+Pvxa+Zg+SUcsn7dXV1XtdURKluVE3jma6FJ7uuEzR84
u2GMgxDZuY+El7v1whT+3Tkc2UhlGaGwy4Kzk+oJBvC52l+pG4XfKGgzoVjDPp6gLkoy7UxKh5TJ
c62HGbvIzpcGTu9yNag41fabQKPxfolLoJEVX09OreaSvNL82BlKjERxu8gNp0M9NnjoNgbfKlGw
ey4kXx/JqQjN6lmvGyhqXgUeO+8ifDFp2UFfZmoiCm4izxGlxD18tfPAX5L7Vy5twdznHhLd96gm
yfKLR0jWRu+RVOH/P++YaLNTzBbzRJ9/tv/W1uLVq/FGQBHdd92wKXgOueiDudvVNTzuh+bOL8PS
J08U1Pcc+wQeOyBYyk3TreUlbzhysphfBsGqexSFrI1dY/04/9AHIf7ao/1HfKAndfZo6R33m5TV
hVEb2Zy2hbtZt/fNGOy96xNnBTQ9BbQt9Gabl/pHAUTX4o/plEOg3l0BuLN33qbQ25WXLtft4ORZ
VQcGGZQa4RZGQAE4qbFY31lie7p8dR6ptNo1o0McKyZ/hAOAF6nuRp3vJA83b5xB3Bog1O9un2TU
KEHYNX/N6Pa+l8eKi/YGAjRnZkh5q4/1SSWPoneBRw04+3eNX5uXDPLebi6gAqFsnHGy68ayQLGz
XucbdjFN82o/fKKBfNUOjoPLaTWuUUm00QYeF7Tf+f2fx6eQXo43ION424uDNM34ndBm4hR0Ck1+
Xjp0WB92+vCEO91BDOXCkbZux7Vl3XRk9p5icyjRUzctvbs5DBpKgiTLkkAnPk6B47ZTlc2UmWl/
UrR8HjTmvQzCEV8TfLbd8rZkD4XvJRNSb/0qrLHjoBPKLgZJIEAC87wQpALU7d4y5q5z5ZGZfTvD
w+dXCfSMBACoEcpHx6GOAMaG5v1AUGEvPJ1gSi6EP/0xUjlxWMLcCVF5D2LnefFYUsT6Jhe/HGbw
VVElnPhTpLPo1Y6uX8I52A/w6Tost8OUIUBX53GBNNqhGUMX8QoO44nriCoU17wWc51QAxaHWRBE
Qjgcr2j+s9NfTYXtVSm0vlkYzZmZhYXszdpD0kuU05k0EIdjd+emjW6ScsiNvhBKENlkIbweRWsG
3dO0Ek2o1MLwI3CValNIEZtIo/yRYtC8nzEhsCtPtvvcR2gtfnrMGmnah/kxY9jqkJPH/qw9wlan
VK85lTgpBbAC81L+eCQTh8qIUfK4Xh5Vya17Pk+a2o35VA2YNUg8HaVIW1/E4SduEVJg2wXQuRaY
f23ckAXCL3ouqjH2A7QbsKQfva874IO06Crwszqbog4djVzrc7SDNmDVImst06Fwv9JBbUWMNZWI
Jp/LHWpXHEfmPXCNZnt1KDWnsd5a6JVvLvFb8b04V9WIKM1n4Y0ULQxeiTUTJvut0fhS/saDE++d
I1csRYnYdyM8k2vBf1F0Kvgt5g0EFG5yNMLHWaIBn3SNWV/4ULtoR4JS1tPKX/wEGB5g42R7pTA5
typCPCGwXJBG7UAM9rLJ5eRJmVLL/4jEAJDhGO7HSwOcX7W/vJf86t2YjQaRpA00usKMzZD4i985
oVgQa0UUbPtHUVFPHxLl84Dowo03nOtnMy81FObUDalNS/KdUtoJwSmhBI8Dc9OiR8lSHzX5ZnM2
afJEtdZzvUBb9Wd1DJI8l8froLsjXa0rvCHW1yTnWxcLaUXgRj35JvqjZSzxY09lYkuilbNsb+Q7
Zot3TEicUUEosVpJYxHDLJS4ayRGyPnpCwFioHyg8POKCJSV4C2Lg9Dm3HL29uKGda+8qGCcLohC
SR5wdlK9f8XuamdNiM/JJXp5pV1foUgZdBcqcas4VUSSIpTX57ygbAjjp6i/KCDdxRcM8/b0omgM
xmRcgZKk/DnP75YwR47rWJhzgt38vPk6zzBQ6Zk7zOmACrvAno03YNglcDubaz0QVln2RLfWKc3E
kge73vp2cKU5jh4XFlReev99aNnq8/DRgQYw/k2wD5OSQ4Q7jN4FxjYx9xAxvo/U6FRF2x48jaVW
5T5/Nrv2pSR3PbosT5gG5Im/IsPBTVxbwmKGUmAubjWWIFNjli+XGo6+kiI1SX6WGHCfaQrYBSKl
wrHZXzw7sAW5cRQEpYrwzaXoBFWhY30BNhU01ADGAkxl8e0DbiVeDD08g9JfQLfSYuv+Z+JGq1uo
x2S/Sd+7fRdO0OFWJROqZ1lqA+UiX2SVwBlnaDWh01cJ8FmopLts/VAjS8ZLuDEn3wp8vxI0JjMg
tLpJYRuW1DoOywLL8wfH4vMdOxW8WqWlCYckrYYPlNWQPL5laqvmpWRT34OSQ2HvyJYQpXovqY4E
MwW5iLZLqjxO4yJzGYnij/fftEAXjVIkD9DjWSyuxUN9/P6IiSGeERyvSNs72gGoMJkqTalX2INz
YiZiVtQibxh6RR121ZHVIFUym3BbR9WlBF2KCV8Z4Ha0qSg2KTithbdn6I37/1blvzHs0rUQuX04
w15X1cTVXhLBEpCogbzqqcoJ/FCk12jwHIJK3C75UxX/q41P2nLMKmX1Im7ljyGzYduOfvtWAEjE
mRbINv2pcP+oor5i2vPIf6a56Y+QsmIrdb8luAhBmIQTmC9FD43LV4+FGyG029bbsYcy5SJNb00C
DKWy+A81PxVTVm7q0Rov03kfVsRR+4KiC2VpxKcJyPtYIkgXY05aFRTnt9Hf+b2+nTHDU21Tvq0E
SYoqL8yLQfq0iU5ws9Eky/88WCodrAo1u8KPuIZSW3D3W++v52pqi91dltv2j0z1Z/WQzzOx2ROH
6ZkzdwX93uOQ3DrThSp0loCw419SOIDeC/sDOuHdwwQTI1jpOnyuGpYjqDJPc1ut7rrvesONvn7X
QnSCRSxhOdFPc/yOeBtG6Wl1WG5dqIZbsAwFtZhuzFjftupKjZwGxzomaIJwxAt5ptG59eQCFHsT
nBL5ad7udSx5IURRaUPVUA7oHbWzl5SAWKIaSNRdQnItj0TKaTaiaVPSfoMRcVEm2gl2HvWL3Xn2
ig1ot+Wg+tASxc3Yf/hdLp3Gjr6B3SE5vteDdiAb4Sfv9Ju7Am48unQyPFgUYuaFpQpdHoJTgR+k
R4J4tEi4f9XOqDfrRAWORMABshTjND5mwh/h49cJvJgHssPEyxtQKMDdEsUVeY0eMT0OSBDRzs1G
6PULBMXtsLVg9l84xC1vpe8mlx1LyJ2kOF55emn+Y03Z71EmSoU5wBMKDIVJEO98XSRFiKUijS5p
jxsC05QlSOnaX2MN0RM5npzzfwv1uY3d4CFKkwYRH/b2IOjely3luyzx9EVrprCl+0AgthjhGSFa
Crdq0I6u9r8E7epHYmw03ThgZ2SvFANL+J6W1dsaQ9r/Xf22jA9M6kAEgN33ObCn4w7tgWa4A/Ia
nAG6yw3R4+CBXThL2JKtStUyRxh/EzIgMAW6UxLp9tP2EAiRbLLsHQ+3nFVLjkRNMoNgIAjyjY0j
eFT69NrPbLq2X+RoqR+O3OGzaJJpUv0omVj/y1lrKY/LiG9vZ96aetMQxEu92NuZoK4vCv7iJxtl
A4RPI3aHiucMJPHjpBmjp0C0FARa5Tw4jr7jiTA3uvSBzw4MJCcIn6S8CiqaU5NVYMHeN4waf9Gs
iaNQFkQ2wZyqi7t+G+f+GNCRJ3YnYd4A35gUKtu2rodQq5agAn7gsq4vt/dGHkowaqbpQpMpozHz
3XV5HdkY40IovGhknYiJTcZT4BGpZslRWKOZkeNKRPtaIFRgSKE+ymrMMQ9y0btCX77lj2cjWZmk
Y5ibNm//xIjy5OR30jWpOiJL69KTyrzwTYzNRrYI1UkX52U+R8GcZwqAlElDOb1+FJG7P9bHqTT8
hCnlk3zA6um20ULrcJzPYmllxKuitIAVHtTw/s6RFJuooi/wcNfZUPLLP2Bb50YU81lEHWFYZvut
f9HhgSd0RrfKbaHE5UNhjHUwc71o9NLY1wCjsWEy8Otd8+wS/w+yifH5GU/G4gRjYWE/xJpQcuso
yEqjhcZd+vNCqwXhwnYKBpAsRgvAineL8rIhseawdj7a9jvHzxEi8eLAjvWPfA4GiXKW5GYeheGd
YykTptagOBsKHf2f4gjuD0/VE+s+7E+v0d8yFhgahsLolb8y6TTZXMPJARs8/IJK0nuaT3yCgRmq
OQ5zx3CLUxnFwrAmE8i/2g/miZ6FaBNZ6OUsQ1QykDnt6TgaLn8DNyoP5Q+Fg5TpteGlRbOlNLD6
0AzrlQ9oKijpHFFzVkXW1PhXt8D3FwVVXZ6nmopMj/trqwFhONIrE64txOms36NqkUjOBCUP0rxx
3vq24qYTssePA/4W2Kary4LPXCWrKEbMJPVEXI7AhJFZ0Du9rCXjdWhURUkPIOOqdp6GKBfYcM9m
1o6hiqKb3OaCg8zoWQ3ElWBViRSF7TmmnuspLzs5RZ6e4Wo9X7u8TlJxJwwtSUoi1NY6N3Ec5J+a
UjzWAB0N+Ne3qbihzr/yZHO4UU9qBRusaPoKrOVZSMH7BHuimgZruDCanCAKHXg+DLX7egZxNf0O
rG/haWgNPNls1wTp0K+HAVof3RhuL87PMfnC69kL6yFVheEBEGhmLNjOqjP2z288knjz8TTI4H9u
Z0LnmnkT/HuvVYUjc+8IGlP0jKVLEem/+N+wdT3ZLt1UUPHK+xPsjBhIbXLLwW1XsmqvTGvYzzEA
xiwrTF4rL7mLD2YvKUsKzjRqfzcw1Syc2P3od149YM5v04ZGgzCkoiKBPtO6dlleEAFX9yK+MlrW
F/F6CuBhwaG6UtM3JEClagHPTYh3PDntR+vmEKBrWqC1FtKnnlQAx1gS1IbySTuiSnZtNEtFQinR
WrALpzr5VUwC7Pw1fTqDVAVWYr+9T7TvAPr4kIy6AxrlCrcqEiStp+jMI53rab3L4aMzAmp8M3un
R1iu3UNszd9c89L03rRl0HC5lghAvrKmz+k19OG45TFA/OlWpeFyeDtJAUaJOw5v6kLJBZmvDUdc
P0g8GiZp13K8JT30Gap3JX4xaWgA3eDyDVD18pOx4ZGzcq4Q+YF1hygfScYRg6UdTYAavi1k62iL
AGq6yvybJ3mxsqLqYlhy9Mg4KXw0x/YLQzh4qfR9XBh23AgMfHPtLjeVlwBfpd46j1mCkU2F5lUk
xPETgVv65Ip7/vX4lRWbmxauKnOrsMpjIfyblQLIYrKw2noIYh2kmVmMSBMcjHLJ9DHiafc/Kkl7
w8eDRT9/+vYc9VTX1DBUpAuHTpdAABJXTszV1JyEr4NKi4nWKHQTzRtXqwMfvtXuZlQGgtmg7cRH
9W0Nras+SVOnM2zh+TX+jzzQZ1oTVtfSubMa4wZyM7nWUsolLqPqNhOWPRlV3z19mxEf6KvaYHHG
QzsNDqv7FAPMBIBwid6VMUazmB67ePd02En2RxqxBvt8mHaN5AXoICvRX6Tc9j9C2ctQJZr8Y6uO
g6gS4p982tfx8F1rkFruxUMpuqZwq5Ylgp/Mvzy/HgiQGMyKL4JQdVPzsiuSHedwDrgTrT2XAAhP
Trm6EM248p5MXErNPbwyCqrAdAVjcTe1VnBRzi2lL020R18JPlB8qoN623bqmwgpCzfN3yj9dMQi
EAxjyCCAxpG/u6FuY3IeaPaeq7q9gl3/8gI4mhzvbuP8FtcgKpTdhvNWu6icoBdxbx/hQSLfBNYI
+8A7I3v92doXjayNP7VzXqb39soxO2trmTFow6fYDseLLW/nsVsQvMrv2O01WluEGd/dxtbnvky1
472pYjsgcYroWIYujdQ1w9Yb+m+N6H+sxIbi37WEcmOCN/3O96V6eOluX24AxdrkjRXqM0rqCACq
N6IIpkTuvyabO9Bh2bfjO0twFJzBQWioGmmcaoJNNVIJNUvGvBtzlLXeMxDhzNGuepV1VGBKlYwX
Q7Ke4dpxCiZGwkbvn50en6jib9ypt9vOQ3LI91c6Kc/uh6bkmaghC+IIxBR6hrj8vThIULcvk6/3
DQgF4xj4WwbPDPqHR5TFY9IIjrUgcuu31238A1gdx2Gh8cGVF5UN5rajeIM23WTEqYfEIwmuMUKk
TlxrNFIjL+C392Oe7WySNv5Vm7hi5k5f5ceybN++yUBapkcD8lxeL7nJXkS3FInAN5hLCbJr4O6P
YSs2zm0VBgDlJVZd+W45LXYaj+QYxP5x2hu6nBubMlcUU5mwtpXnG27BrVonXZ1j0R/Nt5v4ZCIr
+GCnttUs3Avovb9ukXIPWc94jhKG8WI+XcZCb2NpTQ1fFD7HoMCJts4wkfqw7exVjeEruZgY/HEh
5bZVUmnHbEyClI4mbBtOCZlx7rMO/A9M1RvFF1u4FdE/DvoICDVsEJXLnH3pZRUcA8WUD13Aqv0H
RxOwtrZf0/091HgRxcbRdqN1fg+02X41b4s4D5gUfcrKCJ+X89UdcoYph96q80M75xi+I/YBSWOc
7giFloI91sKHpGMbt86z75mw9J1em4j8AwBa8uHJbux3lmmFDyebJ3w+mQzMsnBDK7/XpQHGTbvE
hvCYbmwoDlKu3HwzmBsd5a+OOc8b6xkQM+tKZ5mBLOFWg74vsoW/2B6uGzmmpZqPyVzjrrilVer5
2WL3JEReMslh8+MXZQVCQjczMbae8cISuzqLGR/b3D/9TwNgzT6ci6ny9BvyrM15xzdIZgMiCJjC
lbn8W4Er6gaLhpD4Hpsz5SuzXNelQjGPxyoGmzqppSLInBlO3miQe2TMa2Wmdx4JlAyOWQNfCHMs
fdc8ro4QV7MNHjKGC6YIamqoSD08l4VVl63gaWlrACNOwS7qa1Pa4iIWNkjF1fr+6N1vzLhwJszN
DOTjJmfPSNo1NzqF3B7flQTebWo7RyZHEhwDsdz8VsrYkyPz1vlpwRoWdXzRt18B04LDtpD6qBAs
tGf+E8dFE2DnBs876x0oyS5OURpFQAMYyrh2ZISipOhDgBLonnr7AnLxhFQBWH8hO+NsX6AV4gXi
KlBcVOYV5rd77JhGXKJJ/eP1kWKycAu7GYS6sz8CJ4Wf6z918eB4nrk4srb6sreevU3LyeLyUfOf
XK0Lte9/BNdDSG6FJ5OKPkZNz7xiyOrSK3A0h0IY69zEmkSva3OX/HYKeFjfPKi0NapFlvAJY3b9
wQRRRPRrmidqvqvqLtgCKaHEuRPRN5QbeLELCaII5x70EbXIiYszFMIQx2zcHYvRpoo20b2keu+N
yTjCpQp9auYIfvRktddjZZdeMAtineqIaDy+dWbcO9HLE9z3DuP4ISW+tUaxHlvUZ9DLtKg0NGMl
oRB1eoiByOh9JlHp2nMdaR2StsBag6uDrg40NkdlqFXk59eHWbgQHEi3TLzE9zadsLI5pyQa6N7q
V4wSNdVggZrlILhRVBhIVOJA7STmzn3pSYUqGNTOI0Tz1s8gpFOf1vsQpnOwbUsXQYxC65E1EViB
paiD1KVMVcV1fYjEYDMB2V/gRGClNQP/e5YbYAQjdDooCXk/35CrkbxYW3LLjZsLYeHtVqKiHMNB
nK7Y9L8GigJ0penPfi9zciiCgzM/gXfhO+qrztdpkOBoqu3DXENHptPLGv4brG3q+mKbKkKOzjbk
Drey6FmPA8eURwfl0x/MBIOf8yEB3nNZDGLdZI1sGhmY64yFGP08A7TT0bLDToRQ8KcnZLAS6oOz
6JELmnwzZr19gucq8i6GbwY0bQ7ZrPumTKE3rC5nEc13r65/dXSF4av98IfVZCPJ65wLgZkX8RM9
1T+5tifIyHMHEPyFRSthvj0hQA2E0ZdWlj+cE/2DBbebFWqi9Bf+aPMo5AVbmH6RqdHUg7EsTe05
a5+AQDd9cMSjF3wQEteKr2VNJNhb2fFp4o+jCW+n5vcmHPdus3TWXUZdiw6jtImcrzzo9kh1JSZG
QCvLjF2G5i9qdinhzXghSd7s7W5ogpqF4bGlndF27NdFCOdHvOEchTLkT2JhFAiExUP9CKcVAyyt
887FaT8Xrjffx3AWoMzgwlW1dX/6bt+3jjLnTZMB5LP5m1yt9MO07AKNQQdTrep8+F2u6gRX3soZ
/2iNmsGjzZbO7rvBtjhJlt7vbIkkDV9g6y3crQ2DDGVMo0XDMuH4bDdBp+jP/SoCIrCimw7+hJZM
ASD2TFga8nmL3nwf1SNzvxEwRF6MlNIL5pQ7uu10MYD1VvE7MtULaJul5qgf5MVVkLxd2AXR0XCO
xsIfAhmGX2Bz0AaRCU3dzUkBQ9UjjEdRuaF6y2u+KqMT6wCP40Uru509WHOk4x6fWDxIrP7wgOgw
DW0xX5b3Ia3upCPKf/ZFA0SdDAikNLJpfES6RYKCe6h8A2R/Ho7EPTRzHPdOrlkOpIK9agMqUpkx
rszLxK74YtEWi6zRrT7jL+iMh38bOaU9uPLCOBXBtzgfztooZ9XK8fImNkvBIZoYWxvQj6pcPG4h
1WNLZcPRzr9lbMiqNIgC6EiWi/YXXrOZwXjA2Uzr4umTChkfeRXKm2MWytA/ZSPJT55zfQXHCh3T
V9zii9sUE8uMMFbKHOVKThKbsH4yre53qb6KtySfFR3kUqto//3raYmB2yOcFRFrQJ05c++bQa7x
5NUsROFn8EgD7Lp8WCXhfoU1OwpnoOKPEM/mgC77MdmVCl/6R8t2EReq18xQZXq0HHcdbWS2OsyM
ybzMFCv7bkwzPeyMuu1sBoyUPXwnYfGMa0qmW48YoPx2rLS+BT3/W1ktBTRTr7FA13Gv/FWcy+rm
fEHzz/+Gf+7H1nvLzYgxY9/bnD6jM6zTm3DsnVVbsOXBj0yfZ97YLV6JhY8fWT0MGGjsiBV/0yn7
IxMlF00YidAUuCoR1yimXWC44XbunjmlYPJtTSOo/Vh2RopzJhUbADlk5+pjW+XsRwCRM8gXgn15
ZLEjPr8JEv/BKTKJp3+sk5MR3rEk7NSGzZLZNzyUG9zerMKR+sCAf3z9G3juFu7E0SN16GB9Fs5b
pJwS+On5Jb6cTcukrxzSz2qk3xk7YzLKAywEkaOR2VS8eX+bDsZMuctQIMqZUnqRfrnrbzJqvpQn
8lTQ1Yb5gaw8y+Gip9HR3UCPN1fiyUdaWFAKfzpwTATgBrggn9ZtTb/G7phOyJ+Hv3FVMjroxS4m
aRL1fRtwOqL/lw3SdDhhwwaOyo0Dt4E2R1Gdph03pLB2xJVHficFqrXStjSz8pvF5QRAvoSSH26y
aEWnad0Ijy0aEEsBM4M9p3rkUF33Z3OSQ1w/aHhkzJGz0EUd5lIp0jjV6k9xoY/cJsB4fMVcjt/D
YryPRKHlqvNOn6XRgBkTtoKMgNMdoaGRPRips7EhMk7ZpqxOxN6yMqzRMWMp8NYUlgbXoL60Yri/
vQhX8IO15dt10k8F+HqCoWXlNAlTRQQTrO/WzfcaqDmbBojV0DnhQkdmogi2Wg8G5ZEVGONtDHy/
LbzX/dzAeJLLKNk1X5ZpA3oplcDxc4yYLH4HE8g5dq8LvFwiNAYmpmfVnsmdJ11WcPVq06t8r4z7
+cuTMbVUFo9neA1nQmvC53Le65G0GQ2ZJTtg9y7aTHJIFA7B10IBrbMcWTyx+st101pIP8vz8WZ9
wi/nd9g3ekIm9PFH+gX5DNKwbyRSNKc99vYTOBAdRS8Cv3EW8OXJvJNuMuYZmqt9d793lOZmydUC
EidffrmVuIp97z/f2cB22Djcc+13uMLwsR5OI+gIhRJYoIuiAijshvjRevW9kfPf2vSzJPIS7IWK
LVO68NIvA2CmfueymBaERfR/T0I0Z4vrEFmCAQK/OwFumQTXU9MdkcjPxggSKLsognvW/gs+I9SL
OUwCgnoIE7o9Uysle5weCTvLPnqDniwaEO43+D7EbgZagIb5eccKvLnS2s6YDU/gJ7/p09r3hz+R
zvgYQLUYTfOTQoceICVvMB1mKDJniDkEyWigfWMWP4rPg+oK/HpE+BLAB/pzZXbOBmCFzf2RM06Y
B5ZXPgAGoTgdToACzre6iGr3kYrDOdNu1Vd48Oeb3IrQRJMmutoLGvmXdE5WgGIYsMFZGr6dJCmQ
0/YSVBZs4O/BbyNdy/7+GHDBEH/V/HSyo04a9jWNVNx5RV1EPyIhWntj/dlazQRRKlhimMJG59sx
Yb3TIyEnl5KcSNKy4CUEXg5F4s44vHVF/WjN3uqlMytdArLzV+TcZsAR9XhhDBGdR37+aYdIvxzK
mllP4KcwEhwW2KeusOgLimeyvx2R2ssrXV8kNxx1afybyz5E9E0wgwnm0wYF+aLSlgE204wmVVgz
W0fjCtjXDi9/pNxA+qvSGYvIN/hJeibSbuBIpqqTgk0Ja45OBJP6GjAt1f5cB4bpVGB4FzBBBH3x
moNwCltwY9vqf3aB5ZiYbOcNPn87B/rauYMLJMv8Xyqvvv8K62aAcUcBkcqZzhIYdjFVjIR8EN4t
5oWi7O7sYDZRyz6AHKA5IpLS0m3+LoMRisE4sv9nUpvp22pxlEgI5E3VCtJk3Py0GykflixaQTGO
0cxfefvF+NR3GD2VysquiMEidmzBs6I7cN8accgautU8svT67FPRb6F5TLtwpeODuhOcUjQXsome
GodcBgwr9ydZfFZkCmRfkG+4ymttKv/Yc4d2H4a1oemMDyUp64xYnWm9BYF2tNZjIqPlpvW+AL2u
/5s3o/HAplIT+1KJ6DsmS2+YD7tJJbE1d6hRPYn80Icf46jw9M+cLpWNJzn2sxkLVsg/wl+MYsYc
I88Q3FlEwYeRGnofxRgmjYbx1/+ujPe32MvIc4AXw+EGbnwr6Gy7Q7tVaqj5aBRXwyCMdQioTQGW
DmR//B4t/wihiGmhwooT4dp7VNPOxrKCQxh4h8oZ/KzxWhGMR8A1umx8ytUXgAxsPB4stXT3nbRi
eOM5i39IkV5vJZjfKCuyfIh6ZYIwK0HzUxFye2MaUTz3EtO2KVwBJ8hzEwqopypfRB042IgqerU5
tVe1yVO1B0cJDDb6Zb2wKvS6IhctjhnYDJvUX1ahGvMKtWPigf/TzNisJDZbuEV8NjcLt4oAEsYP
oCkNV+pHn2eCS/YcTsIekXTZHMmqboLqqAwaUJm0z7sDS6AHcxR1yhFp0GpoUytAAz8/Mrauv7vW
ZNHP/3zhWKjD/QoeKrKHwKTJ1lR1Xr+uG5P092hcVwZOH/aGVJlG91uXA8Ciy6pJzxix/eWZG3At
xKvji97rbxuVYq56ztmCJ+asmAWG2O+2Wu9e0zLsoFGpayZHaJly/vCrqGor5sA7/K6DKTOKzY34
ymPFfcjGyjxJ0sOQ+eRyPF2IFMoegdOs39xpcFOU/gus3w+dEUZ9mCKBulbYUMuv06OV/+6xLcha
s2/McBhn+uMaur8Rxzbx1WkBXhwgsPOAZIkj3uSggsHZVhDt/JBKVAMBDUx5jSNncrFgDvcAmxl3
44zVFfwbfLrUrUTH/6V6CpliarfIRcmoBN1IFIMa+YQ8pKic5lPddCrNXao6PRXRFhwVd8mDl5wb
kau7N5FCe4vHgyygIEAvzcc6R7KNM7Ld/j0iyQiZTOTY/jYliTTTL/JkjWzfmiR89Go01voRumSv
MhT2pLN+eUwxUhlHOCXgnmJlvlRKECx0YP93blPfjUATB5G8Ju6czjeOTporlDl+iCX5qbcn7OuJ
0Rv6p2ADmrGCbKfbrugu+/6ou7IyVUG5G3odeKacKQhS2kN01OBPKHNTl1JSefB0G7alxC5sGN8C
w02LzzbgQ03M1mgq5ND1Mu2QtRvhLh1u/yiHFfoQZs/YzPLDgNDf+bBGDqREh6vekSv5HeDS1NwJ
/6W8bc/tj6rjHHTa/uqjd+6mWmXD823S7dO08cld+ahYtj4TsNKyQmJj4jgvrWw8RBx3X0XSIl9x
rJ4RHtsBBu5kI+bSpbjjm5CdsaJvHzUnnjidHwqLJ/U4oQQ4zXiyxmesJsX2MvId3Io9B6acMwl0
AMeIiVDEk8GqBlXpOwW6gUNcStjtYj9loxonNY/j9lOQcJJSPfd+6tTeVKa0oIa6ySRL0MFLOQ5w
gDJf9n8zck7RrwNBfTuGMA0+Zag+PVMDcH909BxWjrbZgITA13ymXIm8GKBH7yjEa58kflx0VMF0
tXEfORCmYG0lW6EzqFIe28F1VrTQmeBPdWqu4vX47E/gpPwkExHVqGdjwb+PxZ6a/XG/st+s3TbZ
KK5R7UBW0mAE9yFWJDlSkruzoW85evnRRZPl7Dun7SbfULKemBB7oW8VwR+PS9BkU5KjoRkFI//g
wBcrUNujDSjLJ/0x1WCTr9W8pddkxjs9rk/9EgmEYjmB30yoWbvlDmxcLPOVcyo2w0gO+Bg+D7JD
/LSUt1GgWB9wZbcpPrXAn/iOqir4cwSyMpu2Pn7nFMQ/GE0AHms8NHyyyzrFPeGcJZBUwdjcops3
lCR0SEGlCfXUIoKRBPyfrhD02aL/l3aunT64p07RPihqVwzA1MinOEQ9t+ZFiXXCEI4D9R0vUDp4
8aPk/wzbRqb4U9ZdiEGiMpKBbsanm8G8eKZ/HqiSw9mXT5fyWLE02gABsQ4zByy78JeiNMM0kPkA
5vbds5bgsPIOyRChmB2kEAa0jl4IcqlJ7uMcjtTvoe8p6qqxLHTIAXL6tHPI3OIEeqGFRDjBlWu+
CRh0W/UgWbLjdEFz6HCov8jLi7Xo/DbMHiIr7feynUGwsUpgFxGflDAqY8NHotv6o3Pm1586aCIe
z024h7N2cmsUJNoUhnW+LJlZBq2CuSn1sB5x10IvU/o1caJ8FHsbweOb/qzpIktZDXclw7xaOZrE
Eq7GEUs/59VT7I5fsgK4qpX9UiAm87wZVuAIkLe3090jgu+X0znw0JdPRrALsACVlRdVqIV9vX/3
A3cLHR1l8vr1R1JiuEmDlXAB7aFDbE8qPmk98nDs5c2IAmS/RmrR/nQrJ+Nj0Fb+STDIdy+T2F+K
vEcb2KADBJ+Y9nFs7HdTwViDjhEKFOJ0jLBLQ2Bigl21oMFA5mrFkaXvPk9IMk30B9Q4K63yCben
2rCNTVJJMDV/3+V/sU1wyaid6mJxqT8mpkjksRcD6Dg4cXcXiRCCKpUyuzIhzMN4numApVXyGa4n
O/PtfW+pgx0TzTn8dd5zI2ZKm6IR+//NCbcFItHF8nd8iCVNg2jES/7h0XnBZTaAN8pGMI2isINg
wt+tNODTFHGVxDEDj+pga94l+o0sJzsNAOIh0KmX9j4BsYUJVsUANZ5neXpQHrd6W8UiITNjkSCR
IqVRRL1Fywu1LZYnSF4nlRj8dN4ddl8vHZh1tu3zjTI2QlQqGanPiZ+rIAx30zexLNeRLE8sfTTf
pEwoEXLQXrQinTQP2girzJ1GL6D1Gye5irCpt7zOayiUHc9+G5O750jR290fXHHI+DwRcPkAi9IJ
ooOzT0mdtgKSfjzr/UsYAmZLTuIwGhM5GkWtYqs/wRXOKV0k4li417pqavQJYyenZfPF3wnWnyX5
RrPmMEWFmXBVJm6iGnOo7PaDJyVfpIBVlq5w3uDtYglD9mE5c/KZ6hF6BtvLDYn/MElbsb2Pp5z+
/KwTAEwOWYDoN3TRDvvNEop/1x7VsZIRt6EHnEEhsj8HwkRGBaLEYuqDWAZsVT9v1RnstJ7qecIv
mWfnBREi0Ba07s7YjSkP3xEKi+uIYgk1sydvta+zCo9L1fSMLR1EGypfyPKFD3echXsYaKZoqpch
BynznZY3VWdekGTy5Xgq6/9Awub9BKW7HacUlyKaYXgo/UgOvB5Al/EGni2AvtnKqCEbajCunYvs
eothJVuzBYmAChE2fCjtej1wwPz/C1JARjAuHvtxOFlG+O+GAei/Q8ac3Db1xBtBzFr7F6yrubTC
5vwN05a/zykE6sY8Y4C/e8xlKgOU8gdiLL0ldAwSTRlCb721lTujmBtT7JwjfmHMqseUn8TkkcPg
w5foN4ik9/6PqWWkNcPYsxVkpF3s4mbOoiMihiebPazJZIsg2sEwSxWT5oXL9MbZ+CC7aUEi2h7P
DRv6g1xxD7+6g4yrvjJWE54wgs3lMfFeUBjiHyDEIuVEYX7Ply18Iqh6FsCHu2L33w/dGknWOSR8
uK++T4jqW6bTIGFtGOEikcLG3Slnhh+eDPWaKkTENN03vFQqD7ch2FjGtkE26Xxg5hyOqJyPOeL4
BtOpdoqZl29SIIh56INOAVT+wcuQ19gZabSV8VBgKTr3Hey6HCskWij0JNdqXHov/WDK3PCdmHku
+bXEEJyb1sUF29ybcGFHshGTty3Zw5g8q9hWzFWMNvqmNVDqF9zex+TtOoFhcKxRYb6lM2hXXvKe
K0QJMigc1QAdAXFJpTxYCqoElCVvVlmxze3wtc1OazSo+WKQIrhZ6SwCvekQEJL9hwAQjHQ1eu6T
DlMCCwo0iEKhXyTY/gLq5jjLWed0G+qymvpYyWnBRY5eUOQAB3NZ124uufF9xTiSGkb+3+isUFsi
AqNoB2ICE6kAt857cOk8Q//gmZgB3/OzUz/vyVuzCY48xfp6G7YR9CrHg5ZN/7VsyYQTJC+9yCuR
C7Lx4q0805Nhf1cyCzma3L3cap/V4wFdl2gb8RjkO3TXTv3L/0VXe9NeHNJW6M+GQHgiduthUGdc
aHaWn834MqC8Z4TZ51v05m7soad5XhzrjFvGdqPFdPyEd4+VFTmUGjYaUEDGa9O9Z0zdRWQRs/He
zl2V57Qr6O2XmdY6e/XAfGzuS1WQDQYpABbBNQY3PrZgxXzAXV3yp70W+u5Ddi9xP+htU7k/jCWG
8zyCeaVRsoMDHKxrWkE/BkV8IdWb672S+CHkDrGPM/hcpEvpQrqs+PILet116uk0WGthHqufCpAM
dFHK1MFJj0DwU0eSbGS1cG4EXs4qe0QH7zPZG16/ieT6EQMwN+tVOVHZyDHWjG/Y8BDxAseNBq1K
Ppg9+6K+yffb0MrZjb7ViOcmB9l/x4DfM6iZB4YrZ0NzINQvNDXjSdqlgaCvL3C4WozcFBgiZdCK
akrP6j8yk6oEI9qnKxoUBVpUp1QwseFuFqzm3pvqJlsaMMbipi769suUYW1k53DivFMkF+9oytHe
NkEH8uwu6Ae96fgPDqAjq9+hseI9ys0szFp5mK08eEMdedap2l6b0mZKW54jpfZAaz/ZtQhAfqxn
/GxAbmhMP4bUsPP74vw+rnQI7vtDeo3NO3rmij/1uVbcNi2eKCXEManJ13/qa1NWJ6k4m8LO8A4Q
e7bTYEFpod+f3O/Nx5eU5bygRLP43W5lhEiiZy12LjNtSot0kOzo8635Deus69qkezh56UqNC4Sd
CFhWSFizUIOeLl3MmbJIBu57dQ84qFcnnp55/b7oX/lQjLDf//tTYOOqdCodD++nuBnEMKEKW7Xj
R3LZq9o5PMXQFQ3BHvaB6Jtfs+NmJbTjpD+y+sC1t0f+qyFshFUasxemMYWBp36t002yif19k9X+
UbmHhH1Ihg2/bRU9us6v+4zibcc0cOZhrRqX97UeFEjDbNEU6RiD0GUn+dQZabISb/RhHvOdtRXx
jmxlTeLfZpGsW74GAfqIrLijTpV7mA9Vnrn5q2lPAIpQU1INXSBCqb+rSdqXLlrPjohiz7YT6zWC
ucqizfXAtIU4DpOfqVqseg32wycuiGNznHgm+YZk0DJUU3UelX0vqdx07kokfQdKpS1qooI1pOaO
VIjAfV9LHZQlrKUnaSaeGYU9jPBpcjEXJsJOKnEg+b03ihyWVKU32waZTdib8rQvFl6mnMUgIYHT
lYcxI8t7dGOou2RaEtnl8jrVILMYVnTv2KCGTnvkPRZ/Q0H2d2kJMLJ2Z8qbvtCNIUKsxkHwbSvg
HeyI6PuGuCvb8v2G1uQ8tawOSj8PZ6rFspJioQAxC9HmK4ZxRc6PSbvYBTwOm6vP9LxMPLulKWVJ
Ha5EAOcoIQMcccIKBV8emu8waAMk+Ga8MMuLN8vefDMimDN/RIDzZ+nbwrouSJ0CXt6aH5xqzlTA
jW/jQkzi9xWyS+48vgQINILaSSXST5ZQKoa/mSv64HDfa5SElQ1cQzXo7POgol75RdikzM88axjv
K23AnpQE1QoQxte2thajdXgtEgnT/OJqfPBFii7sVq/YFncPFd5ZEuRuC3M8DBM3wqbvfhai23zS
dl77cZxG6C6aJoj6/dr53LtgwKVHawCtt7MKTkyDMvzP3I9+UW0gu0A2jTReLCWv8guEpEdq+I/t
16dYyVHfL2q0mUHA7+dk6BzCCZncfpQqlTRbndEBZZ+PsKKckcmExfMRikEV4gLFhg3THbBQsbU3
Wvfly7R5ttEzqiIpuIUWjbGPNtZf4j06edxu+K9O9K8Eeh9sqyRZOMaqPy/teLuwwF2Ob1PM/7Fe
9vRzkPX8i0Np7YIzgOED57f/IjWRTNx76wV7i4gSPPu44s4Loi6xpIsVFmmlIYQHiXK2QRK1Y9ot
C66X4Dyp7ke9K+nAquWbzJnsJ6YUxtW7JjQiz1ZRCdn7h8YmaNIRm/WV0qYszgWzrrcyHyqrUM/0
aETPPeypbuIBWuW9waL3pF1O4VhYiCCF0igoanBwdj7qUHS904ar+ftQO3YIVHd2b/Ujtb9EGDSn
6TC+V0SbNjky6fhA69W5PArJUcnJoTFbj0XfQbpXkGcdaSiiCVzczf3pY9qTjUhI6zCm91xCpB8I
kQKBJXgb20jPRVJoIUKvlzxqRvM4MCiI96w1/7xiK5GbnNh+kPFHqKnJ/S9lV2KPggQo6WV+8ij7
pV13iYK3x9XrnB6HH2IAw9y5t3Vt8vj0iUZnadoS1vQyGezr1CPkPdYogMoDZPm0WLAjDWpoOfuF
D+NgkQx9uMc1cA75Lt0yztAl/0nizxtNR9/PvYY0UDlLac15oYk6s1Ut0LBhVWJeNrbWkpQD7Avt
4j5QWVAgqW7a9WRArArNq6l2qi1E33KZ6JGaY/jq5f1ooLbGrgDYIAHv9ZYte5L/TuTFl/fpXJ96
qez/cr8oM4aSAPBT4ePABv0+rxApXLiO6/u4J9DBnGh/GyiyJCU3d/7QcrmfbLwdki+8L7HbUFC3
/cjjbzI76MJDCJl8ipU01cRe7vxJDkCRnDdQizmUwnGxro7172CRwJlh9zZknNUmWcZANRn6gHTj
4PjDFP6PQ+9Ys/MWvDz2zYbbNmYPEUSqkeGrJ/hSzpK86AisK7FSEXqEel4tgqJSFo8LRt5uV5BD
MGknNVDbAIDD+RLTgx3x5vxIAFYSP1Q+tKnT365A1w7KdplW7nugPdX36RR3kLjqf0lI/ezTWJ0p
COKbEX4hc68ajALt7zbEYfdMuJicP4B7tUHd0yMiVzyJ1LqE9nly0AP/FzpeuYs1An3BNtUcd14U
P1fQtp8zrKHBcXV5/yehd0IQa4278dF3AusFWl+eM0+1tskGBVVI3uYRAfBh8wylYRZKAKxws/gV
bbc7nIAWLQ+MimY9NKtwas4H54RPvV+L2eU5hhtp8Hg0GtE/b1oklxsHX67l4DXJMRgX3DsSoFtS
mCNHk1PMqm1G7jOVw7lXtzwnV4pddv29c8crDOG7+31ljOsuahLQP9PHJ/CVQCM0RXka/pYdHbAK
vG5VLlwe/kRfaaei9AnCsY3BnoNAO7noYQFNtj2m40pmlDVSiI3bF2kk9GMT+b1ftTyONk5jYjmi
gNzxve68bkYDd8RRn9dZlnzw9BgXBOletPJOD5eW86nCKPfjtlRdmbOVfAeCdfykhqbvs8hk7Ze3
oKYCd5YCj6ewRjl8tioLQR0sqvNdmfpZr0hnrpBDX2c4hVsqAtXjZ/m148Q4z9nz+4tDH/03hPg8
W60AGnn7N7+C1gZQmQYPeTVcdvM7DoByNwJs4u8QYQBXzA4eyKEmqaRFV0wVc3vQ1RujFp3j3spO
cPDPourOMYzDc+Rrtn/BvL2bmhwrfCWA5bVSiUm3TutevP414HHO/iBChmVVrXqnDgfeBRpOxGwh
jZ3bgeo5h3jdRmdTHHUaIB9zNf5+3MtBl6n6KGFVf3bX1fUJ9IPCWKKbb/WpmY2YACDShw0xsrLZ
BYcBxAWYDvyGevzTmE5fBnPVYf7oTHmrMwA01g/I5y9b8lGRmwwSD8C05675S1pw+HucBQLcvYZz
RH6WNH+2rqdGv6HVX4W1WferCI2WwfC0oS7ZdrlUSnKjJRkqIyTMk0ACRJybEajrMXk/gCboVmID
T3FKFNjApuT0168KrNZeZvSna0HGayBiRH0pMR7Glxhx7MaCUh+A/ELHElQoCLkWQ6CyIm9ysWiW
KbSOssbbYBrib3RAw2iMOMUmUxsIqC9qVGNYtjxsFyZ4nvqgQw9K6It5PB3Jbg1aSySOwKzfJiLZ
1tep9Mwp0I8XQXi5+V7vk1nfKuYql0asFLQzDQFpxEAvB1sfA2nRj48Nn+Dcx8mvrksYZAx+ga/m
P3AAhhd739ihbmWp2aVCbZfsp8FEhuzedRvrGgdivG0+WhWsxhl2EOn7+/15nPgpozBJfVQlX6sv
SSHZjuMunYNur2qrspVgNX3nPZdFiOX3NmwjIqsmGBSI5XkLPyGMX4/J4XOI7+yuiPCtRO/5DJBi
DpFqT4HSH+cRd+S6w1eHHLqdKGBgVsA9saQ26Pq+DFRqfESKjc7DSbabceBJN0rN62DveTJnUnms
6esOYwbWBkHxi0yzzH22jc3ow3R36ydYqD4oNgJVnaRz0vnqJAudH/ZIWDlfWGdoQs7azqlV56cj
bSf7a+RhVLnPJ6KKh7DhqE+sXtujfacxwq0LtZou/2EwzSfSTqQTv7x7nUrK4zCfgRlFo8MUYjS7
5dJRB2c3oKao+wzQsssro9jBH7cflnow2cuHfE2TzV0Wuf8WCSntxjhxkywdOj6aUlncI5yu3fPS
MgkO3uhzYjFhpqvqDeeRLfTOZhHuXrDTTXsd2KSRt+hLnTx9fC6kwhCEJpRQB22g/qgN/ghqTk1i
YZvXsX/KOElVnsLtLEVATchUnPzAq9iAldnrsnGsi17xzTMSzffqF6nqg5+zQf43Sq/uD/I6YKPt
S1w5l4FY+2Fcae8Qyu7rPudIZd1nm7Pvrnv8VriQeXWq/YB1E/0ffcXw7C/N9Cr977o8T9p3cBtI
h9SDDFwatglVi2DGstLzRWmUpLLtSSjVxs+0kzxZVWFp33jAj1WlBP5vPAmj2t0hLiQsaiANBYae
n50mNk/h7DZnnhp+P5SGFI8ksYRRRvWTq2xBx1PehymN9fu53PbRlZmDrod/n7fc16HOYXGqDp5A
+d5HFL5MO2rwsdgkSUUbtgo5QI77fi+tCrGnBzyPl4sL0xlRWRDnGVo3xN1pipJZen/hG+7qRLAF
T3w/WZP1EpP9po3i4rNCfyQWPvQnLjodqGxGiiNmsc2bT5R2OQtsYGR7GDBcrf0kYMFW6EcvnFOS
moerxoCINlRYjzBIViPYWshCtV5gttj1+mnUVoSBC97D8FK6TI/Z4cSLPnvaEfWJcRpp6mzQ8QGc
WIU4i6ArQoWA3JK52/yCUzETneLhSjtRTWru6SJ29a7fPfJXxVYK3wsySRGSnacM6LD2QsdHW9eq
nZm4WLKCxGwIXXFFt9i6wXG4Y4ZVxiR3PTlkExjhoK/q7lzOFbueN2nG08qohMALF5UkyUpMSCJE
kfRWuY26zBKpjIzuxhnGAEAtXbEep4/fv4Ju3GTSvil2baYzXmY0TPko/4eVR5W2uh/mCq3Di58F
L3kcALA4XmhWBaNhMrV7Vb8QWA/5gqHmUKDQQ9JK2iltG3UxE2TyBQQFLeE+IzlfyfATMpsk7JWn
F5bekIhK5g3ISkp5ksamOcLCEYjAK5XEW0P+QHNI5aey9M2QadauanMqd/oOAM77xNx4tBRIPqev
s2qJdxICx8AGv378ohdIZYRBiDVQVcN3vPfWJ68kzQzXsJ5I7gaa3aoYqJzE9iI1gqd3umi6+MRq
20w+QHFlAqFoRPod9i71oVNyMOTa0j2sGeyjQNkesnppGMDp2EnKtVzHEBbOK98htofBW85+UIzr
21OuaBSwqGm1dXE140Xcpnf6UIX7qxX82nmOeoDURaN+K/G8xE7/iTCz7JPNjw9O4BCOV/Hfrvc2
B7qoyDcccpS1oo3itHQaHpW5mVPVPgsGSIjHNIfMI0guhdqGq/6WViIQl3tErTOxyYmd9pu/9MZL
IxHlsUSgB9ClZ+gfviIONozdjsvQv+XNXh8F51JbdHnHsP1bxtOm88Dz5ub+uSVPPjI88RV6N6VZ
SK6Ky2VKSTMLkBWWFptkEhJNDF8i4OpoWTlJ1QjMsGeDo8X4tAHBfQBfDdUdFhOjTFqmYSZs8QS/
nY2Ivq6XZM0Sltnk/8DSy5Qp6IoDNzUZYW327u23WfwAZ2YnetNy4NGCUIcbFzYjSehNyAvcs9rF
pRxY4TrZJjXWbLhNa2Y+ZdwX4r85DlV91Ai34YemaFtACB3V0fhKFdYbMsvSKm6Xbs/pUc4k9xnQ
HU1BzXUeaQazobXYFmRXta2xqlF49zMJxao0ZNtQaKm6kNdOCOJ7m3eKhcrwysX/sAuiCN0vWjiR
z0oE8NYSRIl0BcyJSewihKDLE+uPJaxUQjGNATVs8H4kQs749R5z3fXhojTu3BPxKH9Vf6xvYoQW
7ENCHIvBjmTHLmBcqbGcOXDROlTAWiFjGNdQjnmDEwQFFazFb4xyTq2sxuTIsdNkW862VJoVQk9p
G3HxjcHDRn6uy/309bD/nzCfd6VHX0xJhBOQvG6v426ULUULbTLk2fvQ+jkAhFnsueuM8uL8zshF
oEjhFvIBx9lFGR5UbAjuO3mBVlgaGvj/+hBev5Y2CfYBD8OCIZzZBfieMgqpOEpH1hlkHG20ruwI
5wZSSLKMzS2xG6R38cs4wTmf7vYuAWGhhl5Nszj92Fi90bTI2LhZMRNFigQrOLkYOsu1w+dOQB1p
db0b1HfmC9AyTlEhYvs/cjc6n5xiNjLECWTfbBYpq2yulK3cOOOYbOlnf1W4UMa8m1JEEsWgadfe
gXJBfOPsF0Vs3ryr3FjMmZ2emXScWCteGcgoLFuz/3c9HdzgJ9FgAUJotx+/kfNdk6Ubqy2UhaOZ
0DR59+PgKru1GNw4S/crdsydy5ghXuIFhI2iTM0JavD8Uv+0zl75z2IXJ7EkhcOvk3T+tUFZqj1q
K4cFTgUtz1sV0nlFiOCAo5TpREFKiMPfLAz/aHs72IPXT+bH/3zJvLZwsDVZtdylXeqBAOEF3aVk
NM9T3r3h5E5HnOQl6CQ9IpmHLvmfcrAxyIdHvBukjhwRPaDw+4hAqHvfGnHHX7KZWCHgXMSZjy5X
ZFBHJ5ewsetEorPla9HSQEvztMJVUBVkiTptucQkyURzI5o9uGuR3OfjK51ihmlhiJjHswgkOmOg
7vzJpl6/NMO14wq/fCILNGzWOjXh+ONvvAIVNcLM5AqRoDFdmdilRLNGegN+CfOjDxTXYL+OCmMR
nk9GyHEEyzlYgb5dcm76ltCMfhFM/Aqkkcuw+0ujEzzY13cL87j/mSOpUvHB2LJcrCrMj+zHQXIK
8FY6g1t4SL0VKcvqXdLpl2bnTx5iG2kAEu+xP/jInh9HWMcbAzK4MgsvFlqZTYsrLsnrPgdnLNMR
l2laFSgnxp9EXRVor+/q5qGSp/ZDlMUJwa0VXNzaSYYNRk2X0Zd5VG3gEMqYADGE2d88lP4j4d+q
3nCFCLZcAPWebekln4ESIC/yV/X7GlTXS+Svok8+4CYRPCdhKX1czKhqGk9t9T62MWNvUzxE1YWj
yXZHQPF+lyiHxmpsyVsAs8sgpe0zPivObEelbuA59w+3cr8OH+jk8CzyBjRMg76D2U/ucEMNX9zg
LHcReQnz87WrfiywrIR9fPJ8CUGPyYIeGn+z8uv6VpL6V2d9ptLtJzm2mCB6gJgcHeskZ4nq++B1
Rh0RdMXV/c4ITM30jjaBc6iGYesfd8hSuU1m9VbFVBVydqJ6/OoPzvlwHKN3g0WldpQnaDPK3Ywt
OOU7Qvev6MwYIaqt6eCYZpnK5pdHS0ym5UI9Jirdnj7JA9d7HqZnF3ymtMG1bEuLMqPkW1qKR6hC
aiMxAeusg9z1fJWyZFljwgtt0M/uIay9hbB8D5jEv9PmgzgnP95tNp+NIp1bFz6tNQoWo7KYoxXX
AQNXHL4/IaaZSiGVRjCJfEOYoQ5vrrWYCiABW5WRv2+z38bbhlq0PKLkXyLFRuQ/wQEYt/YJ9Vhk
srLlcChi/uxfq5Vh5F1cn2beC+yIamqkMD4g6vaWO41IcaCRQNyOJR0xmzW9+DqDhi9Mu6gjKj/R
A6kHq/3/JpHGu6NxLWkh2dgeWgWRvvN/VWbvXUPtPGuXeaoUq+fVjCSjSZ1MkViWwlsL5DqkmE+u
VHaRuZhl2bPxdD0XatZoKpCe/AH9jD86WFiq3dci90/y9UOZI/R1zAC/7WK+fxmYwnWi4gFr8Yv1
EWa1eh0aTn4d04obaazfCfDwpoVf3e3x8Jrsmko7NALlqcG+RuGh/tfvOwMdiJvjDUqkds5e/Fdb
af5Cvfsb62U4uwMLVFEo4R4eaklV7M1Rdgea61dAkdtJNHD/kzUr5GSuv3JJlru5x3LSpFSmRCbx
TY//WAUoKsr0pPxN8o9LtiMJA87iDK4xdlVM9M+zuT7/B+MITLCy8LviMPq1+am7W+jrLXMqBlxI
lfgC/ZQMl8w8SCPZaD8xVUrpEX4JjNGcqMU8gR9QF9Zqh89kDw2QgnoUeN/j11GSLKEDmmm98g2E
fiUiXcaRJgW39U60hwXFf8DuE94MOU8GY2bOQBIRGHKZ1ZV51TpwePzUuXHqNYv+DrCKgWu7P9JU
8K0+BDRgYkEeSc8WWrp8EmzmBYSjSmGNMBWjnmRTky8RdIYpVuXaMSY1UUpAC+zGhljg3Fax00Pr
EAq5AQJNTqsykGB84yJ1alUsoZ8U8KyLs54fIUYBhq8zIp1rPR96VvXeUHRwZ3jmFIC2Dtcd9KES
bA59OOvvgJYqXVOTcgcjFSHOndSeHgtsjZ+VGw8iSOQU5Z7AKgJ2vpRmAa+nx8j5qzOGdFz5DBEg
AVjXFLn12FOTxPM9eZ1cDwUE/1zqGpRSZx+TcuLc+Hq4jQivE4c/f+Ko758+fwZEsxWaeGS1PATg
JNCwEeQS59jYKdtlQAQSzNf28dFYSN+qJBqyOukXaup8AVsc7FMbYRXyEGbOv2T2fUcKIHAifzaP
mW/yt84FPZqu9sJJGIyIE4LC2M0oxvQAJunh6YYVePmVnvxlV/dMCOpts+E4jPb0mD+miH0M45H8
NMQfKNj5mRGYAw6U3kgpkPGIEt/b+haQqcNQOq0fJlKM7zjbEa44hw79ghXO7eWLsec9i2pGExa7
4oqEt7RiOAvOciwWhxWJTj8f7Opd/nCfOeU64veu1iv2+Vn27ZGVhLfnsxnYDw5a+Mw5KBUYRy0p
mdK48OLK8hOD9JU6chcvOTxkjOBFfa8pBaFj/oPKIe+i+skEOkKjwTXDgGAoyMnfdmpsIP29RE3/
9kw6mgoaqdoAenhQO4V9GqwezC7DsIIyyVZ2AbCL7nGoxlco6JDcOTeeIKGkOFgwyqm8gKaCXKDu
Ls/K9eKcbKgtrBMOrZuIMb+KEz/twCbmvTkPnwqp1xNIhvtxDe4vh7s5BQdkjovSZI6izjv1uwVe
1fP4JatkVymGmBjNIvCHEAqk0HK1o56HCPJuj5CPh7bwGTxvdmjjiB5w1PcdwD45LHXLIScTg96d
xiaRAOHdfsEXExW+RcHWaOCeyCHyEhVDqoK8gGmLZ/GeSgzuTR7WusjKF88h5JsFLjGDThh6xNEF
LBWzeKku+/fQRUa+TVrYJTenNdbAnozJuz9/FRV+OZticFyyb7O9tOJYlZCHtkpli8Vw2tRhS1xi
ARyxH8UlqaxIb3TjRB7pYtdWpeH7zWh6OJLXRKUmIs0+iNEtyK31vYMmYgUF+u6ufhR+6mfDhT7R
R+SsEjF3wfrXnvQtfgHFMkfXZvSvXtk9ftk5z2Xs3jHp1WP36dIaPknx1i4xftfNVfgBN3XA3JQx
sT/oubVsr83zDgx9gUlsNWtqE+asc7xJ4px1b+2uDGRyTf4byBiTnmoCGY5KXAWQRsvWqV9ueU/T
+5a9Y6Afpfxd6MxSS4Rx2vzf/tCSBXPPnEfghs+RWreigEylz0bPfPslzOc4Ro+dtQBRcsDXVN0P
LB8q+0ORmxCBFk3eQy5uDL7uWqX/Bgvzi+WyzO27Jnorn4EceEyHmY79ErMoBjVc44iTiS/qNYJG
0GMxL41ZlhFs6fX9p1GGxBwqyiwpe13nTdy3H4NGITz+WehK/gNi8LxBTSfNUAbk1ZHv1yk/vZTo
c3kegnV5AURKm2u78UzID7J/mNTdYpIVE/xDFzS5wIRIJ0cGMX6gxuXxE4tdutVcHNu69UvKuXVX
DJh/IZpEy21OTf32flsxu6oW/m/SqeWStRiVQPQHGp6221MsG/3B4JZXSxdeSECYhrzPC5SCV+3j
ddKQ8/z0MY+MNz9NkgWDwijh1E7Lbm5cph0biItuwF/U34ShJC7xStwU0LC2qj/97Y6C4/GLvcXd
02mLzZ4PwM9V4sdR6JM0q5cpzVXtb3NrCcNAUEDFY6oe8A9PFFH0eoGGtyosg+K5xQbIdDkKNmdd
GO4NsIfY6zzwjfNE2Rcqo9bDs/ebS9CWieQ1n9vGTeFvxkwcyBslc0VH0C6q8G853/NpLu+wvdUP
EEpZkAYwmAD4sUwtJrRWrEnt7Nkkdd6HeNe1++Uqe1AQvhHCVIl5hG3NFF1SeSv0UAM35oXHishD
Ab+vC6nRcmKxjqMnGquOTAfMB0GTe9PQ4ea0g1G91LEVc5wJoO72FAvwbfqwurq0uqEJpOD2EkcT
QqMKI+spMQwHi0rq9VyXsMcFe1s3HaPFsL74idtxcVJrC2B0KPcOuvvGLnAXHX+effr5zGsV5Ihr
4fdXZejH83vST4dHEG1GIRyXBnH6iYvUTYgucGnP7dgnk5a1W8RCKba68J4uzZXYSUIegYseU1Xv
wx+VRUD2TwQ6wEQru/pVZYDN20NXk1T9l4o5uFKRmeK3+u6jXirAZIDU9GoZKmHMYgv4oIzyLnQf
wkb3tuYu13fR+8avsskFAVnpx7krQO6VNQaiJotzg8v0vnD7XqigrlZGpNffl8Z6eYrymsSQhWRA
g8nxB7Mx8iN9YTHSvZRTXNiy0lSwaA4BRQ+j/6UZYXbzEMSFv2D5+1WO84/jPNzZi319K2E6brH3
9GUH8vtiB9X7j4w4RKFHcmTENdmZyyvmpKOXuBM5L5eY426lgI9MId0uk+gdODP0BeqWZzlUmt3I
tbsE4X2x12YU7Yr8jdPbJD851N3mXbOARHO0qdZ7MFcanL6FpoY7tIehIkmuC0cxj3BEDM6ZZ+4c
hdqiOvL9fJUlexttpwPLeXqU06Yk0wQITufzBoCk+QHOftls2ZnJ8kz+xk10/vtjrzqVetz3Rtsn
hT3XvEGAocTt6kf6Py45IeOIJAV1EFCbjJwzZL8GbnKb6gnSJ2ddJ5QqKmRMqhsxtwSIBsN+4oXy
D1mxfiw6a2lZ4Td7s5Wlwt+q56PS9n794No/r7rLPO+qFBzMT6m6y5voRVVVfePwpAExbhFfkNke
piZ6KNNNYDn7eYi6YqjzKYb1q++LbgJ8k875Cf6TXDqhlaiecbLuEn3veofyv0mYnZCQlbcUoH1H
QLKVPvvdSowzBk6Wlq3veK/VQstWiENwVhqypkTlpzUqUVBzjnu9tNgeGdpLbpOBJZBWqJWZx2gL
M6pBZ3HW7NrSd2sBDH3auAT+9V+LUzasVXpD5Ba2wR6u1xEDg27j567EJR/F7vNq+uNSvu44r5eT
w/FJQ6o19iXFpLIIJiu60rkcg1nwzuFYJ5VUPgYawphinxISrmC5xIhEUyxw9W8WWhsV/VTl7qQ/
/vqofNfl9iuFTpZFPGEI6UVHIYXtTufRPNThhLaIrUp2WuoBhc1AwDc5MNEFbR7MB5eXuAgVDnRy
kcCyhosxEQxUuW/fTJNaseiREgEiqUH0cT/dSWbMDNYVaCSyopcW3wo5HVMKKm6LfJLwvCwNSsv8
zB6d+hbhu0eUi+rT1poKz9ExT0hA8kq7NFGMOW5BjRKOGoK6RxXoFomsGZVGiTqgzXZr67+WT77e
stCHorm/cgkkjeerEKpYNVuwqqGUSVNe8BCd78pIjYtfGJoa1H61e4guOPkqhcCT6Yt+RexLsJT2
Wj8X7+w0Fuz4LfdYQVIp11hdGjKuoV/KosrnsY+Vak3RxOumsQMiYIhZc58Sb0yKx/559ZjZe9CR
UATr0OWGBjDnSK4nZCA++P/6JP86n9YZmMB5I5GrYRX09yvQBKbo0VTGyuM14AxXR4jESKssUQJd
6spp4/PmS2gv8M9F6QGQsk9qvLz4kK3XYTvnAV3QPjRkV2OEvdvKKT5FF5v6hv57ftTwMY29J8fX
l+kea51dtKQw6jyV0OoLz6oCcEHQA4G96rVOXAqcfg03J9aSXHZCIu28UFbKs51FNIEmOIzCUnXQ
AHeQWptLTl5RLYSUeIyEj0xwjNePDLPlyKvl3wFy1FaIa7VVJGPmvcivjmQE8QhWkDSJX9o4Wi0s
OBSM2RlYrRTCjxAfbyl4+9aGTGowXinxHhoit7SvH3KR23wNJywDLcgov/brmtJNJYsiDR84s8a3
mdC8dXIfxVmLFX0+nGEEVewTb94AIEwWfFbRy1P6A/I3wbvu32hSEuTyKyG7VRt17uTeOoUP4+DD
BrpiIRkHlwYtDGtgxhYZ1RgxHip3H+UvFXP4v/rjLB4+2F6+CmzftenRh+eMEP6M/34LTzqZhkeC
cq7snb9jlG8w623qaNfavbJyAVt1viQbhYrHCNKSshNtekk8rGH4UF134EXfFpJyMjVyCKdaw23g
Ou47m0kKwhYmEOqRCN5QYZaa8kYn8izEk90K/Sw/QjwI/65fcF2hY/MYBl5VStPsxytwfA57U2V/
GE+8KDL+cumvMCND3ts4LoHF1/eCzL7E8L2o4+s68OJ0mKK1CllxXJlyExiB0sDMRrn1bAva8mW1
cgWxxy67a+5jehrkNcUbwEKQv4Z9OoTGGl/M1MXVtHDtBnba84kqqLfF9DB0DXVKilJCgncDM2FU
yhvNJ0fM97PUMrDFXEphzNsiIJZLcJwqauftdIUVScv/yeMFY57BMTaU1F8M6nP4FuxGNnvbhrJU
+QArz7LAKH/tWi47nWB6+WQtfLp6BHgQb7ozIWMy0d79WEZhCykwLWX40rS7ZnBSx8kFWc71PksF
01K9ruw+JHKdE2U1RZzwhDXjRSqyaJdYH9RMxy6dkrkeEyTw5WKB75NujZPYVUXUoqBEFQAOy5MQ
AYBGqwcwuo7P1Y3cu2EGFws1FUcsp8tlppwNvFKgFIM8GHyt+HzBxiYY7REXjnYWYFZfYsV5Hotf
uyOsjkhLeNBuxBGoaywqojkSceE4jmM0mzf1VRo5c4LdC1czfdmpgTy1FNwhPjfX78SNigkojRQL
1+/hg2SSd8mFNKLKUvwdsRkn0iu5tktVo6QWiqApIyQtVHWK1JGBDbsRlFX4IpINlldoNURcS3D8
el39TqgM95Kp7f3EanNr3/d06Zd7DuutmZzD3gBUeXxg1nIUecSjMDNaG5dmlYK7fp/1UvMxW5tB
odz/hX+b7dF8FnKyZQ2lfs072cY1pXihxxTt5qHvwelQamQnVC7cEVjZRzdRgihkYU38V9AUcV3B
SV5tSUbzWrEtaGVYWSuCIC50pgEMuIvR/sGhlqHRbIrkGTuVNmrVniUteoXjTzjV+Uijjh7mPCih
TMaaHVXXA1LIQD3JnfDSYvA1MQpZYW7wcYJ/ysNF3CEVEB6VlIaV8twjdIn69VLBSUPVuEjT5iZ1
hi8CLh18Nhv90IJChHa5uX95tTq2vcEF2i+cxvWncpQ/bcVVXHs7Riwf7eMVke/RBQjq89t8ZRlw
vJuQeHFWDLHfsEJxxBRMEHbZ5o82Lagby0LVDheQWxr4xddzU+Jh90QGaEnEg1xxKOc/+HNXcpmD
567b7G5ER+NwVSuzbySe5Qw+WymmIyI9eiyYrKDShR5a+yVtu49fQPRRjWbY75lO63A7KrNvzMWY
6mJTrZ1cw9d1bTQ288Gad0th5gY6JFEdqqwZrmUyizWCbYsuImsvjIthEPZ6H1wP6GL08i5XfDaS
fy4tjfBr2JS9uegHiK7StmDBWJf/f8y74ijEullwqa29Ben15uF78SBaQzBTcqf4tmBHDnBYexc3
gHSDVC+TgUV7XjmNl9W42dAxRkz/e5urYlj5iQ6tZ2/kue8UVUalSjCsJYNgXcvyJUcTypyZq62T
Xe2WubTsPPhf01NAOuS39i5S39Pg3w7NMcV1K9h6zTBaxgO8pTtYqjuDB+69IU4G+hnHq6LxNV9Y
XwHr8BZ9Ip4p4ghQKkRz1CVXzX0kY/OaYAze6VQvSCuDuwCVUJ6WSIrs7AuK/r1PNyFClng3MrYo
vD7yQr/hpVDEUSqONWWF8SVtkCji8EA4kj93AxUVfzYiS5n31K3z0r/zwcNnkihTEfF8SakBSmZL
+z2e4aUx6q1DGLl/Gisl2v36UoKmhVbHQISHdllHNv7EobicInM2QTW2lnlypXfeahI9rsi5KE4j
lVLZ9rUV+nySuDbwj6ltVDdqiMd4eG0uwl5GjcU8T079an994ZlDxwDo64NkV0d5u8iJKaM4u2sY
xR5VVCf9hsF4/hGWTnA6Cd/9D12exT3q6ZgKYXio9Xw9+HIPQ0mesFll9W0J1inNc2SEOiGA1MC5
L9uBg1E3zjs6Zg0bKA3rBc6i2qoI/e3VnrhcNYLDRviIyYeGpnLKHjI/mAdr1DDd7sdgnDOwo1Li
OTl7J73oAdKEd+1uWbYZ910YbRPEUF1CkB0yxseayJoJx+wceWzpdL8wCgb8VW2nD5RVp40CMTuq
90KAjn7tOeR/z3w1hwqbSA0TYdwTadbTfHBuBc72oU1OgXBqvbx0yJOmzmjZ6P5ovOU7zZQDdQys
YoBSaOUVaDTUazAbL/u7Wf6K+XDogUDwQ5tI6LA1NnVT/s4cFbTeTosZr7BHGjsyolW6Se0Txz5s
ED7RADEOFMSVZqWc4glg2Rnt7qfasKutRv0RqzLJ4S6ZXg0vN2zHIW+Km/e0CfdbSBrn/HUiUGge
Tsvdk70dpUwUR31daNWn6o5wbzKkhLlNUuKbzXnZyFavYRsc2ORv5+/wvzMa4AkuZ0wv4RBcz5xq
LXINq9NfcQczQekX6yZzsYe9ojVvfA1W85Xa0z1BDpHNeWMVB0TwhN3SvnWxyXKfBWG5Vcdxov6X
gAg4tSvfTUQQ2eabWeWCNQjBFYhtB6HXQ/gusAbUsyLeG1FR81AAPsfg0dYU0Eaen7pTA+D8yW82
iHeV1VCeQtprhudQUKFDfLLEAcgbW+ElgzWpxCoYLzPC0LfkOkEpfYoO3RCabPxeg0qkm9sRwbmK
kKwnzT4FLJw3ZUUcauJCgY/Hog2H0LNIpYuJ6lYdGGqve5FpyMdx6VVC4lrI7cyWFRXT2FYmXkG6
3n4ufXf/JrnZ+9rdJiqRTw8mNxavDG/HMY8LrGguGrKOioYFE2D0ZBGuBhzfOi0aRTeVhiwQQGl9
FM7ThDljb9rxdHVfkd7CtC+CQh8/BCZztSFBNysIe2zAYuVtrJh2ggF/78Q+0lqGuPWmIElTKmrR
2gFGKqMCF9flj9wRNf7AiPu5XRbdd/sNKO1NyJP25hrFI9A3TMerU2hy0l31/AmvvEambcQ70AXA
FJxSxd4cZx4VCg7/R1KBQpCwAX4I0r6tMBb58Z4Vg18VDpp7EqZKG/2IU0oSvAU92WEtU8sPMhNf
jQfD8x9hKCaUaEThmTJpmGrnQ535jEDvETQVawxeFboEfmmS6SPR+Z/ohvfG9Q17GbhgIgo2OCLx
hdTBcLr5Ap2S5wcYqEjXkw3G+ybLMhfGmF/vy0I++EM1Fn8XsfPQRvtHNo2A0zZA1d9LTYQxzfDr
W4gKVn9282PVTIm5KiXQL/AoezbgLDKo/jcF8sXkvlRJjeS4CWqAMWmvtgXp4tMtauuudlp9Ud2d
aFLZfCLAcFqxck7HF/GtCW2pFz6ofeqhkG5QvrS9YjR8TokvdNo7x6SG75Qseh1eRV3rtl0H+JgF
u8x911QIJxb+28gGEo1TDh/tKKUHEY01m+XIcZlwzu22zMZK7ZfpUQyXDeui42VEnfgQ6x27rE8s
F65rm4i7pJw+nVRbmozsUjAONP6ud7pj+FIE4JTeYT/MXm2cOI7PSLV1LUrZ1tDamrSoRvNcTqqN
25JXFRQZIqflin+BpDuwQ6KAi6BOl2Oy4wSJv4bivgf9Y9Hg+lb12tbgJX9UHipA1hfPiiFLg57R
BE8XdD2R6VYJiTyd+rrB4iyV0Pf60cuPIzMgTP5Kz2Co49oE4NZzozkgc5ikiihg7sertPLiYqbX
tHvumzPrHIgvgj3RjwCJNy6ospH6UHSdMs4Pf/oWHcMAJvms6kCGRtPFaH01lXYe/u4rhkXrx8R5
f+FO4Uqwxh060kWVl5rYkIM7Khl++LaMnqutyF6cbTWg4PeAdn/ysxW9kB/UE7XcnCmF1zvNIHM8
1yiKgohbeSCSMYekqgToU5LNdDyaTzafWZhCjbQe4biBs+VsGhv199IKD2xExWN1NDlWKiqYHPnf
S/HmhdQFEjstjXzzFajbTaeqWMt23Zd/CF6kOizQQa2IxmwPGO9RRRkyu09AMGj2axRvA/clYwI+
gUzN/2lETjtfmwKePlB0sW6FvdHLSslxTjD6A6jkcVrFopzlU8YKx8Q5asNxwWpCeHJGICL2zK8E
K9eePre3+YElZqz9LeRHPSYOpt2Bz/wv+N8M/oqHkWbU/+QpqDgyKmtJA2py3p0P+RrJ/2t7YnW6
W5QkvSelxx+T4Ix0HiicG/F1agUp+NL0gAo9YCiudmzOwg5w9xIk8OZ2+GoQSJVrHDgT+QiQ8Zf5
+gmx73vPT3dRWoLFeCPCSf51rz4tvp9o5DcpkFHDt8JTqEWZthHzGrMq7g0/NeVV0CLBb1qwZdVh
fXZAFAeNmnXdANHR8Gu598l/oINtX56fmgD9VquYgl9yqxjurPa9J4v1MLrE1/XokSkGb/gcd20R
QBdU59ABtO/MhOmMNLEofDqqEQ8w8pBFI1X8mi2OC0YdmHfxlxvz/ZiebK2K58EeH72vj0x6G356
kUg2a9BkrmFBh4FdCwk/c72jhYgkKYJauj+Oi0UbjMDxx5sprI9Ap0TeMXSQZZ+5TbIfgkuI5tZD
RAu+Ugv+piqWA80x7P5NKnn7v3uE7ybpPO3WlMg4Ce0Yp1I039UrmCHNxwFJvVivvy8BX7Xf1XoC
w4gGTEmLyiYfJks89uYvp0TWQvVE6SJFBIRgVjiI3kUOKIuNxn4pd3ywJi71WSwYAbJL7gcXvGsY
ZUX3ePiA0ljlKL5vfeKgNzgnQoZztY6AlUPIkqfS4gf4zz6RunC38oquOiZNxqli3BZ4mttFEMab
flTxdkNpguJJtUAhLPzxXOnKlD+5ge+wbjHXLoRkdbLpiTigN9q8g14u/g6c1SkrQ9e7qgoNGkUm
h3ULPELQbAoe23a4i2y5CPv5xcDZHk8LPp0m6vger0AOC/mz+qTYjBYPUh+0ARKiTZojErRFpSCJ
5Tjx8hP4zYJzr/4F9oBkUKYOZZ7hdR/l+GuJE/fmH1tUfOoyPbOWWa6B0iGjBdaR55ul1zuLomXf
MxVwa16horGMYyVjAaphOFSVO5FcM4ybFL20tnwAfNwSFIQ0cB6B+FEHToux8Yv6T+lGaxzKYpT9
mnQoXd4FEL+cnAdjuJu9mSCG2mKSpqdyJdV6ZlM4+8A3jXfFDJKXUmXFfBM5hSdKmVBRHCSiubeE
6U82BYpvY23iqDS2YQOkYfvpuv9MJ1CZ+Wq+Ktx7aKzY6iTN5NCyCHk6C7c9RUTlqZ1OR6UxKE9v
latYLo6Y6+2RiezLjfbQ9QADubF5nUYtJLOpYPgDFxSiPsLKq1vFPVAzLr0lj1oo2cfZazcVm9dc
H50IMivz/ka3T3JhsqCPagsHsqGLyCVC/VcFm+Nh8j64oQqFjssLfuff0hmXgPFnuGitZvd8mHZV
AgDH60cmbEPqONJ2BMz8RadqMf9JaAfM8bRM3+yJEUDiyLBCevFeA1pBDAcDXTJtDYm2gb82+8AC
4Vgy9eCMc4yqXtE7tJZlbXQWcsyh9AiJKlDUOyO3f7Z7XFV6yJ3yKy9L61/FLU+KN7OpuEORtVLv
fKYRW0JXVzFwrdEn7ILAitJfC5LA/HR1gOeNfhSlOAT38g89ngv10VQNXthqU3z0HUi4T5SIBSn1
w4jU3Nc2cZtubjFXV2A9Veq/FMMM/dCrxXXfqmJm25JBEb5eWfrMcm+k/4L06KuxNVq+F3RfPXgN
2dmO94aDTRvdANB1OaIcfWDw5sj3TajLxEkpiOZQKbp5JsisbDNFzwQwXFGvr3tesCYF55nDaAPC
gH2pqE9hvgfGOMp1Tf8kE/v5n2qqEEhvdvjZ2NTYFdFQ4RAVAnUP1xSuqIEzETp54sRT6ggs+z8D
m3h+noP1V+hbGLwjaqgGpfdOSHWURRSui171Pyv7e7YZbvdF6h0tabvmOFvvPUv3kFbWhpgHc6PK
Q5vMaWvDRRzbRkAfFbxyb4tMMyMk98uwSpsP6NVt1UtON1hTdZNnH8d8FFXIKLNRxnU5Gc8mMMpR
KX9TVFlJ+ZE7hjoC4pX/DXj3vDmOQtGJ86H9UOf1XD3zbG3ZbIbr7487Fuo2/L9zQz3RvXvL/hcM
45P0AjUonTKbu7sQg0KAUqL4k488mZudvHIwxiaO459P3H0nbVuqT341j9uDDkkz22xjDn9dkSDp
UHzaDmcqEKoH+qZWdkeI5fNTBig9ixIo2VwqVsOvryNbW/WL7rAqRFZUqfPv32PfBca017Xja7Th
VDAfX/AfOR2dldf7Otv9zjrzlxwDgyP89r2lVmOXV2V1YrcryIJiH9MvxKnRFQKHRDwydAlW9ePJ
h86bgF+uGgo419VYhQ5iKJVIZp4sHJCC/mC5Oi1dTYvFO28mtWyR3cZU74tpwMDeyJouhZdxph1o
rfTs7++ZTm3ZIJByr2ARDqxIl+YGORlc7lytN8SXFRlpOhwHFmKZG5fdwPGgzfnJRGjdNzBgHX2z
qRJW46EQi6MwIxy6eMwAqrmFsWr8M3zRWo3QeQxWASByFu5Kg5zJCI45A4lPWBM0K8sGozpwW2uB
kVznG3in0PCa3DZbIKl1gvEgnbHa9Jihzcd2H7VdsaseNmuLkH8MhhxL0Iv2Fr5rzrE2QhAKZXTR
VPgFR6RtTq5heKNR2KoQttxOFMX8wZCan+1rIUnwm/BtBDuV0zbzlKVp4NUYOLUNgmNLFdWUpnzf
7TkMTCEXTdR0f/ZOIICNDqTlO6bRO3A3dL1cpd/aNhr8o1LkBe3JVymp+F9PAQ1jYtU5TB3GvbNy
32Dln5KXBV4vxJIJ+PoYtEO4kDbHbohuYHN5w7vx1hRPQCNz4sK6MW91QcGSYSaeX1bxRiytlVZz
xgErzMzvn6wOHhMrw2ufF2qOhz+vHmeHKOlNGEQaevBoKkwGUOsU4FAdubszLFwaAN3femRxA/OR
4nDWG2/UzSA9/5j5gK6l4KbP2wCi8yevSzhiacOYmO0lweitk4Rz1Y5RQPaNIZKD9L7OXf2zSlba
RCAQI2RRxLhX/bl5H8rQMf+L6rw71jeizsKoLfMATlSihgIw4+/FjmlGVKx9AFcVuxwcodGidi/R
xLq1U97cOd6a8brMWnuaTe53+Xn8151j7Gu35LF1UUR2ynOK6k39i5glbiKYAZvds4qoah7wfK13
/Z2+hiB8MsMP8wbquhubSiiwp4er80S+t2m+4xdF0pc/zaAAuJZig8mXX8ztjckxPH2UDeq0sq7l
fyhC/zCZFpIu9tExtnfNKuzDXHclPlPEaLmGfA6FXlAxBwmeYD7wWOX5HuBU0clZZWxxFlUDP+ed
h0xVwN4hvi/rv4BeibtxNsRKBwxHxD1DKyVkDb3vvypS5ADh7d3w6w6RQIBng3K3P8KG9IGwtB8w
eIfs43fE5ysZn/uiH3AnSk2je3moDnsZ59hY7gd3fHPPia8nORidLYKRA5ztZ7mgRtm1uJwgfmFJ
dBCRFVxODiNxvJIyIFYXqLEFhYKgJ0Sz/liC4sAlkqjsx5wSYODJK34mTJoL15isH9ice5L62asy
zPnwFGGpsliSvKwb8q/siWQDFBIN8OzZPHf2M375aGUe5yPt7JZgkdkkgOiD0uR8PTKEM4OwU1xa
CPbxfArfW/I8ZPG/3LeoucOvUmH9ipxd/R2jspk6KG+pQFOfCUOigsDsbKwAY2jEfqCCcBjjKIRB
xNWXJVmqvV3n78nl1o0Vg5gHdQ+KpISnVCAvxe6ta8qLm5OqgroY5ICLznYO0QXbt27wX4tPWfj8
7a0cvwFIPbmRfw/TbUgWrj1UdAza58N/1vcGBNw8BacIfvufLhWj+eiLIBd0fhrYHO2CHdgh0eqq
o8bnsqNiZ00r/m/Qjs875ebPQqds5bbtTe04PFpP1gcfQG3AqxaGZ1spaZFw9rinPiIZuMDD4FN5
Ed0gJBDpXYinuT8ZpEgwILkD/oBys8RFAaKqEJHFl/xoDsJxSKgNCXdHuO8TMp8HSF7DN/Agbmyz
J0963KrQOza/NeKPld17xPZV9+qrXBYglUSR4tTgkH1d9O/5JMnaLM6ecrVBqgnyotZRpsKNLkfJ
9VazgfnBNakU3awtwNhtCFQElNjMfesdkxnPyo37BOeM4TcBnrBmT0rlMaHqASJW/8kfUySzACuN
xqoBHO/Ia+WtgbW0O6xuGx/Qy9Ffg0Q4fI8xZEC2xqu9vT1zCCuyMrNyxCR4cup3K8JPpGfob8+y
m7no9X90VFgiVPGZeoOneB/liypxLYtO3TtfV+rRGSLAH0sAr5k6a8pVV4TaqyYgwbtR4aGV3BxP
PGoyOOeOuzk95R+WJDWZrJyp5fD9P5RGUASLO2ksKMFsTpz07I3ds3WCrtggydq8P5iFAY2e70g5
UdV+MdNkwZ9Wu8ZpnU8zBvSJ40JSZlmGtj6jkXYEXs0eeZVo2VNPPq3jwEg+pGViciYZ7w+5S3yp
Hir+R7Njcoc9Dv3iqoYdsKdwSl5C2W0jGAKC74SiNjndmD7p7acN7shmAbpdNA6ZCIIrmmPsGFlw
ms7Z1XGJ0o+DaNZJJY5X0eG65E99AHbzyfjatXfra0Zkc7jCrK2SLt3zZR57F+SYjBlUoTWjA9Mv
VZXFLK4uViPJp5nVCvrDHKZ8b1SKCHFxACE8dngkBXQ+p2T4Z02YgwTnmI+T6B2zdJzNu+4GbdHd
i2QHH7G/W0P5uEQlarWZRHqr0jWUbJkwvryPRs3yNNE1z/5zml1OouHgcqBIehK2hjhK3l4KMCZ8
+SoROZSZCb9qq/gspZCypb4F4aK+kRed/iJqU9VWQuDJxMXzoQiFtFvuidHaKl3ef1GMXsbnPA3E
fQqrGQmDsxWZlo4m0gu15HweDicOizBTsmrZjt+r6Cht9yX0Zq12gFRIU0Vu4DJ5xS8+PtnQLeor
KDFMk4myl1Axi5Fg2nDJTlBXOD+bC/SljrvesYTq5VGrx0A+u3x7unh1STgZHiQGY4X8ulozUiWw
oFgJ9ac6C3uO6Y+ehfuEAZILUjOwZRatHESR7dE9jHmbDJfkOKoxFB2Eo7JAxTlSFpWtQTAe1l72
2Yy+vz0/nVVw8E6IU6Q613brhhxrfJK9ZOrvP3hR2vJkzDQM5EZyqA3Uyfzcau5AzId9ubd+SJXk
thi2W2b4WibI80bKVTRTVhzQ3wZjOc4lt0OHm07hrVMpQsXibXf/1WvD3O8Xj6Kzb+XdlLrhvpxq
wF4fn2GEHovLJWGZ/YnnhjKkS5O4TglIajqG/PA0n4w2TIgmF8jtS8rW6+20FtaMpTSk6W/JZfck
QPz0x0dT0yi/RaufjGPJXC1Ag5bd9L07dF32keL6V+zoN5qfm4DyDfV5VqxwbpntV15H5BlsYe6f
BIxRJkrWIuZySPartvXADtJ09t79y8wgg5IJ0MdpdosjH+Nu3BmRNhGO38iwyI6ygsXDlaBxIRd/
hEoi8KFFAAzCKCIGni4NAsrpC5ACrrd9lY/FIi2e52x2gEToGlQ3o7BxpM7r9NALqJ/zgwnn1qoC
4kNAdi+JANdsTCsGS6X70dYJzVKLjl5aw9ogJomp534EFHEwL/X5enOSugf35VM8KYrmAOuf8Svw
CGNwXh03+IB6pytB/snuifL6LcfW/7yAvJ6gmXsZheY38qjuPA/hs/4GGz8kwBDkVaCt/ppjh8u7
sakPW3izwPcSkPmzxHq3FaRY7Bh/n8IaLd9fCGu4f32StnIDTHkncFUgkzxnFdieLDApSTBVKtf4
HCiU/t57YzTPQPLXPUVVGDdmXu6DtNywItehNfmLV88JYFM+opD+Hbhm+3wmBpcyC6eHzNcm+J/q
LeAndtLDaaQOSzPYWoTFWuUM9St5lBJB+R2xZ7z8wxGAhn+KekLGS5k9ermOut4ALKQYwR6W5V9B
8s3IsG6M8zkkSOJXc/je6dKHAEInCUyfAvKmBWU48sQ57X1m8Pog3CimM1ua2RMKuHw7F+hRm0aM
BgrSKHxGmQJICjpFhQ1v2rymyzsJzNk8euzw2h+f3jHECdF85/dff9qVHhsl2B+UuQcBdzNPy00h
J0TOnjGxsGAApHTQFiV4LyUl6U5Y0w8RVje9gWNEJjjvig+E242C89PCar/IbqlQQrvtAgBlO65v
240XgrRpHTjBo8TIOaFkd1rUTtnI8QGGi9iT4C919ymTNy5ZfhRMVGcdJawHcVfJWSDFoy+PUJcC
p6bC8cPagYxI6U1V74S4jsZtO2YU5i6yXEY3fqP9R2HjzlhHpC3jJNIvio9DyYe9RZG2q3qxA/dj
ZLnz8KkXiva4eBVaoJPjwTiX1vvJTQNni4iDWer5pac7Ud6tHR4jl53CIzvOPaCiSIP1zW3Ghb8L
8XhxT7d+xC5sRy88cH06mMxAytUJszOKn/Tgw+v13srsIqkCTgiSpvB4XZLvrxv1HctqCDBic6AZ
Oj3phbgoK8MlxNbvP3ovnqSdiwg89VXIsXd8HYDibuVk8e8pxPlaAL2oNV8W/xeNo2vCCXn34MS3
3b1swPFrwXmUOeQ9ORamPVHQyE4tYADE+ulzdbke4hdOG46RAp0tLIoTtyHQNx54rhKnmODRM+6z
uA2geTmCGzSQQ0kzu2ljOHZRjW2dmEsyzdoSK6OgpAviGB31xuyYcWmONvAvlCZFX+zHQ1lj0JqP
OdmHleWSAy7khFgf/S+XgnJ3gfkJQfJkXUToMAGwGT9KK+PYvv2XhZZGHuNENXPF9iXA8WtNAndp
pPmh7c7sYq+lCxRJK9y7F52OD2rKBA+7f1XSZtSDl64CW8huPvDwsWvS+fsz37pSBH8QaZnXZDy9
yL7ReJDDsHtYfMD56eRrbcYlALFbaxba6t95ML/ymH6wSmBLJFzteAurOG6MQG7S3DNxSQNNNfe3
f2V/XCcrAO015cxmGyohybrZtjxifZcLmG/wragDmOccr7vXkl4cWkEdmzVTWH4eNkiuuVvX9EO5
PlKbFwlnruz159wbs3uGhhLWlgwps5H/xSFF7QkpV24YrO3pqnBJcED46Hel0CisiANbzwczrQp/
9y7x5X5QxzdIxbAKT1rcBc5GtuF/WFjp83xQtbiuTXNbcBTI2jAeBBZ4vjEWpEOqQ7uEY8xGV6tW
PTq4QaDZOXN2ReEn01DQ1dnSQzasor/42u+qDOV9++P0iQqCLkKMRaZjOmZx37avu0/tn8ghxIWd
YvAa3U/5MDnMmw+ykCZoOR9liSqF/2lz0qkoSHaNPAFXK5ckPmYDxPw5N55Xj4MFrx2uDL9ubZFo
wneInYDlJYIm9P91OlO5wBxefRqVAHFpNNn6d9Vpn0pOoSCXdpPBDqVvVsFmY3vQoNomx+6xex54
XIWKeXDWXXldMBQfzCOgc4wVDtj3uJ8XoxCK63wi5xNV2Xh3wOMkHscYznj1F+NLDBp89nqs/gTR
h0QMwLOF2MGdkmb9s3qJ8IleRyGAyr/4OLf9QAZXHte3ACFS++AC+uNPGMd+mn4Tnmj7pLjM8Xpo
klAiBMJ9smDkyZ1nfv0eolDrv0nk+P0gWWw+SEC/Xnq6N34d7VPVfCZ3OhKEb2vbfeCmeCa+rFN3
vIPY4dHKaAznVQhz/ulRW/4gV4owvySN6cB14bQ/WbTqEwu4JPWWyeKtA/BGe0dWYEnuHi79VeAI
olDPsPO1qwdMuDg1wgH9OnUJ18D+ol6+KxYiV17WxgByQoUi9Z6q0HDd35D65P4szgFs7nfbk+Uv
Yb7eV6e9FaS79wG4HPnZtioD/cbNnBfg52h2GGa8kNnTWCZhVAxwpCeszL8jFOJNLjzsZCcVyV1Z
7OCCr1ZMNYUF4lFWYzEbVgR7abyiUEu1b1HsK4shIXuo+nLyadLlyaLXUt/cChzCJEsPUEd034A1
BJSpstTH65EMaGEVouQGlmheAD2t1WRSkMG3/nt8FiRctJoBXkWWJvYzlWS9EYeXkx4U0sn2y4qZ
pm5hH/QR1lsPqOwagZs9/sRk6uhvyh92q5WGf3kpM4gj2/3teMd6Hq3u3o3NV9t8sCZuFEe0MY6P
TxQgWR+Dgr8L+uqzOCuVx8+OQ4FxGYV7bEVrPtAEZyloRq2cvIB9sx68LXuAc8PltlgyQrFOFQLp
JpCaTmF1Pf1wlG//56HhtnL2jPVrxbuxyjN3186e0CI5jNZMCOoBnkmLIXUmzDrHPYEAjih9g+Hw
WmoiyXZl0FaJmjf3uJ+Mk4kzyeWxO2oejvmaus2zX5lw9nwZeORdXa3gwfDuYqTJeX4cB8L6gzjl
LqDZbC2iks78BAXz2yjTvW8xeUFKQo/PCsBi5dGXd14LO69vUkZjYxCGrrchI9vvjeBBog4iXhRo
5YMfmoxzo+zxHDWrNvSXgOn/IAAX9ymQfS9UD9rqLTko3LEE02CIONiutDg17juuNUK1YIJkBg0c
SeILNSjrIoM+c9cizuEw62gkYf5ZYxWYBJb1Ihdgx8Wd6EbdNHVXtnNrd7UVLVAqKsfN8j9jAphZ
YR0ABvuuYITF7DrJFpuZNDDMk8yhxaMT/Czq8i53qepqfq0ARU9j4yr2Temyf0wNAxnLUaFWks/r
ONdo6pk7zgH0hzoJsAPk4qvvINqKCFBcODzbWWZy53MSQmVWWfruuLJX8tMAbZoqdTMsiZXHmc1x
/2nt7rrB4xqPzNvrvGPTt6z/8zJJFhRF7No9RAVVs32qaJc4wkZVysYcxTECNffs1Tat3f7JjyqJ
9IwXTvU4Olb9UkZ6bcYxUrBPYO7EPzan8EfzDooF+4OQNf32bfQbIehqQ8pJ+aJGrq8FplXgOHQz
rYFqHBebo5eR5NlVYJ4h2dhrquP7X3zP9vhuYLKza6HOq1ZPGOQUh964fGsgwyrG4HrlfNq9KT6Q
cL5xDRinYxrYnjJAHIwhIivZxBoc9R4JCP1Q8t4fMFgltJvNb5OaMVURQ2EKuGcUHX88DYnU/NCZ
frTIwAx3gwqvdMa1XaVu+SqApcEvWZOubQXb0wsUElyvvcl9YYF2XC4uYbL0jTparKDdUEmnZT0G
Kd/gW3qD9IRW5FJkAbu+Y5TIvsbMsMZbzpS5GcuANPcGWUKaW7Qayi0WmSkaoqAh8c3dTTECJKNs
zKeR3qBsymAbW0AquK56FWXWX8ym7v5tMl3qSPapZG6UBrwQZ8nH3vGLZvoVMfFV/vFNxYLhAJsJ
mpR3HYSWJRmfd8qrg8SimQBY/tY+yFH9K8sEbEggC0CpqKS8j6O/z/wEbboQQclYTzS/WxrUu7nq
rRHvHR8c4UPuHuxkXA5mI6+tP8jVwkKRgIcyuWLKHBnzzJ1NFHOcgDJB5EA8+q/lc7fUjIVmgIZP
4Hpru/ZHTIeoV7SJ5Xn+aP35RN6LzucsaHDpbdSMtErS6fB0G/Fks9xWH4RGPmW6AxGtWmPvAARH
vOHMLnp8RNHwbsq1VbxWIk15FfCbQkhvyLEj7BUMi2Y9K/j8b1xKzVV2ndDDH2RVIVNOm8Pq/35Q
tiHEb1oy/Vl8uBLe5vHAu2xCGkdoOzvvxpcCYHC5pZUPIDnmqlYjmqm6tYtd+XIvnQ6cgApa57+z
UKbxsoXGlI383F9ZOHx+lYmzY9o2LiHzUEpJ2VVaoD+cL7+pmPcr32Hdxs/oBtIf19Sx9KaNIPI4
GL+IUy/suGQb0zbcc94tRP1bVZTYyx11pRB2yinkCbvoJUxN9KlzvsCHz/oAdMTt3W4p6Drlg5BT
zLVociQZGssD2/ep4ElOSPZKgb5LhvQLRuSrkmbRcaYjKY1+ENT23EHBGODWfoyplgpINGLiyWKI
/MSL8eiF0cEUbDiXvDfBxErNZ+jomLQiZxsDzceJRgdU0mAFcPFKfDjMvLkFstjZfIRFQxKtiiYH
UcTeO5Bs4ibRByghH03OmhfywzV4EQQ5HxKzJ1QrRHGW5nZyE8ZjA8kFJRttDE12GokG+ZYxgY0f
oNUOtd7UVXLS+F9YEJ0cXD1YJSixa/4pBeo3RF9EznYaC4t9YfP5I/qmMpNP4TBwwDS2PLoExquk
bdZL0rw7FbtNJ1tfgviWc4TUz4J+mV95wevUMAe8D7eFjwPKwIsDiAoBeHIc4NLbsGuBOa4K6zMY
l9iZCT7BTWgWfwjIZhlMhgq57JH0/X4vszugG8R9GkCSL9c2wBKy55QpBakNCHXRWnSxqTUZm0ro
69hDOJ1HifIjmyT+eWsoQZgIhBEcp+BiFqA7PDZSNDq22PrEY6GmLwNcorNLhpWcP5NMxLhNRVvj
AV92Bsawfv+DrmNqbg86TxZwSCt+lyXGcCRP0r/zC3ff1chqAFMi1uVyO/A8V+3JrP925puzBN7S
2uDlerBaPMn0GCs86jUpwCP4cibNFaVBgZO1lkDd662yU6JjLkpgBsVZQxnPdFvUkmxw5d4pxLQY
yxnr+QCX7RIXS7U4Kvy81ysM3tM2hPthHaxXEGWDDhHs5C8WILtGrJWsPgDR5X0cieo14q8KND8+
ui8HdziBW//HU2TdxKpTRr1nEsExLw03fa/YnozL0oe33W14xfMJLUWzr2aECJDa66N8FGUJqJz2
vAeW5cqywa+mp693ZOypX8CvqoCgEr01RazJySrgZ422BdN/eHNeya75O8eZywGVSgdZvSK4ES9Y
Xit8Hvu0NHDYdLz4Te+48EhYXJ8MHjxhKAszAyUJGSBZqPRgqH/GqEOjL9V8HXCpQWAdH9/grwMs
yDKgrW6lEygfIEQOacdrgqqTYEd6lMxKv1Ccc2yZ1CqigdSueHjsyb1HNi6LNiFwJ4SzvL3u6u03
9UIjFTCh7Bb1M5jtR/tGooOzD3LGbA3Vsqa+ZActnBhD4sB8iqtEuwGYWYJErymObcfkMrNNEPAD
2xVqyvYq3Jcne2xRZyTmkJMpYygQy4hSyX/FbohD+zMgI0LGs8d0M9T+IUq7WxX5IaxYiU77Og2X
11Mv5d9dME/5Fcck/rpiImG680h5nE7DeN+N3vdNtXrtawHpCT1K1kfftBQMRtISqc+9UrnaKcIm
LDkIXyL6VPKg5onJWwlitJJSprmHUZh2Qhrhmq0VO/OjguzWf45dqHkxsnBFtE9ojKcAZPWBIVY2
80jWws6wVz20SZmAy/syVP+u7rn6unW5fJMuUrbyoXyCuHmOAH8R+GwF4mY4gM4zPjVfzSQf7y7W
Zkf8UkiF5E6cIKUQ+iuskLoQKE4/f/uy324RweEWcUKb+AirO/DdhRkaDtD2vSSSjZ4WSKJpu6Zx
vC/P5cCJ0FDKMjnDiEoyhTHf6ZVVZ1v8nJYl8zvhrB1Sr9OI8oJcs3tkLhJbliFPy1q2th0kX45D
RFDBI3rPKSGyA3scF9DClxPSv9z2uwDr7ty5EcOf/6VoHk21edyW2qRPtOQGv41gYwXPBt/pzZar
ajIR05TwDXI1zbe7pi7P6VapWmcAb4E9EsrMl+Vi3FuN16AsGvHQjJR+KZSKB8zti6KGEcH2r0b6
YVArHsd8ZAXTLwBTIZ5NjmMzTUOp13UCVlVeZf/kNZXLz6Fg0S1AEt7GB+SD4l2M3XIdm8TnLyU3
fEdJRtrjKOxeYA8aGwZOhHhECSKzxHvdCHHR7K6ffblpcp/zsXpveeQg5DPE+vHCKXedG1OzOpQH
oAz4zMgwtOv6WUaR0vDmhA3eJ+3gcyw2G3IKeBGs45pcPjT6NVq7QydvWZ6D/7EbwkBoUjMcyVfu
vvudQPkA+Ms/Y1W1stLWz+0Swcwe/a4b9Al0PMCunKzYv36VYKtLNUu/iSNmlEMcaF5SUtRe+O90
0hnM5y04ac6IqfC0sVF3qmA0esyWZ0TatlAYafpvpfpJKs8zrFFymk1oTxzF83w7HrhtCfAdD8pP
7ShiQii7S6pTmqXXo5ChaX2/RYbk9Mf9lj+X10tu9z8G75WUoOQsng0eBnW89aa5XT468Js93WCn
nu24yXhQuoodoolTmS5SQpmMJyc22ZhPlYHraICoQ8Ck+jCiQXARmwzbgneNjKF7EKDW6xDfJ+nl
PJPxfpPW5okmRIW9m8i3uqdbGDt4KwwoNb2/L7S2WVz1KmOlkmltPKBZhBrqkL6qSMgSMqLXvBg8
K/qiV5nb0YOHDB9P6xbWd4VW6cID96+YvPDDiCzkuB25V+BmA2Od1QuCJNwnzyh7EIBZVn4ASNbG
/7QlZZcNfjyKsgOy5MENtPARysj/sU0wvjxMBpTyY/PqDhnnQY4ZtYVe+4QxRDMNpRmBqInyqajL
5vXsddj5Wy7hBy1qvfnxig4GALhQr6IFLEj/8gM62/ZS17hRAQiayOQABRI/OUlWjzv/1lrdX18R
ifD8af5irfbuhgLK51kaDKntTFqbBunMjz5QAOVbREDPwRqQM2YLhkl7mXSbw8Di//hjIZhPW6ef
5P38V+NnJdDNFnf602BMkIDuUrtrF/vuu6mClOjBPVXssJ75UzX1CnEkQ4diy1rXJ0uma4Ad91Hj
ZkvWgFl4s1A+HIG11+F6bcAYjV1dqKzUf7rU6D10uhQsjbJqn7OxUwky2yslJFli8MLIuPN0PjMJ
Zy0e6KTdHFYaV1pg0M8mwA9SK18SOHXZudFYuYGxQJSs82VDSfl+ffDz0Gm4YF1akRoTatU2250o
xvU1JnCGO6pAh+e7ITvQbN3IRFIaL7wtsRKnhLVcEmFgiX1IUf2m4cBO9mNsH/ITiGHN8FIGCSi2
PkU4Qi2ORj0L5kNuucOCI3LWyScy5Rd3BXyqS6j2eTlCPBfPHR46KQ6zsH2IkeKGvKbiksGRyart
WKduZRXuFGr02YMKajtDcgVSYdoeU4Qm6tcfyF+PO7qNEmT+OezdWzGw2aSNAsikcR15HP5kFGKD
7oRHpnGYfFW9RMzNg4p2u2SJT4rlfCJxK+djE+ZaAeCTNn2N9yyic9f6u15yXg3jVotoLsUe8Ql1
GcUji/SwYBiIVDybtYBJVxdsxerZ2jhyR4J1Vi0GOVoaOwOfai7u4dE+7yG9JWaR7dEvs/9m7BNO
GFJnyujRF/ckWmFk4t9v6GfO61B+GFIzmrNtZqaKDmqzxGGXeBCO4/eTSxeractMYG5vqwAY6mwU
wKrTo9DGFg2wBu3nDSvRlMkdHW4G9ZtovEe6O/DPEWMzqQv4ystPAYJlQYTvC8oeZ1wRGEtaVkp1
QHnzUbPuJf62zLblsmXhUacL2L6jauhPGpY4kvPqRzcP9L76ZvnyIE0bSs2FGRhj5+f10WBsjIg7
0OXsIL9y36k2KL3FiwuaCVA7wUbvlm3O3rfB3aTrawg2us/R4hQXfKY2VNLpnw9wU+KxU8UhIl0h
WAfSv/kwUVwcMC+o3LNGY1LPDD6pywl9EisBGis0U5Lo4OIaqEXjTQc+6SJh2LgGWwIx9/7WWaG/
CFoEriH69VuVofiqXi86Ahq8QNxHF4EK51nm2jzWAGN/mM/hAnCTyVLqzzxyUq5o626FS8Gk7yBu
jNHS1K59SHpkJxj7CnmmDw8hsBYB94jwfboyL9/AEoSlMm42TySRaAo4EaDp49RQindt/29qyJP7
O/Z8sWVFWbY1Ra5JmbIHlEj+2lvqo5JDzgfY9GJTHQUS2sKVqAoXdGvRInbjrke7UZPbfuNXud75
1nFw2GidA4ZCFwjGhAJ8+0pD2dADrUX9D30r95WPXpYfokWmeLMFm18vhVObBgzod1gRAFerJqEj
jB09smJXQJfUFzw3Po/wrEmPmL82wAbKV5lDXZEeQ2XjZ2M0tm5gstonoNTkDfH4R5lDIE9qVVXs
g/b6iNok/hSyi2RUyRyFVJrFWFEdHH82Wouz6MoOplLpYNHkSXmMssMtTDvt/bCk7PxlGQFOWePd
pQaQfvzw8y+u5ZcLgtdXfFLRscXQOVKjF/YH7RUugzGC00yyOfZ0kQ4VWo5YTrOcNGECUgOBtt07
Nq61HB6XMC3ZzmlCbU7VS/JOVW/usRcq4J2va2lFpM33/HcNwAmIkiTC+TKvRQ6q8iR8if362nJe
FNN4i+syAj4p2c84+mI9jWEptGMce5HEBjoG9MEwIgHerobKwm8O62dmO0j9qEESGxXrL4G58SWg
zLQy6ZiweqwO4+2eY97jFJcS4GVmwkKpidVkG5p73lX6eyRYJlGp/iVJtQbaL9J/ezNkJyuYCIYn
QLtueELU+DABb0LSBaL8VtggDSZy2y1sl5HDNC5Cx2m/SjWui4GEPE9drYWrCN9bkI6+srjqxShN
bdmCE5mebm0d2nUbQzJqzfK5+NbRdrm+PFU/5zcWS1ROZ0z+nL1lIpKDLaREHiJOkkih5EghitxW
yFII2ZwHyOBm6OaB+nxrtbmEvgfAiSsd83KWYWBdFQMsZmFvs5BPl+4KwwUZabblMMKm0ybyIJ+L
4WbnyMPL9uHLbPGN5ZspInmNACHdrTiH/y0k05poSnpovqimlFAb1wGVNZcLPvcAamcP+dX5N/FU
6EmyNpAOeTAxhB2HSy8tlhVKPYhCiuptXZcXB1WFr+iWUj0mLOgZdfugciOxzHkacGMXtC/MHGct
JNBQ7yMCut3WLdUE5MeDN82gGu+CQs65hcvF1bL6n93+4zbu4DvnY49T0a0NeV7vzD4fi3H1daIT
/KC3UWV/Jb1/2KL9So8L+/WMV50EzwZcLP9yX4q4wDbUlISZBPP2kocV4hArdbhR6kr+Ta+urCqa
nvSRxJXCMv4vij+qw/La+bd81zrnIQPuaGs+N6QFgyAi7d+iUl4w7vUBd25NpR27whLNjeK8omwy
2wLvblTvHGdAP9BAnM+PCl5VBfp/cCNSeNXax6BIT4II9mg6DPTBmAOVOndMyUum8JaINYIm5Pxd
Qp8eOZtQbswOnT+SHeMXAZfSngqTFukcSS50kUJJS4zvYYlfihu680oUuUnclfa1YFoRSjPBGXfw
fh6/FpH3BT4O0/Fz1ibn6l9BgTHlHv1Nq3PMLK6P5yNE2XTRyR1VGUCofc8J+R5HHLCvzu79u3xm
GqKEmwW1egUEul8aA0xk6UYIXiwqq62Apb9P4KvDURzJYvF1d+Q2AYUnjioKyRkTVFfUrqLBDk2L
Le2DjubJaFZf3pzyrPg2z+6lHADwbOGW1NSJPqzaz0eXoGRL5JjRJLfjJ7+/6LnQ1hYOm6KuWflK
/lfuTWu8MQdM/Uyc4FK5QxMFoIyFCEtwNPJvX3FnyOA0wqHzaVw4nChDqWCv+bwiUQK7+LKFx84D
ZrrFecoMd1NvtFZJPfFv+U+WR10DAcLfZnceM85TajCwSiUvSDfYi9iIYiamebyON1abWYKRETY5
owA4KXvG0zcMBUo8ZYUkYEnmMXegTJzfnb7aLdLEaYyKT1EgjW2hHS4HSSrsoTGx18vdCZqnidKd
2EpN0TWBfYe2JvC3e48XLqfo2Zb7YOLnJjDIxjXnd0G/0f0OyLw130quZ4r0/nSbx26xUl0SFc0C
NHfz/ZxWKQ59hLZNcMha5TmS7DN9Q3c8iMuGVcP6qPRNRAV8BcJ9wANfqKuyzIGoR8KMVougbRAO
ksyiAo/Iup+S51Z+mPdHKfDgRCBPmy1R2z5ZsaNDxYb4bqtnA/6sX78LeXe+qE5AIi53w4Wr0soh
MyfD4l4Ksb/7Tg1wDsvsfhjEHxPWiMncIMr22GJSAwfkFJH20hzVcF4fCUEKpDFEi1oKv5MwRGtk
qWfPfXzapEwHEHLX4xSoucvzrhaClKfnBrJG4EiuG10kbj7jBrZCO2EWKqjkL//TZ2fw+YBpWkv8
V1pRLYX9On7TcovSYPZKi/Axuc9EUkHtK9w88uwA1oZjRIqbeCDjaJCd9axR8Hh2yPDO/KkuYlG0
vL3TwnRRkOd/5Fa6szQVZycOBSrmc73vSNdqr33qSJhYeZWszPB68PytrD+e3uFET/aL5tAJYCUA
eJzyk6SyfmYBPbp6ZwydP8b8w2ysmzVp/oPblYX1EcjHNLOaQjCY6/g7Vlb0CxQYq4scHehwaoDf
ZBB2eFD3SOt+Y8rddVHnwejPX3U0INBvAEXPQDT1zJimubUOv5G3WZv40TDX8vSGt1eS0t7rMsEo
Urugs/AhSlBSARJ/MdFvLlNY3Puhz1M2zhMs+pyeGkPnCiU2G5BaGS7FO8YT+u29snOMNpXnTw7/
CNVK/Xn1ui14wbJAcptT1oOD1dSjvo2T4IVPaxoxXQyQoWKRke1YUIP53WES7ZubujLTpRbQqX+g
Mh653CKe7s2k5QtzTUyjXn+Pp/iJyEzud64h5KWZK8nrRWJvd6xV2HYtWboiso6F5jfA7nfIHHCS
2o/+ORaTq4Xchv+FyjSAJJkR2nt9dDj7jpPotD6ihRnNC1zslnfCUXWTWf9ptfPhrjOcyaDTBkLC
6b/5XcNfUIEhY0EMay2U05p1my8xv01KSbvZjS1NTONkWH1KOU2uuy9g0hInANvF6KLT9uh1Sv3C
VOaS78JXITa46AfEd9RFX4nJ28xe3RGIsLGkyq9mlJU1P3E8G2bx0K6M1iVrzSSWS9ruCfmEOxDZ
WgrY74UqVvd970LVWxdzIDGw5cFdq0s7LxlzLTBHtIm5aEMM6vGAj7cn5kln5xRVd8RNp7BWAuOV
TtO8bV3mQrNEpre7xFl8YDNmYXHR/qEw/HGz4DYSq1XQYjnCBAdPfHS9XFggIzqQw+7JtIidrjCx
q9LHTLCh16KH1Mj/XDHCmZU1WYnR+9401zMJ/8iVURo9cn4uefOhYRLGoCDi5lM3nUM2RZUnD2Ic
fUohqmgkulx8iGJNk0ji8lpWSHoyLnZc9QtAbdTEof8mdCU9idQTgtIyntENmCMnuwCKAWgU//nR
nhsigJZqvGKHupd24n2buW3Soop37LIbS7W9a8RWWUPasvkLnkUBREN4v7eWuYm1GlXTjbvZZXDl
TCGxBzyYegACTkDVPk6MRryycju/7M3+KdzVthUcJzx66bAbcl2DjpWnxpR5NzRhMggB4gfDs9LS
tJDcYHLbJ+1ddnGRBNCpZwVpII8F7VBcFNCHhhOTC+yyS7LyyEhav80WWXTelojfX62cmUOIN+EL
tNO6y4y1AGtNxWlYcmhrHDHcE1QqqItOn/LnXMoKC/1hSOodPK9tpQb7sFowbRXqk5Zi5YFeQL1P
ozkS1nzIAosIYObhTKB2WGkjp3UUv6C9f75KZm25JNgIKfCOZN/BTpC2YuAnLPUwiNKVGZ6NYR7S
UJWUGyiDpZ+/wSdgtgCAvUjdVZAszavbvzVODYesF+bzvXyMAbha8DOxTRkfxbpznSyTosRfJekm
iqrEf01cL0MENKqrL5YxUUIzTJ3aO6nNv3mzyXgMGWoRxhio9IR2jOT50pjIMbt7Shy3EP3fQ/49
dLtFBKHP+2m7PDwePEl7pbipWQmpzxfWrRfoMk/+lWC70CTcHv3C60e8rUr7u5VVMs0avUIMY2ud
iwT5zldWChJiGAKJZUu9c6f+tbX/BMMW7Quk9cI6XeHWeXEEpmU6oIQ2ewDsHUL9KEPwW5XdGoLE
vP6+f2koJ62oLr0qvGOTmhfWrR1NY9SCnEYVrsDbV5cI9oUPawsUg//X4NCTDG+crZr3vtJB8GwY
gYtHN2JAgb+imjC5YeKZvZdrIs8CSw2qyM1NWyFjXRACajvP6M/EApOaX5imED0e65qneP92w/nw
E9vJatQngnikF9NJ4QJR4WwiSlVBytRqXhPBd8vLj/T9290Iz3+ZsQZMXhZDpqISIsofbehAREvz
D+8EXiii2vPRX8jeptu5x9CRCMLPOFFo5Pv8ntnpwyqA90MuVmSnhImXS40kCpLIyM5qaNdYt5r3
pOgqlBIUT5PEdOA3wBCm9av6QdX+MlOoeT7OIzx1ggu3fiYZP5AvecjFagJKTNO402mubU21bdGW
vWhQDq+e7tRHEPLD0GsXGs9mXVrJt9XfEYi9WCztI34NXYK6wmclqGE0McEPjsz3BwctgSGowvq4
H42cMaRg8Vg7X3ktlWU9bwBnysPUZFscdWpahQebq+DCu+Gn6hwR+HS+HeCToJKhWH9bz57N8Dhh
Pa8dKRAIIFOGgI/Gkp0aKPIsHiHn50pE9cuqyjMKYFKE/n5uTYGZPYpn7zHYH66PcvP87+dhgXLy
JO9Ei6SJ05AWMK3w8iCnpZ8vlMWg7LzmBQRoN1cAR8s1mtyW6lcIkrR0yfUZdUbaCHQ6U+oK0+ta
jq+tlRQTXhMfT70O02oT11hfZZnZ9G6LaJa6iMCKSibxjd9LtpHFuT/vRwSuJJekzBwSSiGprKpi
92Ic4FEYhsr/7nHHkYtNc7sDBonzi5X4pPT6HICSX9oKsCZvFpNqwYH2otbol9z6wiciqdjeaklQ
fXAnYkUS2TvAHVAonTPb2zivcvddmzloNOC5Xq46LiLqStbXuj7cJEAIfyRkZMj64ZaViO84rDmx
ERSxXiLPXEj3HxdsdYzVEmTNQXXd4tKN6pl7uUxWtJSbT9A/ZtDhIffqP+EuggeqF8dYLw0ptEDV
in/dzvleSOMW1czW8tLJKpvvRI+ziObHfwLBvkyUU0otd2rue5JIqhqFI6Ot3/eYnR/vpXaSkijb
NXPuFh+BMcDudW1d43+mN56S1atQhJXTwC1TZOTMljEO70ks1vzaB5y+oJWJEXJFOM2qi7PW80nF
M6nU6I+BRA5EGuDyREd8J99msLh9HTkjPAtHcci3shn1UOINbH/FCOtAsDWyzxjPbjgY043Dkq6k
tmDEFdjRi7ZNalM9Ai2EayOfM9DbqqUIYznJbFwSZhtZMg6U1ehXWNqsFopjqXgO/jXWiGhlnLtM
GVD1al2hjediOoIL4REVLTrDwISIqVYax6LY02xsGMwaMyNIwhDayLCg2FCF2UVZviqLaSdjxraF
mzgNHbxYR5k+4d53upj6GUs/0upGASaBYniCjm4HGxBpP136Fc+s5CFoR/6DeA832wB8ESG/7IYM
WJ5EVCtcLcXMtfEi9MRFHTEt5x8hrXny/dHdLDncZuVyXbozN/U/+QtmWs3jWjrrsaAqKadcTCYZ
LGYx6O4lvhNP225NhV1U9avAQJBSfjW+qF57O43QyzEk4mQxRKdcgi9AL2Z4vaKOKQ9BrQDLal6V
kKZWn4pljU6neIYUZjfun0rqi6xwEPFpE/sPJ58A1X/P1T9Es4b0sSeHPgyD8ey2MUPYyjbB6zlw
6cDe15kwBPfg+ncdJRPoyw4DercFPaF15UgY8XY0Lq1FBeOp89zB69yNq3btZkWF2OXqBcwwvXwF
IoqQSP6ow2m6B+uRttBs931pqsRfXMsiERbzJcoNp0jGjAXGIuVoGWOVkQ1BA0ly1VEHURP0nIbV
qpO8xrqLhi5k78qVCvjDsQpKtDvib5tZ7qf/J6xkQ9JYdqn1GAm+DQSDfZnHryu0Km4fI5wsq2Dz
UUmBM5fGt0pyLWy6U4nKqG6UCSfUmL3UQHoko/qHiDtp2c1NbqjNmAA8Q9pu62BUCXBqTSMTuuCc
IavZTIhqufmsD2IlzQCK65dRoRFzwchnDRaDMSpTmuslLrv9NchO0gj6RgJu4Ishc616zLhv5EH5
FPH3PYlMSHzFqqijMtQ9CdEu+iyyf+ciKGwCYDiuQmVSR80XpchQa/MPed7WwPJ47Uh53fBfuS2g
JKyjtsFucQmyNSjx7JvSXCgWS1qFqUSj1oK+SZCPNHILS8ZDNbb+mmIg9U++9wo0RdBafAVFMd48
rLStfk5maZQJTjTBkRm3BTfAEm0iOGc7ZMmTr87t1xaDRWwkNZa7JS6TobeYHo8zuikfNpYQ1M/Q
FMIoYeBKLcf/dH08pi3TMP8YrfS70y//0ME1mpw/Vjwz0l0ry4MRsp/iVtaov3EE7Rky6E9izcze
3ORpxUpw6ihzzXWaIdDHtwzs1L7J0BgO7UOSUg0qXLkWqkUwkbvFUQXYo0lhb1W9jLflLCI7brhm
0zYUh565DsKI3Z9tTlE3jpmaoc0uQ1s16taOlyNbkMsp9u2aWAxuyC4yIVyof4YBcA940MlCRsQW
3rtTp8c2L2G7iuznSgET6VMwsg4ApGFFqdzlhmtFPN0JWyKFmcpzrOUvlGOWjstzVqfRTt3u5lWo
pwuKxJ9U9GWUOjMA/RX57dpMFzR4VJ4X8lfA5UQ79D7+JhQLpPLxnbUZe4szAocPNJClwT63X8gS
PnznepYkF1qYPxsIzmggcLdiGRvUUmXiP4zYb5OIbTfcrV52joPUUwWQaImOwnxUMh4qmo2ww6LM
80DSC5KhJm8TvsIx6L5v4TFydA04vGYfEGJL8TvekhfcGYAgatn+rZyvwKcY7xZTLu+BD3j6UM18
c0chm7TSvwf/0oc482mYMrUEdrWfNz81YmWrfWHw80ZkyXU4QDj+S+9Brr6x85gQm0rMiHQVgWQe
MZiEdo4stO/PLanT71IaosiY6oagJcI5gpRLDVCR0N2LvFJpNxZcjr+vFXZbGyLF+BvfRInQknV+
nUaJCgEMBd+6PVVgA87u7GeX22R5gOrA0qY6siGE4aKQyOK/G+CP+mVHnERs9tRbq04MPPId4acH
rYSK8ScB6t52+mPcHzFWjgUYcnlWkZrB3ydA2DnOP3bULlUiE5E69+zFjrrag0MUuLDW/MvI4aFU
NdtMCaYSxCON80bpjW9Z+q/Yaj0PKz8W7LDCdSKRojfQhMoqPFXJ9WuMA3hwNoZZGntb64sqogyg
rAKUKKdDNWuFoX74xanGc0GByJPLHz5FvsoPmkcStVKjZ0o4YgHakshqOKDGepsYQXmbL7MrQmrI
7C0LLMgYeGwpfJxVLSX5ie1C9rCqUz8GLFMzxPRDcy8pWW5de/23aQoQMiNT6jkzZbzSKi1+opOZ
2fipFHkIJ7Blxsspb7xyHjx7dNkKuCiunEKQtpF8CZYXFkt6/Vvudv31v/it5PynTiuBmuSI/GeK
z6fV0o0oQRpdvYwN/262WzusC4bHno/nWYoYAfGTYYIRKIxdyDrXjHTDfNUUj3sECXnNugAEp4Jt
mZot6+QdBRuE7c7Co1ML3noC69DVkpRRB1/FvEZ7VJdvmhEh4Q5wW76tPRJvdSd9FKJqmo1LYs/i
VhQlm3WSdZxfyWeU1yTqn9fxgIaLE2gsQCV9heNdB/82Ii+TBtLKBfl4EYF8a0ApzzqStuw/AJT1
TCPDjf/xxpeR+Hnd5wWpUpWpMaD2jdopNy8mplZn+joT7/ORIKyVSK0DmjuhNP7QbpFzcHboDXDW
UAYgNR19yLmHjOJkGbUDMpqzsZkUCSmaIHfbpsw+h7XqiPpIMcVbb+0/lAzW4Uq3HK+Ri6QmPOvP
lSkTJ8QxlmQsE/f9LGscPveaJ8yjv2R7Yxf0QRWaJpLQbuzJafPP+ioqrweqixHcmcy8kF8EQQ73
EPvmbFE/DA/oPjam+inkX/dY4heGdDNel5JQhY08iUNdvCW/0I0XzN/O3mZd7K2len/NluImDuwi
P9o8PH8u3J6M3hi1I++evOKBJYqTz08YdJRWSL7SnIRJUakJdqQrW3B72C6Ktej+lHVx8+cquWaB
EUECjflui8Cyp1jAAdlLCkEOQ6gDqtyJ1HXJ5cod/DUv+mkK5DTLd+5mh2jisyz/JMGuitKpWhUa
GwyYSFmTAsdk9+3gNS2Urjb+9RdkesD+SqGS5u6AepaJA0H6t0SpmFMewffqHTFUZWqO/h0u60LB
vB9IzgDezPni4E/vj9lJR/pBFCzAE+1OMtjdItG/OQlunkJK2C/Id0qcurcw8JQ+7VSRtghitUTY
QLWyOY88vvaRjrsnkjHv6JsarVr2wf0V66y61o64wx/raJC//rYP+tOJXDdOjgIilXmbrGCeIzil
b8gdcK9MKNuPvaDDxLH2hP7zSaZx6ruUCXrhrFeABvHMwNi2+375r1rv+lHX1jToN143HnPze3RE
yzWHwfnc6De9KJPqKeEyRnRQNmMtiTCPlOjVop6Zvobao14mkSOaCpvDRIgjnSai1QKkD8boV6cz
w54MMyncTj3RrPJLYuRtzV3rV7Vlo0MteNUrRo77Why8qZV6pOYvy1J+dTAAQTl9kc8XMwSSP1Bo
k3yju7k28/RS6MZZNpC9MP/OX7KHveXNjZwKHZto54NMce01/4nnI6tmrGoPKvtoYDvTIJxjizB1
upBwT2q55Kjh/asJRadCb88OpaLw9tp6YLieOvM+Q4NiQCXohssxnfWuxRZWCiajf++ODpWOyW83
u1bhL2ZpmNeLXnAoOZtR2eCRy3EOdcurqNi1LpT557c8ocVhAEQIYv/lSWY3YdpFhjXwEWnQip3A
z2JuJRRWt97gDSWycFN1rWj6Yi55QgmtCWJ9saer+I4+GQeAPhB26RXE2e2mu+PgodPct0D10cNL
wKEDjoDFYK8j+cm4ODmsnumHh7tBygNzMf4tci5tJilXAfWh0vnM5+NHMqZ0HYBQe78Yea7p1ywt
bdBcVbuIa3Gk2dz8wuwH5crKVYUnHVVFmeW+p5uIsiw9qt5KJhl9B4JMaWW/gJdBFf3kNMKnW8E8
oACoxnQgZWmaway9BTRCvwldRlLOIh9bRqKTHzfQigxVJ1/dbr2ZzLfaVncp+WC/PohL+lYgTNBu
sxDXwEDs5/rDf1GGClQ4fq3qhWumEyytXnizZ+COinprlCqYk/WtDTXdnQYVTitqc6JJwAYO9z6P
KjebvUYI2MizHl3OEimu6c3YMcMHNLlogzf3R4mbnxTXf8zuIdotFL/aOOEHhQHuZFQGoU1BaNgc
PwrMhwGpu1mMwXUx/dAAa1hfRKggKkq/T1hzTAZMoj+D/pv0m2FLm/mqaoIbJQG4/mpT4opq1exl
q1xhTI9UUOJZUAokc1IzpAqI7lmW5am4duPIfrzgiPCkrMNJCEa/+lMI2k4V3+hKsSdBTiBW5TnL
RZ2uBiwNhf7o0bhTUxXNMcAgXRM6aeer4+UX48/U3GhhmpniIT+MrTy0j5sJWdLsJFenqqP7zYJM
iSVppaABR7xG7RvqGLOYTktkqkvUfQUGEpayAZiPvT6GuWv5AS1llg8aCwmLBK5vKCgn7ZbjRgxF
0poywOIX6wx5Ejzm9WF+Um6gBjU5G5QaUF/OQsxZwOsftQZ5OdMxkiLazifEGKkfEgv+ztAGwXMh
b6wkTWjkIfv+gsp/v/d9l+U6ho8kHlJn5aFjLQaXsFnYrp08vsCysRjM0gJ8L5UsEn84FbDHQBKa
VLUIb/2GqxbPsjVsoO0lli1x1ficQEavgGTxQ87hQVOkFCbjNFOTMD3XZZotizIhwHL+KThkSprH
jYuBaeN56PdHCcA6yQi20+dDEPIqROEEMa46kjLevUUVNDBDvoKlCPbj4df4vB3CveIHMbsl4k/i
q2HJk5DLgVGgCkmTfu1evsNFJXibJJGtYpRYgCFmEKmB5uWnwQtaTynSHYlG/Uv27oqEfi1K756N
dkfGNSYxdDEqMBb8j5UOGRqTcRojaMpfOPJjQemds1x+xSGA2LcD9zMnrP+IgnjTbFxxOMGTO9yw
ZCnzuZ+lxRO6Qh7+LUcrro263NTTV5AkaJ0E+omK9yi98OZjDp5WmVSZUIg1jxcQYhrzMY6HOmn/
Yb3bD2fylFO9DZxcYu4ToSi3RskwP/ukFK+Iwa1khAXgYOFtxRGZt+740Zvx8xEO3G9OOSWMN/uk
9nr8uq0zU1lhSYtHEy1SpM0C0zKh/T9yKePV1YT+n41mQrV9EJFV9QJss+Xi1tKMcVcLTC+jZjSg
FPq/DsyYlYaf/PE8jBex25D1eUVIyp9WhCbor0x9Lye/NUNfqXUNEM9yFFgEdKNkuQNS7lLDk9WC
0KQda4h1EVLwIva66JtHnUg8M/vfSnNMaffQlF97dFRI5T+99BQNk0JxFezXm6pyi66/GRWFeOGf
jSltW3YB7SqldJfr+ResuEpQRAsdxH6NYUe5Els7Q7HrbBFtd8SJpXi87yhl5FpzbS58nwooCcJZ
xLapQHZzMcOCCYjk4y9NWtTeKaprkpN/pzVLrn3Ik4hPsFNuFXcjFScsh3Sqk1EFsSNFgrrhfQz5
w6yqTAT/MsoQoFqPfFK+JDO8KU9bLnEOao/RVaq2wyUsa0OCh5g85RNzTm+YIfYFWU52hQxCh6IN
EUeWOReKvp0TKO0wxvgAcnZzZ3dDhjK4ooPt090wQbcQzATMht90UUWIg6jro9RuuRPIf5oXqwNM
TdAVdT7LiRei19SkeQ5J54HcZLNNy2agv28hpvH63iPe439GQhqAelZS69w4XAf7laufLeOkclRx
a3OVbNYJ0MZZNV5TWltNb9BIrjVhIoDtShHb6ONjouOE9ToWkVBQLb/7qYJfXekzPcTAOHBQfpjy
ph8jtWDPm1WwBlYUg+SIWo0rIKj0yEKsDri0JiDNo4dL9asgMOpBejeu6MRMLIy9gLpOPhmVfOHR
VK9LN1JE7aZaDskLzcYmqFpnydjkUe7Kgon/HXdJYiUO98Qt551CQHia2JHUH7s/A7qkQDXQje7B
T2UTxMxYHW0zqXRIaNDDiNvs8pPP8hjHHjJ1WTh4pTrKehKayMscZtUt/sj2ikd6ogooMlj3jfTJ
n07+PSECjmcsCfn7LuTQlO1WndMypz4uJ25h+S/lFQRcM1uQxB9vW2faPMiX9RQF9nKKpj10B6yh
ES+3nEfg2jas4iN/yqEXR+KkS8dCkxtXtccfuIlFx4WE5vJHqCwbICv5VyAqu2Xu8yOP8leZL31N
vBfjlUmaDb+tk4j+na+X97L3GM+cCAtrApUWYX8h1XzwTzUpln2d6zhpCcXlNlY9/jgtlAC+ZgaA
98cW3zMDG96dxW0olVgqf54cpgKkiRGZZ7wFe9FlxHShxiuKYuroObx4ArwQKc5k1JiwF2b1+ZbB
qHtNnRxhfoP9rVi4gM8j6ZTDUwQsrmSV6CMw4yBeUul8a6BmK2bzkuXI5VkWLX5JxIDrJ8eClNYL
FGWazT4dIdvDbNVYEQ/Csj/HldvAYYdlU8IisPNYgnEsgjdYGUvghLBzkRXMmgwDPd4ncFkG0gdA
HBpFo4KvSXFXki45/Cp7mx89/0U/Tje/ze0VixPxwozoCI7VNFnqHjW2h8Bue+jEoAYHINtk4ogC
KveKWfcBbg68oegILBKDbKNo2XdlY7j8YzmbJmUJCVt2CJIRk+QwaiyvMC/PmN29bqD89G12CZzu
dL4lPG6MvDN+8DxqjQAJewQ8elXOO5+b3h1jK3zY6ow/5lzJtnMyr44m1nOIMjpWP2SL5cyMIDjM
pnOF+7KOPGmFI0S57SZ2Da1Zd/BgIxhQ8LH3TZ8klByeMOlJV1geOvSFqS5M4tf9QGdcVzy9lGQ8
m5eC4XNRmwEkciUGkBaGZ9YVYgqUxvE81PGYkb89eKUJvqlP7LfuTQHswggB9kLqlgl1lP1+6pyq
ow6Lpe76rnh6L86fBnyWgtalxq/5fWHdnILBjef+Ef6iZ40s7IKUwBz2YhEUs19oSzWYjWrN27tm
oMBlxOg2530ZJHzl84f80mycHSU21hyruWMbZ+/fx2sjuFpgnAQ4fHdgsbx7EZLTMQA512uj2vOQ
dYrYqf1pcUOrq25gz3Z0kFeaUc0Bgo8lgBjumybjS7mOc2beGrMyHlmZgi3fHR9ignExQ6SS8flk
ITAJmbercQ0rTFil6iUWxNWyaIFifEXkBefu/4GObz0KnNPMt6ANUrHn5Mp/RMkrhdR3iBJdjdui
jFBsmJyrTSoJg+ari6Jc/7QKypErZ6IWKkKfWJV37vFZI644h83N/qIMrhSZkRyRwvR6OJ35PUGZ
+GsLaNAwP6f3R/hALnpHlENEKx88w0G5JC5Dai7fbwnKZS4DgESOrkiHWur4MEcCoEJDmtaVCf6T
Jv6rQRpyORW8NhFkppjs4A1jczAkqM0BGSGcdVOC1vXs/48PcM199rO1Vxjtk/nC9qw0RcwcjSX6
4Ir12wlub991rXHZtIcLLlGVhrzVwp3+3VTtXf++kwPrBEee7yaBBkkRq/mcms3jbMd6ws1CS5X9
nznnsmXWukOxdvZ5Ljhc0ZNzc8I8LAhtjxkNkcVWqs6jfNbkJ+/Th4itzimEYqsgPT/rGGblXOLD
RtDND5lS9YaT5g7P6KACv0aoux0+rfISTms9w60Sqx1+91/Tk663p4WPg8TUQjNzD7zYRDLUs1zB
w0zKsC/2lPrHX4JycvRiuw1tszcrnNc8kIGuGiC1B58meBGqz3aL5DGVts6S3jxylQTd3qBdd5kn
8gKUm89xTNetCVljZvRVgt2kK+zps0YaBqrB0B5fUdrJcBgR/CyMA0XUMi+J58PNjow2mEy+fbnH
v+NsQXh/pp0OApSpURluQhFfRX5iJ/nrrZgUGrXPeVi3jaw8Ya8MUimhK4Wl19h2KFQ0k/vd2jEp
O9wAf5l/4VkrBrqbFR199nHGN5apLDFrIxhunNeJQR1h3nkYy9EZ2RaJ9zBOY/NFpD+G923AcNXV
7S/tpoOcd+X694s1RtzFhdMHdDAY4XmcHuL1CJZZAqTeQ0cwDlOfBYKz/zVNYlw6i526wIB7UHN+
ayuTy/gSHXmVH6ZNOJwxUkXyYeT10r7Tx3THg+cXr7mI6ByN4r64wOa9OwcuZuug6+NH6kRSHbK0
010XkCYy2j86zkiXLr5ZWTnDGMR70FroBgaBhqHdQKqW3trwc+GT+8A7sXuZaFVWarbe05sHkntl
Vqm4C/MCfs47vHqe7zjoM1xE8jhH5jmotPhhNCGm9+DWoNVIOOza2qnt19YmwW4iSm0Vqk8hwGVq
zGza2o7+gYTjEcfgKJ1Na2CH0SsyQtE6ZEroGMfjCh5oXk4lp1FHlUz4viowNAB1J8a88IZccnFl
u+FyrxP9ueJLZYxfj57RNYjS6qeaCumgk+8PemwJo/gZ/r1GyCTGme3RwnIx3k21+1ckvCSdZ47r
x06VfCJhVdrO+eLZ4rXCifaxyIhu1tYoGQ3/D4enKpwN9yKomjJYfbL7KN2o3j+HgVLgSnok3Unz
W6cdiRiGyn+rKzpgnBFsAwM+wEYPDsTAkHwHLbIOGPEd//Furf6eAJBGssjJgRtK2QiCDn38zhPc
vvnRLUwHGWeBWALN/OQJiHepUp6hIANd+J2LBG8Q+3B5xtuyDCaeJagM57HvbC/mAxS5grDr89Od
unzyrw40PMg0BCbpKlOwkgUbwzcmuVZvbUIPUcf5N7Vy2BpNeYWC02vQ+rEtPa1+rTG+k6Qb1R2G
MJjRXrVqUhR6GtVkUVLpm0gXmi3fn8x93btJzbzmREtKgCXKcYhKHB7/vBXC30j6o0eEnu0K4KT3
gcdW+ec0wNTKRGaAOrOrP3/qTYBsBbiDsyZSrRmZ78jhCyUSlsKcGvrBufUp6jJuk/KyfGpNcQJr
27KK9vDUzz3OjiyJI0l79N6UJ6tfVzRu7s/by4+7y4U12h6idfRA5LWvHA9Bffn91M7wH94zXL51
ZwB+QO6cpUWP5T4vZ1OCoQmBptZa8wHCWYWDc5h+BWihNTSSDJNpI4BjKcKbqr3PNjVs1CEH6ubr
v3hzliYWtRodLc8TVTMGicLPTPYdn9h05dlIuMQTsajUXx1APX74e7WUqn6TPKBBBE2OjeejZhKK
hfoX4LLnqGIVKNLbmPm96CCRAytofBZUPm+dYJ4C54fUG8SQrgF+yxn5/+xJUC8V3OHyo0RwyaPj
7niB3Sjva4QEOiR6YgPxdvYiNl6NkVTEgSOzTSTRZ9/ebEOIXCQHpoRP17BhJzxlGXkfHlPMmwVN
1123E+aFUWAm7AhUO6lAgRV6irHq4V/L8WLKObA5DVuwZCH66I7EnGPhjfW2dLjpjrEp2mISkdQb
dyZ1nas7n6sl1f+H/58jGWNaMooWnAnsLqsTGVPzkeKp7g8Rn1oryoYlzfZ0fOx0l7dIcPoiWOgh
9Rdd+5oWAA2wd7Wqhm+ALUDbX3LeWYTQ2DmratQYs/7S31joLmedON8JwoCEKFRDd6K/SmBDYtvG
GOFLX9TEswB7AArfiARbKkBPu9dfSBD8vW7bSl1SWkKYZ0+8L74fL8IcKpFk714rRhnFoq5MtMVL
mpsskg+pPYiUNA4PT72yEfZrQEPBkmYc3jbtJjbia8Kz5xCMRHtgQrgwfzfR6p0q3Soz1ZXG5135
wvlWZiHvbE5vpomSBFKY1oJPxF4Q2KW3b+ngrJ43QlYdRgjmL/NT7wlfrTZzk3OG08H8KhzHIzJs
TvyeGVcbnNmGGiuUwOnw6Sz/TrUmN+IJ6YgofU5vVjmlDwVNoSu7rVaDj3nUGao7CTYTQkv3qKz1
nZ9Eqpjk9b1Y+16ajOKYSdPKDWlF1IzdjKc0rsgjDt3xTzrH9CiPgb9evBYPl0QllGSNpTC6Mcnm
PJ5Zta5Nnip0O4nHiRIo3k7O1oSMSzZW2wour0+aSIiK5pC4c5qLWAA1dzBPgAGDsbBE5eYPrSzc
Au96dfQ14IdQy10KjoKCd0ThGF/m2A9vaDeMXxI6o+2YMGGRJZcaHZpWr1XD7JLn5VaRuM7UdJ+Y
QI9hkXoY+ZSQIRfEdR/eBiVeN6B+hgpkCYxN1SBL2PxB4Bmz/OcNcPIjF1RKZVV8gEgMU5ScbbX9
ONQD6f2S57Ob25Fadbm/Qpxwd41iGe61SInC8p3qfmonjgc+AzAdL34ohiaQUMc3jDO9tr1DCW3u
7fLEL80uR2AnH+cyCSFgLIKH8N+7pvhMc37GYYMqC2xgXKrWatA7lUlFrBiFr4jEGzdvybJJMnSV
G0YYav++kWshVsuVTcPRVthQwDMWHt9g2XukFKCve2cjBulg5DctubuhTPwhH2sAlb00SAdtsv7n
C3v96bZh0KRJ83yRkTiRplvQdREuaArmFOVXfl8K/JQknxApgyFmexH3zgOzZvQOvgicOhMPK3bF
A97hBfEH2Tz9ITr9r+AYXYnM2pNGWLAnwxVxRzdPdVPlaNFkbUK2hCbdnV3JZmLP0ykbQsCQofFH
f8Dke2pqsLphVAf7uCHlpsWAH3mRVxcJ9QHEBZ+yWVcmuVKdOzazs4OwxZ3pXCou9tI3jcr4BvZ1
vhIQT++4LWjsp6L56Q2V51TxyrLaXCMfXF0KqrFR2RgUvHUuzJWxdT5dDDx+QjiWyfmLKK//eW4r
h9H7vpij9v3XIfgf3shq82ezJcWZwfOi7JFcJk2ubTjx5bj9laCaRw96TRPuEKXtDIuK52YJx6Pi
RL6//l861Slan42G6EGNj+/WnJxZR7obTUsAOhtdaHSuKuvoFL/bBLV0u3gou7VDYDqycQydx3YL
OPpxvxk/dcXTeq2/0l5TfdIapw57jPVKULw/2dSGJhxv/pszQ5L1ZsI65YWgNq2mhvbg38/8ipP0
dBdCFo/mV4jJYwN/x+52X/WV+IEZDB7NQnu+XOmQrZb03rbxC5j4oMs9gFbb9ygQ4MlnnZO3wBIi
QksWSMaxieesuq/Dvs874HNrMwUpwdyFidaCOYr5OTQq33dsRmcANFwO8wU68p+4q1K6W+uTklzN
zsp5hmyX3MRuH9cf3P6Ua3P7l9Iwaq3KR5T+t9B59T5VjNUX9nb5bbHe1G4x8iMNY3EaQHYwcuRp
w52K2qNzcpgP+IWzr/A4hjs3flmdkJR/RN7DPutztCQM7NyAFHeWGa4+4QWKY8frrXRhxGg9Maw5
HjQDclrf4u6Hq8MMnVXAzrJ6/aaOMMB8vBdbKdCbjEThHMIHm2a5eh4QLVREgbPbNS7mxP5XlQ4V
j61T5lVXViiA4rKjnRWLNGJx4pkgIVoraUUZJhLQiYgU9k074jlWfI2ZnnxonSrNZVD3tkProBsy
4vi1MoWKMQdvK1KtO9oOdkcEweSujAuWZQVIqFjD9a6v7LZ7ccVCv64qNJI/pOSe9iWgudWddxgO
kuf998LbYHBbGlLCFAjUTI9dJxemi1mQMvEetEWsMJZMcyEwgtGnkcsQrT2OapmpvCq7JOQo0UG/
G8bOjpSYU8aRlcbI7N27f/v3HxAAwnlYENHQp9kjEj9chSi6bxnexaEHdR1sO3Y8xhgBBVOfDKNo
QQZcR0ipWTL0NZfKCLVbQXqHGalQgd2EvFHm7r1h8IwvLBUB9JFTO4VRHRoPSPwDtOXsOEOYPzap
KYPcQVPqx2adn+0X0HFHehwJpy3NjcmQDe5HyGc2HjBpa8H4hejw2A88Y3N86ULOBOEiDEPPJaUz
U8+nsMtNVxdk9v/esELoN29/+X7ARyDLH+UgaRVzLS3evtLTMe6qCjmsi358sXYjYARnfF6+3Hdv
AHkb/6u4pSdCYmyt2UkJ92eo415QRvwun1wJ8rOuVAEJSe9aG239pj7GYhtxpQGi3OS9c7P62y//
eJc7RDYnucbS69Dz2qUs8xgvF0ZaRVjIOklAwHWXumCldV9gY9kmWhjKRgj7uEXGF09Py8e5cfTo
sEyxG73RM+DdIMshtklRT2Y0POiQf7OaK0Fh+WPB/jf1/IRotHb2sWBBkcP5iv0DVXqNuCz3/ydU
Q+vUM2RiuJdXqite8ImTsKcxrvl/NyZAwdnOQfxgQhOlZ/k9j12wcplp9zs+Ghvt1zN7R7oUoksT
uL2eEMYjZZ7dcUJNr3CS7sf1NzCHDIxFS55YbZBGNAPGg1s8jDJXBcZIz2kgQHHHUgxFJkLjlR1C
rVBYrdvHoRka3LcH/mbvrFwNobNt/0T+BlVRVUy8T+YlEmegLBhYI2E/8GiURC+jhRq5MiWkTYEZ
3pN9u61+40ULJGQgH3uZW/06ed3Tl9sfbzz5oJQ/j2mpoH36g8JSN1vhYkVZOxOjWxbosl34Acur
NIhCgC9jEcSWKXvObTfjVwFhPTTE/Z8bhrXkZ9qJ0hHifcMii+79SCDSVG9dUskcdXXMsX5VU2/V
CUSEYOxBZTcqSI4wBTJ8TY8fVmrCWQsebWhYR+dsDXg67ZFVH4ETknCGmtO9vlVf7hpw+d9v+M8p
wd36Jm40bbA4RCtl0CSbs3w5Ws/YUH//QHJYhRZoDprcQ5H18sQtjEnJP+IiJQoEmJlS4k4qWEz6
aQyV5N39/NaC0sGNcUjoS9kVYcIgyfDBUNp/haPMzfrSKlpuI/i80i9cAQFpf9c8FljLygzxuJHg
UUj/t6c7n3pXiYUzTGg7gaOi9b0C4HhAvyTAXX4BJqHvBwSrJKH46h1d04Fc3MSL9Mbas3I6hGc9
4K8perVEjqFty7eeOInZkRNKIfbxAGL6XZa2nrcLKYyDwygZRCXCmLj81E7MyWAYJ6dgGbXt/XKQ
7w1nLAkqHD6WDiI5M7JlmH6FXEnvXm9sORB8BQtyNEZ7v1b/xafYv5UaiGl8HBtrgGM0U/fHpcRs
rTwWE3i8pSZxAfiwsHhzMLV9vueuhmbvYXRkKy2kPeCcEWNVP/HDRDcpRHNEu4CVNzVaQlhufIni
JZzIeLADGO3pdDCHXNlNX76i+/tBSn6fR+LDgiSIGqLTmvkvfpIKTqVneeDUDx5JWFK+Ynl3NZdp
yKoK9NBJkChNi96WJyyqcsO8Y/RDQsSaXOxEEhZOr4LjeP8tI66D0eOoPSKEfKuR0vz+HmGZxr1h
kGtLKy9gDDzRnNyjtqSQblkWzP12f5shEl+KQcbVjZ9mO8QZzN7djh/KUCfLg/gvHLCR8Hobye74
BlHElODN7dPWlBsEUnMKJZwf0/X1ZJN5gx7igGpgn44DOlQjVEgJNkWBznjAXiAd9chY8Hyi9sTA
BOfjv+V+EggT1oagDUsW1r+RDsHpmfuQps5/AdlgHp/9hxL9X4gBjPuVYgAe32tPtSHcl37hKbZ0
2E7Ogs9OSSJej5Bk3MOc5Bj7u5pqT2D4YE5QeHBhtdY3do0sTIcJHYIf+N++6oOpMU4z2P3NpdAO
9c/BtkQLFbLZtjoQrkiKy1CLOGTY2nV+jTG9A0lA+Ca7TDMTo49jMlmazeCNPpqRctjwdfAva7JH
ZYG6lq8YRyKE8maJWVWixoZNIcMY8I0PJOtQ4Nhie5m4Tk7CslizdqwhHC/7Xy0VYhUj96a61xtF
e7IDwf9m+yp2pvL2HPJ3sJExqjh7bN5HQYyZKGLxMHaJAer41ZMbbQ14sl6S+7l2MR4oxaLvxVHC
cemUeyKs2XiCpDv6Z+YxH8VoYA1eMgEQlyEeYbVodMT81Mbil3gS99v4JjJVBPJeJBy8x/IDkjy0
J8TY/zjGyD3TTHFSnUva5kl5j8POlTu1gz9b70L3ZU8ozrVhjHUTG7JEpmJyQKZ6JKXaM27Yrlqq
bDrqUrh9zQJa66NmQ0NaH7V54PREKod8fzSttyvaugLbFWWR/Svr3E9DbUhEqXdWzf7r/XCeipAL
JREROLC0PYdcq3CXYV/Rt8VCLtm3bhJP+WuJQqxUSLOoRvj1g2RuSGAHjH3SCUhZwQLCrFBgSITz
CHWIECsxkAMmsW6n1PikSnVzQlWzlByvwJfkx2s61/cOU7TRzKvs+L9P1hyqNzRiUN0PKEi7DQWp
BoT3s5V4GPmk2jiroyHKZNEizEPtoKNhtK020UH/+xM03DUkCCv7CMhN2kb9Krs870EHickMlvb2
sB8MMj6MHHBpJENn6CKMFUJCkLWuxXr4BJvC7aHv5E5YEzTUEsA1r7vwx195b3TI+dW2gxJQvCFI
UgfsNmL7LBnEyBQrslAzxmo+H2k1E3gbcOnpK1kbuFw5wcmpMrB1fJ52kf+YpwqZpnNbc1QINngj
JEnBmhpSHdVqE0pO0DrDaO8pV11mRQoUb1KbxnkNjD4s9zSI0Nwlnmk5LhRx2Zpo4Z9lvvf5YqLk
IjA8CGw6FPI6KgZ6E6iPAyzi4U88vLRte1xwphAK2FZjYN1if69PhEjvhln43Wmcthmtdq0c0JFX
Jp4F0dSnfbhM0xDZ20dOajlJPm8f0junfVg1qTdCuvkkc5krFpll4QbNvd12pqpaf6h3SHiqb6Bg
RNJeewduHlx3I7lWD4cVI5B/Ds+7oc46wkT1CqhIlI6wF487O0J8Joth5YP5o/RbDSXqtXFK3SZw
mGw7e2tWvv/oeBdj3XJDij/9h/SQb5BmCxKDRPH87joHQG013wexVGBqxJF2c9X4CGS98a0tDari
VDX6ny7lgyLe/zOiK4rRw2MkXxy1/XRQpPZxmpogFZ7c2Z1UfxEVYLlznuN2UMfzOTAXYjXb4Q1d
bI/G1xXxxPpWMvzLdTIbJs/umaG6yY0lqWDB3AMDN1XnGx3ISzMRXunfv5b9jY9gKyYNUkfk1p6s
OXlKuMzVtRcDFL+mGCNC4ojiTUIn6LXLhGlKBlpx7h4IckLpjxp4wqZRT5bp52zmhKwFVAueGMKQ
lKBVeHmWtfv2AK6oRjXakxRnRyAVBa7w65N5acsHNj0GEFjSAJoijoIGSlTo17P7C5BOwpPzx8h2
hylZFKri7iQN7Ijt1nbahvDWdf2KyttVS/uB+6kyIep5+/2QR8BmsmaX9tpAFVDc3VPfWp9oZfeP
NnA0gO7Y7+Z/akj0kzTEym6tvruSnx93i8DvZy1i7Kuunq8lep1S/Rr0Ow1YijBdIE+W2S5XgWLa
AQ7MqZGS6G3RdPD63IGUTVbDUVswedgGG+BO/w18q+Vxcj7zvVVRqyeW0wYsE05YWkJ4js6QH+oh
3OM7ZwgT7iFs03I3Fru59BhHkXwfeUkfH+nJg4rZOhjC9dTJXdmgLmfGtCbYInN3qdA0G6Nh+b9J
ajcPtA/cn9MN7nBDNeS8OijOjASMBg5oq6BMm26U9UumWUHp2w0t6B/nFB4HpDF3IWZmc1XEbAY3
L8DPv87VSN1Hwbo3A0Ja6aynKEVdIIM9M4EX7NeZuRZq3KDQIo4XZf1izLnGMecuodwy/KPPFUxi
k5D6PZWO2Ln/RE4QFIsJH3Mt9eUGppzVi7jZhlq7oAgcFUBi0VwYC7Nrp1PQxXAEvdVbY0LfnXav
hRVrFsHqE2MA645jK4eYTERpU8wMepYLafY4ipadB5Fpki92ERN401ODpS5OQ9HVUCqexU4QxtWW
jUik1AyV7XKcr4S+nwXk5RcBC4NO0KlmC35npt0Z6XWeCmUfY038IBtma67fdiuKUfb6BbC8iSCc
RLwcYh3AsN8VrhhuIvbjL6laNUEgIl/Ro1AnmtCJA61aNNTCCv10LkV1XxYfcYOgYH3MlkPzIAXg
rJQz+hJQt9T1Coy6zxIJGfAs515hvydhKYkZSAYwZkENae/kH53H0hjJ89xJyrFv2gfvgIF99JPD
PrQ1SCJRrQNwSVosqPI5Xw5BZwxd16FkXZAUwmuNTQTbQXRTf7SDHzzpu2+bycZHoaA/iC55nBRj
QDKmyzCW+EIqEQ7YyVyXUi2hEHF3nIsYZZp0VeDmixKgURPsFvnnYavFqrD0BdNLp55nyEKtb4p6
gGXep4kpTsStMt8y0uSPKNY2++Ao0Lv0OwFaC1Qy5SGbMLl69toCZ0mdyNF+qbC3TRohQU6bDnAu
Jw9vwkIbsQxwSkFICxUqEwU2GqJTCJfiWJOnnOaJeeoj+BKRfNTnWuulWnMLM4IwSOkkkircLJQz
b/Ugqqs3Lr80SaQz1Omh+OPDyM0gR3D3nxPHixiF4G75wz6mLVDXT6dh0ob4qwPnLN0Ig9IC8bnI
SQlxh0qSwEotelZo+JXwKmtG/81VMjzYVux1OIMyeBTBUZYBphVCJiPbl3/UipeLPwu1hJB69fKa
YO3E08AvVSEcpYevDAZk/HYduojYUS/qcu8xz0wMdr+lsapqmYjO03ZM7BGflltIk7OyBhlFRefC
jm1OoBy0xMd9FRUq9ai/HH6qzIlK64SvyW7kHWOnMuAjo2217y6rx0AOMc8tWCz0AemHP2tzDbj1
SkQ1TN/Ye7WAP1xsnWKfEixCgBtG4wbzlogWrKzqGb/ad8chMZsFY6mctj4LWPF4TJCIa7gfgc1D
3oGF3ZAjZcurEICckvLnZ9IQOnZtqqgclmIUyGGbiN7O6N3YkdYKbFf3PKje49WZixyooEWioLtP
V0ucWBy72J0k9SM3Fi3ragLsMqefT49OUrMrUI+tc7RpZrXHrRi9YN2aPS50BPeq5O4Rj3DrPCYn
/UaRmCSY2giiOfNJv+Z/2JgUD7VfOLqx+s9wdQlxKRUoFFc36TEkh2NG3z0SSMxKopajTt7cV+gj
H3Vwwx/st2IQYyzbPmgiymwKq+KeB1/FHAqD26IhxQN6XlVWG1Qb0heW5sWU4rA7mQekqqfArhmi
JbIOdV+wzee/M4h3WHRMxyLCXAgv0ufrvDejDVWIqtYHk8Um+O7Jjhz5fNmhBR2giFDt82RMgBiU
1TmEIrEVNgLN9PPB7oncxm14439CC5Dwd4C9juVOENutk4jXigqhMkkIVBC2edbRP2K2JEXKmnyw
2Uhn5t4rGamAIkyXyrA28lVfZUT0RK4TSau7RmIhIkD6lLoc1zHShHy6/IHO3ObgBKF/IXvjQImZ
4Sz8eYdMPDREOLtas3LAHeHha0Ve9Czs3tZ9wDUO2JgGXi+awL/Dh2cb0jmXQuYo1lAKHX0C4Guk
98FAa2FP6j6B95XRWJR5KL1fzWWb1Qcjr6F0trMtS6BdPJiBX5AVUxxbPFSxOzwr2SpUwuAhKL7w
S+Ji0Vf0mK/cmHVJ/eqh6Meg+7KOCGenUALWZrzNat7jhiwgt+MqZRt4KIfGqS00g+0t5pH9AKPO
BSePzqq7g7Me+bWPqmpjr7+BNOYPZEj3GVkIX/EzuNilMJegqT5QQFkfRTgf52kqEjqXq+4BPt1V
2Ngnkr+oiqGetnFuEuWz/y/W79YV+bgoOJKA8UC5tS5wYSHK8fpx8Jdl94kJqehKJeLoaOumLwxl
OP5uFQxkkuEHwoOmWQCI58RV5oQjkUGhj+t2LA531u984Ld6X0maVOefuPC4D9C1KrM6w+dnT8yz
LyF28sDgeIzAsE7HY+iib//1J9rj6hse7791DkQIJew5ZpgKahl2Af2uNA92EC4+bw9ZPaMzYNMQ
qf7vj4QHyDHovmp9BMgFOoTjPxXJzezw4nAK9BFAAuoZGTaGAwzcxgZPyhrbQkp1vGSI6DZKXaAw
oy+w3PK1u7iZZXGJ3djEetVTKZzoto4U2XRwl1mNbWZIsmlbZLvAlIzHtBtQtumqBwebbdALSnwY
Ow32VLtg3ZXgoR5YKhy3nqEz+CS7556ts4cH2FjrnP/EiTT4EanUaM4HrHkdrJ8w5d8+BFlN0Zse
9oesCbg5e+rlplS2R0XuS8gqzomQwRa1xH1tFqKQlfwQ64AAod78O2UzerqL6PA5cI+utNYN+Yzk
8ko5j1BVDZZ/+4ZkOXLxQUEPfl1tL39iJdlfbynZWWP8exQVHI3d+n0uzWNQjJ3cbAf7MQcaUZ0V
lZozVEPvF9pU7QVxsB/TNAVrGqVj2NxFsONVWtLYfaEf+3Obsc+6z6XzMaUwtZ0x7OjhqLBsXXXr
UB2PS2qOE6tpV1jZT5LXcZ+wy5b8EciSS1H+r/+xSobuE5yBOfNP8xkMbGWzWinJWLAwVVxfk6bi
iPIXFp09n8pL0KSYf7pswiw6IjxhaV1gyKhwWOH23k3AEYmRxOZXm/loc1sa/LvkCkK1nKQx9WkP
Qncfy3DYIUi4B+jhtBe0xkoPRnr4/dYRlygDbql8LPAZZYufIvLIZG3XbRIi8jRmIGPLqgpdoiHM
w5IwlHie2R4xdR0yfAPOSpeKbOyovZKNiMJ5nK5ZkQDVKRRhauW6oT9lHwCx9ksvA5HMeHGcsR7b
0m/JSWCbJKea1VsOcfT8a99dlkY8hNME2c4etH1+C6G+mhyuRZVMdpjf5W6R/uNUNzPW8g2mArUF
euj33UqSheILJvKWvlAduG07yeNnwbiAjp8Cz80PvoR1L73Ad4AJElagWZkYR01fqEOzeYHQAzu8
6Ui0zLyUJ6KL+V/uqfwL4c6H+Mws35HGCgwhEMVN0/vK1miqOmOZA6SBVUfPPYSFKkT3btlPHzML
J99Vynkv1xDgceVg7W+ovm48QkbHqlZXXx+qPJvNWg9JzqbXrw10kDnS3WWuQ/7ngilAEHBMu442
d/fAnlcPqijnybubnzjsRgjw2O7Var94Z8IOev5Q6tHSPNcRVCJ91zf4h0jHm/Z2wlRVz65E9oKu
TvrQ8PDGicMU3SDlgtBW6LJVGF43U7EuZ+lP3If9EzAh+qT26wPcOZ2xQJc7qZ9Fsfj7fyx7Ka3c
DuCyAPurwdkOGPzH8RlBmAfpsuZx3QMLj3hQsz3IugPKSu3+leZnjpA6fjkiVEzeLckAZfGXlrzL
FL3gPW85eBiNlyIECliFKF6mrI7FVVvAC/ZbblXwwA3VBhGEa85QMCF507Jw5fgmgt+29igDQHXm
ypstJV7Sq0JGI7xqixhsQZ5gnW+K9xPJmTbgS8cqBKJryhnIO3BxCNYdXhSZXvBo2XSgLf+kIcha
Z8f+mdui+ul5MlDAPnaWxW5goMR4hXpT3p4T0AojVleRZjSuTKbZ9EqBnSE6xbFCJ8bPqsBjhTin
v8oWk1tBFHl+GlSQ9imiE7jfKzA8XGUgnYCgRdRqYodecbfeo8nSGIX80VnbBCgFNJs//wma9M4I
4ThanzBNnXD/PRUqO7LxUzEmbukAQsAgkq6UZ2ctbCGIBE07+5LGe/Og5Vwv6yrRvsiNHf07MQPq
maKCc6m4qHyhWmMesyBsNYxJ9t0rKfaopL1dh94uORjAN7lGLU9BMyP2BnvJVFgunjC1FRA/cSbr
umBAzPzKIwKtV3OHgJz+NMPEd4RKFctXRbmYv0QnQ8LvyKRETLZA28sJ/1Tfg41/TsAkMYEJXwrv
82k9tAzCeP8Jdcv8nldj3JKwXXt3IAYWUk31J3jrPIaMACJ4aFHcLLt0y+vN01knBd0TIkCQ2j5t
l+DN+UbCQA5puQPT1xzIKxFUF9jYlWQcr1Xqu40feNESxAfoveaj7/raqzJfc+4voI4cLSq6smKW
HLimLH0uMai9xmJvOfHIsmIBt1QdmKq71TfMXphOR+ZMBMuSGY2tphUcj1APqa9jApFQSZMmpf4f
sWHvk8su4Lev/byN4XxCXZj9SiVPHWKIli/xkdzzPRhYQOhJkhq3nDR+ka7U51W8rvWkObODNhe6
/m3uQRCQNXnTtMKHhDe7uDf5a2vhaIlGrAgew9v4faVs3WjJPNg+NKeew7cQKz6jLxx0+iKrGdd2
W1rnQqXj9hUzdplFH9cho6F0ULxJQcaHCYjqLAQpU7yn/3VaNqGRs8OJn4w9dc6hk/doynvzi4Xu
fZndu8RL7ZT2epYD6GFYhIFnbgLil2G3+UrUpAwArUWUbm9NkBlzil2ACjGEWcqA4ZerzKgRZMO5
sZKJgEBKwI5ENGMBiTvw9Y//EsGFqweCmpXd9JrGPdoHvzPXZ/sd1I8zT4APgM80pUMcx5TXhsMY
kx1JgoeX3KCxIXKd2/4Qh6jlVtSmYq7v+iW5C9aa6uzBbBfFrC1ZGl5gBgMZeVkpxa07Yn4JUEWx
BEW1S0xcsuTVJZXSQHfQ7GB81iufS6I5V/2PgmvwIDNygozMoz1MXa339hKb0b1WY5NPOrCIt6FY
sG4Sgb/2qi6ftRpqpompGe6X8ncJoYq1M5r+Wsi60ikLVs4U52jfQt2uK5tfIxcUZARn5p2N82Un
b/AVFWWtzivtkJ35P+7FCWjSPxQCACLt34HksJFPpIYndnhHOCFI0Uq0lkd/rbfDX4tHaJY+/eJQ
WKRxhLd/rp80xOaHTPAlpePvLU8jZvEdOf1daFwz5wcHLKIpblNkBDBRZ40W98Q7UZZocyqfQdgX
/rykj7xGnq5xv4dHxTGI8lSsQQlhujruLSudBDLiRpLj+yobN1DxZvrdjgmkgeA0r/suDMEdNN23
CXiR2RCmUJcd01wRZGRiz1Ytq3Ir73uWZYhMikmX7poD12+vm0xciUWgA9hQaPIFsrGyp6u2g2GA
+Jkz3fT93FCpTaj97oNr8ghF4u4ZH91f3MiEdQxMSQXJ1Ffvte7RkBm3LBDEg5BTGfKFz4dURIWf
2gDvDKgeyodSXu8TsojwDya9/7euqv/p9vtU/+jB4HZfEYKd0yBuoH10zFgTg4p8TE+iQHhvGYSK
9RDovOoorXl2B3eOCifR0IctFV7r2QFmyCbjR+VpmBT9WuD6xJtDVULNcPzI6NGXYpj4o1CxdDaW
bvrQIzCmY35ALBX7o2b0AekLjQCZbx+FV2FmCYf196CsGro517e6Iq/cVNPi+VuWwr8K0GqdXe1b
yp68LCGj9PksgV/wQX8npdatnunb061CW6JFUzXmjI6AkhCC3xz2yoi1EHHVE0w158skMvGnFkPB
23fwoyws37E/V1P5+TZHiBvRaVAYFTc4hLtAFQL0xNqwgYksz5FJHqxRZesPYeNV+8lX5eqGDk/k
6GkvEAyhV8GkSoRksMSog4C8FlObHMHmGtF2olgEWio3lvUZHQGSFcssrTBK3MFFcd9zfdJQaGJe
GVifxYlWYX3iGvXcXSJC+CI1hNgRvKgRw2+gME8J+H66MDfKPhMu/nhCTaq5jz5eFTVRI+K/Asyf
W/xK15Wa0uhLy4Z+IFd8YMuTbrUpPHbGO64pntA+derxDkBjbJnRCJ2y5gqDME3+iJ/b5VtAN5JO
svGySC1OqKd7tw3YGSfwoX/e8zR134UWg1K9iQQPyHfY39p9G7O2EW57oXD0he/R6+0ohtDv1Qt7
srh7nM6GZQNFP0y/daxHUPp5TAZM1WAUK8trqrVLDN1zjAlriWL8BS7v6g8hBB7PxWGaPzfA6dwu
tp3mhzzkwDpTOhDbz3tHiUdgpldI4DG9jeT68wWiO/1kiWpjku2Y/3QHuxXQ+XFHCtvaMndtx1mW
O0QbHE/eedCjcwU00AHST0n5jxZUmTPFBUdWTRUAm5QBMgXbBFDw7aKiVl8+Dp5TYHOipGKHNnXR
k+jc1g5+Q7fb7OQVoelc5MQErzRYE9Td1iAENYW4wT39ogF+TCNGwO/6mZvoNkDjcncwwBx8xN5C
ODjSSj9rbdm5j6FbInnL/QfSRskx1gBJ3B1vOyCeugKnSYl7WLoytFu4Xmj+e1D/4hYpvcqxDXiw
gJine0qJxaOaEdwFwtUPSh3WHPP0vP19QXuQnNmGRHfxtQPvsGrya1BszoPj5ruWf5vY7xVfhpUc
1yLJ9bGm28gRAkh00DxLRNs9kvc6fctvowVCv4el5tTvjDtwETARZFmgKALsaZs9U0NSNX2Lj9f7
q0WKZxi1fG47ZW0j2dm0/PQJOz7g/oRXc20FwqBBr5UlsY9xq6DL9Gm9M9NLSgVJEwK35yjeMRwB
znncmLfV0kiYiv/1P7ZYxs97eKFUWOml4QL3QkmwOW9WSe+iQppk4vPag9jvuJwENU7n8z7UMpck
6lSn3cEMkxzY3MU60o+PJAfVGuRIQLYcq6RSw1A/2vIEnf6sVZsDg7JBpCJU7GOc7H5ShJYgLFYR
HbMpRcavcWBP8pfLASBfjTV+CdezogcNYRCM3KAWVRb+SHTon3tTLWe5dJaEKK1f2hNaXj/9S6fJ
JytcenrJCcUoEHVZBP9ih+lQCsfZK1sVukxuAqm/k7g7GhaCb11fm8vG9Wclz3IVeeIsevF6YzII
LNavjrK8cbnB213gH2dxbqlJxmO5G12N1p7sAaO+huC8RIVncU4XOSHK4O1nWb3R0FCCcZJ4XCvK
+6IGeWJXecYgbDiCz9okB7e9f6fxBFd4QWkdoX1nPGaJfZxckknhPH0PUwu9rtYeeg5nruFw+35H
ibzPMNbZaiv5MCupgzFKluL2cJ9w4a64/hprVsTLOoIL9Sqnt5kNvtsx44hQARagWoKrgJas8cI9
aM/bkc8DoYBdaij+YQgiJxuwBPG2Myiv+/Qv0swJrj80evRTymlnAw2eDYNkTIBuJxye1u5JyXx8
hA/NFuqLucIF1OmygzF5j1mMSeaZR9i8bWADH9nJZwpjUg7BWCUjTvG9C6+9HgNPOHxPOt5h7SAI
2ODHcAi3tNyCmnb/ih49K2a1L9QZ19ttCkEgE6tJCS09qoiJ+e74SMLiluVm1e/aKaPNQc9xTSkM
cDFZNz4wW5EpHCeFOlkRMFebJlouGfOncYxuFdAMzJchoPBziG/JVazkdFCN1BsiPkmoDJ+mbpV9
1M9Xo5mqN0jhunrabXhSKrB100LRzdF/erdZ/gH/8avqp25CZyuxccrpwK6wW5+NQ6JmhGrfT7DT
8OD7v2TFx/8tOBnw1QIxzkv3oGrkp1RU/KOdsgal2tqE47x3IWzAdSAsdfPA638Uoa97xAVtQ5FB
qUpS4YJG0ldsYI7uZUAeau90CQAtG3ID0i42JnnekhwS8ZlJmvqUEWeakgR6R0HmKSslxq3UM96V
a9Sb7HFbMhGm5UM/PjG3BDoEcED54v1fC+QsnrSt66rZ3bRbYM7rp/bBqK3evqqMj9MtjniCBMRm
M+sJvOUnRf+rrhW7dLw6fPFGpdLJoFHs2xR/GaXGz0QGMWJxrshmp1BcaVbkiWx9q0Ee6tL0bWD7
A06Ho9JEkRjMj1xVmBrjGFwmHtsz4qS+oCT1onSRgpVahMJ2/gNC+uxot6DUvZZPNRhr7IVt21r9
zT2TLBmtLckBJGM+LrZD2ivHQcVKrgYelGWrmGLVi/drDoPuAPBF/wp7keJn+O5daoMkC9FYurPp
GvWUSGEakg/A7U+OtxsvG9MThklVbEiAMbrDrAUNqeXQ24NMysTofBb59KqJAHfkmU2bkQ79j1Uu
wRWI5C9H5D71wEVEJRC2WL2J8ZJY+sZn1TpvwyqRWpN87Sk91nKHqPi7MiPL2wzTQ4ZwZUwnriKs
NhmDvFOaf5yOQ50HYvWMc4Z7NKDXr+DkQOQ2yzvRJixUIqjulVg86YHgDumyoAoglm0XUCQn9b/d
pGmiu71gea82sidn0oK2gbRvbKIUcHDi9LawywynjLm7pI601B37el9AgLTYYnMIetOVoFl92SMl
edFPF5umUM1Ig0PdHOb/AhO1kFF2E9Yr0lhEM13nhzwgvFWyUCR7yOhV4XFZgttF6sMXl2MUmqcD
UGrg61nbX5W5EkyOi85htt18p1k+4+EJOgaCy9irRKvC7pkTrkYBzpDbBN5DuW1Yq7ebSCc+kPTZ
Lf6Y7nytRqnjeGmgvm8Pae7qYSCwX3m3em+eVH7rIfViVwD/FHDlTbwwmGsvQIyYPVNodwhIsg/3
vgfD9CwSdOWAxcbQPdUF9q3yRrGCDdhSGsk1vNt4+HkwPN3X5+7GTrOc2tHixdtJ/JEn9rpGOpK/
wuOlLhYXSbVWy1QQyVAGIug+7qtHQqPaG6sG3JhwdTRXW+uygTPxdtgvLYjTvo/mmjnyVG92xxbT
FjwyGNIK1nyg719nOwvXEZdEbkc0GTyPwHOA8NFSijfu3D31sBaplvKc1fVCs2rKKuZvW8Br9wRN
zx9WBcSUSJa/ptwZ0plIsZCQlXu63/ciKskktDRm4h+LjRpXl5fGXox7w6CfGiYvr0WSUhBOMbPe
qL6zpA9A3PJV18BkUYeykj4jhwLMeXHvcxxcRnQZ8rjUjYHD/JdFLoWl1tI5PH1r5R4uMoNIVJN8
vbHyiUI4tbCUOMAvu52tla0WxjOOG+uQ/AVKwqXcQsbaKbcAeyaB9H+aKdyTzqiEfQnYt+FRN1OL
YzQg17k3eSvjq/NfU+hUtSY5oitm1FB3ACado2bDNS1a7PlGjhO9VuzT+vEcYX851dRKLEXUXFZ8
TY8UwfcsGXxIBOsUnKfhBp8GTZkwlr0rG5cZbGTOeVKSflX+uWkdNlUeEsXvjAN0X/xhHGcAJY6H
kyRTWncAvBpR9vJvRznhcUhZdMqiV7+pNL3jTqYGsqCvKMe/fZA+plPwzkY4XJZKu+xX90xWjOum
a3oH1Oad2SfmyWsOJN2hQ0FMYRk8az41qxylZ21KRUWLpj1zul6CahVVDEhPsa18yvMF07gXdxTu
moGGLfcYJ4Jm007C4C0wXuH9ruIK21BbazT10rZBUfq8vP9uOMDMG/xxXIAFWNF1AyEQCHCVU38U
p4F88DQcwJgwEqMbPEKn7rYluqGZczNj8JUXMTg9gvEY+AlY8P30HzwaV64VuNKwD9h9f8pV9B1U
XJ2FgWIeWFP29iP4nG1W6mu8ZjaZ8czZjaiYQPvTxG37O+1netAHsHuukgF/EOAsxnr0ENPlOsFK
KICCrUFtpB/rJ8cvzHllLWJDG1wyr6G6PY7ABO5CHMPx6VD/uSeQKEIgryRvmHtrSmPk54LIN//+
+BWOf1xDuUCJcXEFkeofhNMij3gPq8Smc5gLQDR7Fkjo/tvyUCv7CT8CmDZTCyzHeW7HpRp0Rcfk
MGObD8+r6fp0bDT7t0j5tox+T22YqN8hidpWLhJqKIpYt0+hmYnNzbSyFcX6PN4UIBy0zEELjrLm
Zp9+xsRlnV3BwNoKifb7JbTYYeIGEVPgIjVfG7hdLIyxNHp7/39F9HH4Z7ppamlkpM0afdFtbVzs
a826QEcpFnAPvXV3UNlM6VhmXqJnDSaKspiDt0CiU1PfIdRRUzDyhKpqwWXoVuxOuKlodnCb6ENg
0i5/G0KjwGQhJCNMvdYCa774RDIJJCohTxPwbG8GhaNnfmtLjHV6nh3qKxwJumho6CxEqKBiO+2m
oq0biLOBL5Zp4tAv10xOqK1VNUXccZS9iKB2busn4dR/aRzoAPLltqsxeOm+AaEpsvtsxaa+9WDj
rrw7wwBVW7fFBDw1NkTsmDXzNQNc3xGRFxHpqngkwL1PujwkimMerhuNu/e9wkkiWp7d+yj3GYRd
qsYSmP8OIUrHE4exnki1XMV4RLO1/mLyx715UI2POq/CocRBFA93+ldpkAJv5AhBKdm9aAyp3bKw
1OH/zc1xWdgSQnwfbYDZXk4zYS6+4irEfswTx5w6+YW2Wut48lJ3RSnPufj3RbfjSzKiH33lC7vr
puYen/qiN0gurZRWMXNt2Kbj+nrn1y4HrvP2CW7nnob6U+xfMmepB/qmsAfvNjY2p+pNsgy2QB0S
ZC4JdTeNmxsuatc1d7lKAFrl0xTt+O2ti/QdN217njRcM5VWdasgRTAmlLbqXu/gIX8TNHkN1eQf
s5wZ2zZRp62L0+xJgtlCxMHGJXkF4zw3vwmLtxGpRMQoWBKs4mdVuv059JeKakW3PZQ7i53jwyp1
ew9Kn8uOrrWkfSpmhtW5Z+qZXKakhTqeBiz2BkUetQ7dVfD1UVMuaD+biWfGG7HJMHM8ZV/ZrHeR
4qOsJM36fELuuA/KxMDduxV3LBpj8BW3wSeeC1kVHjKRgeFaVqKHWcJhIE6s8SkI0FN33mfwLr0J
1BmVa5zoxoIo561Uou8ZjpyjAkfRXP0LEPetgsmsUXG6mRCXa+CnoD/Ehjl6B94dl6LPgUaWyeHN
l2bAcnB4Zey1XzZIkXJxnNP7DgOjQyyp6C1sa+xqD3x1jTz/GDHZV6Rm+lAz8wOeFeZoHz4k9c53
fmBxv66PMLtKK6cDajLIUsjyFvSKqzPiQa0JnZNjXmMIT5dNt2Pj8ae9Q+iNNbLjb5wE3IAVx381
DuTcyQLrSfnG2yJe1Y5GZZoBrUGOJ7mKQEznwQScCrysBc9PuMK9SSTmmYe5fdqqK1PDHhP8BxM0
eac+ImU+VuWWnjpmT/7LB6a3+RhqcbfbvxIi8yvZKXMHxbDVCethdIhhfePdqFAcGk0R3PT/DXOz
QIK8rcTDDVQRo5OpuGPF3nWqP7sGd2inxc2fDXG8KmORXIOSe7JrEQQ+vpLvtVFF3y8yaF/TGUyW
aHW3DuZLhEQKg/qGPV/P1f2MXtTV+99V6rQ4lo28+rjITjo4iNv0vFjNyMnKVR1ZZb52rwrFPxUT
9p+0OILtsBDf2WK3b5pOTfdH0Q7C77arRVvun/TBp1IQORAFd4zTU6NDxSC3dDc9DrLIQFu/CKvW
iD30Xp8x3olDtRkwNKWlNRxbpYH1jHkxvcccIDeW/TpkPsVZzGT/fqJmBUTo5PgcmOeIAWZErZO0
gQn81KiuZVKLX4jpbPlMYsb7SlCZnDeSks9/6h6We3vIDsh7XKDVLkfn5ECiiKdZ763JBzG3u19Z
OPL2dxl26/pgkJhJFDBYrN82CDDXmhNs9zB4MORJlfN2hldyWlhYyFLpkIxj9Hn3dON38KpvQ5Qo
Y2I7rdHKep05xrD+sVeMda/Go6wJWh+fvyyjbpJuHYZMwQiySVmf44y4DWX+5vZ5ktypsdopq/Ss
e76v44cApZBzJvDejCJ404ct3LOJOFMJTHlwu1Tj64A2c4EXOqr+RDg5nUvFwuRzrkaJjJS+K/Nx
8HmxjwBZ0UhXUguCJn1wf2q8Z9PfBdXAER4GSwy+vozwqo9vaPILnqcvDaVn/dTj3DjFPtmAMoly
reTU4InG6As702BIx7a2Hn6Gr55AXSaPZg++MysgSUYXN1H3NHyARqkwTnR8VCLHPrGFWwQsSlfx
7kxFU5+OZFHPHyGlAgpE0IJsJac6dREYLx//YHnNU+ER1l7kT9PAivFx0kPQYDYPMRFssPypfVAX
BYgresO5x/L4ORV1sao3TozHInuqL6/+qtoGu6JX01W2mpX3K8HJSQArovJwyAU9ZKLxRpsEqyKo
VOktnceKf7wuG1kYrPygfJqMeYS4bYQFm9Bultml+QcXUTyuD6OixI7rF6A2qh/eWZxEQbH3oyS5
k6cgsLJXixbfMT6BBZunzwI9ZhIGbZD7suKjHzscX2oCadlCLXDdaetVQwDOgLlk9Tla+AsoD1Hr
Nw3jgbo+jz+4DZkub4RMiQtTxfQS53cqYTybD+3ODZtpVL0qEGfXiaxPhRTzew17I+ubnKsqERil
rVKfnAZvzaUhLCCm/TCaedkaNQsMOg/aQ7NDgqGtvuvl4GTj7megvoMcfR3ZsTQrGkDXYcYxUjqh
EFaFy4nNLi+KoV6heGAmndvEXYFu5OUVrgvOiPgawMAYsIuuaiaesD1uwRLl7rERTczp5n0NIoay
jAwHNd1FHAC7Qn7F21S3XoIMv8AMOABB5D4jZUBmKiv2xcndEKb/X7fvS5raHTGMk8HeULeDjDW3
4XrbganTDG7by0F68n3bxm8clGrU3KT632JqJqJQYftLKqYMcVyQBAWjYqOaI2hARdpQywcA3pb3
Xq/gphRGKZrsp36/JmQn9NcyIvoCYfv9BU2x3qHbLo7cSuS6Ol+ciXJhyQGKhWz56SiynwLPSkkx
5gsMh8wbXk3OGZ1o/RelKlPUAAoO7cU2Mfp/QVQvJFtslA9Q1HprXvk2NohjWbEtvPW4C0xYbPPn
RsjatML3IHVmYqKidyhhf5KGhO8i1ByI//y+Fh6/C+3emeg+R/AVn7u+4J5q7BdmLW6mvyt8TjkI
h7Mt/CLZJDbfY89CERjGS4vh5zXrrKYEfhhb3OMNFNxNMcWvDYjH75p8CDNNYX8G9LjOYX/gJ8Q/
homs8edXz4OVfXFNt4dbglxttQ68mxuimHcdppOIYZeXhA5pPxsjpoBkVtiGBd9ptom+g9jmgDp0
2qv8qZ5Pwb82lZLAXebOHs83JO4t3IClI8a/FxWHiZEVt/B9naE6RL/kpgpVAemikRKazjyPVKkj
D28AtGR/9mzLHyik7dNCoHThoCJcns8hpOV0n3JiqEdd0KSpbdnCdxjXsVRiySNFPNOY6yMdDxX6
amXz/0vDq0oy8opnnWulHEBLMSuxsxFOmWO/7KPp7Pr7Xgf369CKIXBt8bA9eYTMPXa1FcoAGoi4
8vtXqNLEeFcI2OTjpnF1s9wi1c0wJOCpbGjslOCHSYT1gfVer1n6TWvNZBoezkrQEDQ03MisI5sD
bdf243xGyt6etBAwXKYgA2NNo9L91ODf/4mfNqtLcDTw4gjItIernALs8zG/5IQMo343Ap4DhNcV
WKR6rEAMZlJuoQaOerxoD3GSsiBUnrhF4Iy0BVrGnaiagbQdJOHuc1ENv0hh5huQyl0fJApdQHDZ
oIBlJqqgXKViRNQNcpaAZ4Lv1cX1mXoEksle1fRFF03PjLRcHN/LWtORcuPqPAAEGvjD649gzwxt
R9lbWIJONRMpGKfQ/Z2wIZGFvPdNV2jYedjOTa3R7Njoiw4hkYyKevNobUVqeoJLM9hQ+T0xJVx5
XpI4TZRId4KWwD77oQD4d5H/c/U2lcNPw/9fQxGsA69ThfuPOV+0LlshImadjoh96f/Oevj/D53Z
ZlqRscl7JW4rsksoPcel1qmQiynG3p2gvm8cL4cn83HHDXBMbitDhejMlJb58ThMvVXP4HYoZGrN
d/4FEOE1qheV9SQ594lwaWZVxfkhZHLTW3lFosmXU6Wt7gDf2XRz1GJRbKlJPlClQT0gnQmYxmG9
piBqAY5hq+svDjWvtYqS8C5w2ur4PuEx7P2ruY3isvkNoVEmb02fOwskIUawhb5V/UXqTUCmMNPr
WMcTV/YWOVPFEnGHsJUZcY5zrSC/zb/RETZ4motethUQVrmrRdOMrS1H65iYJVSc2HTw5DMO7X4P
8PwBMVQZhxZ1IM5wnWibq7AGqc+5jAvNXI2y+NNlVzLXlZ6JHyg/NnEXbkocaMB7MlOut+ditxQr
akEIpNZTxat6euAbrdchPixFAVUGS/xV8gY62iDJzfgNg/uHiwIO5ZEh6e2Hwt0yK4ca0cln4Brt
Ad+iibHPlU1B/oTlygm+DceDFic4GunhNd2HwpOfJhI+mjod5z/xE/ZcTx7Uh/VOKyfBt7k6KWFT
uZPVbaOtJGmdw7N60/BJVQ43gJQAuvz9WzaKBK14PGCPtsGZRAXII7OCZqIP2I4DKldpo6AxCgFc
91x+Wi7tor/FVW1ocUIzmXwnydlspT+17yIIuOSwCLJuLgbAJ+ixxW7zXvFhqetRjp6V3E0VNTyZ
YxhOJqGv0Kr9OST6qLaZhwFPLCttX9QP/sPCUktqOQDtVNH5w5DmfFXoNIoHaWjuvQdhIXrtmv+W
hXfNSVB2jFHRSrIF+4TVCFDLVcFAfTObWLv9TPXPg+3bHomk3mmF+MdXfOL0E7O+f5Skup+0vMch
N/XvjoTe7ud4FYzHLuP63ZebaTL6+hiLwaiNEKPtFTkrwGYWK927HFRt+KSku7TezmRjSLdApUR4
dFqmCvMLcuokGT+xItdc2jn0eaxQFlp8pceHKJhAyUE8KqPQ0djIAtEJ9ddkOydkV5ewvwOMCqK8
Ka6vh9GIePaarbUM+rV9DF6XI0hu2pYOUdxqxPt2/yowSgZb1+7grxQCBhMycem/PsNmIoHzmzpe
tDqYdan953ZnsozdS7v/xsKY8aaoeTHUvMm4x94QPOeBB59oiRJtmk/8057mnlxciU2YzqJt3zWK
l43kUODu1Dh/ICvxuHC9hD/uDIrD+7d6OvzBaOjGm7qKtOQCMzw4Y2s4D2KwpNnuwPdI8QK77Swn
O78d5iOTwM8TxKK40i6RgtZqtGzylS++AwzU/NYDeicMjGwMXmr2hwTFV+W/2Ptro6uR/I6GjQWF
L6aEqNb8z5DmdKDHlMTRy3OUdJWNZfkyNhLyMBtRlmOCACheiLjFBWY83T4dpS3FXpUJ6so4iQG/
ZakAlB4/tkySmRH46ZX4f0MODqm5Pa4Nawt+71KnShJFblTiPKj8Ese5Ah3i7i8aGDtvH2DJtq9+
MFOZhStzaY7T0gWzh6HFB4TyM0/vqzxPJXwBq9yYot4MLHzWmYGFDvFWmfVHwQ+9WB4fmh6ogFkn
0UXKSgyshfNyjGFXwaR0XTHWUfLV6wXmUWrJtmwTPUnPn7xLeRgiWlY67eKNZltdokh6KKgUGiUX
na47yo3IVn+VSh+lTGI6NfHRjByNQcfdR7+Bs0QHbTHO0dnRtF2GXH7sui+3IFpUnpDDrYOc5MoL
e+CfbJIdYvFY62twVj9ad7tIF8Bbq4u2IXtUxdjazAClgE6HcHkWAOc3T637eqHCT1iYpfhY5xqg
+DApIT+dhAf+b/TUOVj7G0dj37lnyHQSGxH/mDh2B0qA3cLrzTDoqwxBSveNJ62YISIpafT27+Ms
6noyFQ+JHJ/c3gVXThIGyhqezz5PsM9mg1OrXzfj8QqdXMJM1RgHRudJi4sL5vltx9FNoWdykdI+
lOpV6ELMqUd31+0r/DwK0bZMAJ3xYQW6YOq/E5FqydJ8vHRYyiswwUsMRhSPdhQ3zjR1o4f/jYxj
nP1D8aarws42imBspl+3Lbxk//ZIAEinAom7OlzvK3gXpWn56aOh1yByH1xZvUGFSUORe+M2vC08
WYzxISL65AaGMVtZjpBHKZP/6RZS5CT3tLL1NzRH1uT5o1NIkp1yw+mLYVsRUl0Q7qOC5hDCjFON
N000Ghxg3N73biaS8Lb/IQNMRb5TMIgRnLg5Di8MtZOl4XjIyJCEE7uS3unCsD9QV1xDACEsv3to
FlL8UWSVvoEjjlu7jAkNiKF7OBobzsjztBecxd5vwPur3VgCgEUcTCcqfV3wlRlHpG3lLgtSs/te
le1o1q/hZLorDbZYuj2/4XsT8C+6kXFtHXWgvgpJUIqppy9P0jR9ROqFoxroYfKLRy/td05q/W24
bXbYG6nf6mv2c8tkSU3LfBavYuSrNsGfGbeBMBZV+iMda5IZOkS3ZKjioqhVxNaKGaaT8ZiwXTlL
jg7wUXDfqJVgcxI1TM1eOp3qghZKfEqCMBysgBIAV79V3tuFca/YU16yeRi6m81V84wRn64nstfU
gbad081LOWxcZY7Ura+pYZOix8rPoR86jVCEJ//H5bnaszyL9wcG7K96PNnkK16eDNGJKGOo9txJ
E8PFqZuFax+9IjteeoiXonqQ6Ai7iiMijup602UN/9mVlT99Tc9DBEE+tZfU542ah5UwzEXpbr5p
dnDBTMVy2X0QX1fqi1hle279npvvBF1dyocbk41rvR5PcoVIi3/CrYKqp6SfqyqvLEGP27cRkRW9
yua/pey/6M376/dEXkpwg4c7P5LNkkFo8aB4pZI8BUPenYB+S81c05rdvCq7bDTeaAZ7sGotwjLo
Netgy9I5qCvI7lAm8Wd8pzeQxJtbu8Sl2E4ofAgaSBv+BkGuTjUbKdt5BtgdKAIYYFO1YMdeGxrs
0c85jjFCllSGgfan4vgJQMVytY9uxcj6HPbAbNvb0gT3LXTEUwEX0S5xmpKFg9FlFjSoGYxEJSuD
tfLkF2vH953xhTfaNfxevJkkjzXqiIbN1yswxXNNmlJy2Dc3x6RSgv59s8c89/krAWkgmt7D5sq4
sPgDwtTAhClxaU4j36M3ixgKy1MANuQ+Lp3jFBY8N8cwRU5naF1Fi2UsQxviINf2n79TcI1NqCmu
dEkBrofsJeCKN1uTCHME5mCbk6H3vMONpacUCOz8koHeiyN/ZYFqEpQw66ZaxJ1APrW/XaR9cEFS
9nWjN6R85WeOI5l7bWcY9p1n+27jmwXTku4VLkEM/ZKZggFXFyqdTxJoUbrnX7+tAZOxYuZ8+H0m
Ub8Eep49Swsv3bKTuf/Nvo4+Jz4L9MAEt/x0Vt7c+92czXyBJD8kbQgY6ev0C4IQ50KnBLqT0bPX
DIn7DQ5NZR3wrEmNZS28eJXeaf23RnugeHN3PvbHXUajpW4YKyqMCMLJfEkdoN2NNSkuOV3Vd1SO
1jX8VzqQHdRojOCPU4laXmDDaEyI+JSY/N7nIRiFSqeQBp88xDPNUrqIY0l5PFCStXwd8eu7L8bT
mR5HW799clmBUsCNf8HnZwHIGPCEWEGxkeNb5SMtT2B1WFhJAOenBkVGi7Zwv5Js/ES1XO+yLrm3
PRfkZbg+iXsyPhikL2i84HdkwqMhw/9Zp3ZnIzdczNfsgUbWxZmRiN2I2waG2X2qzNSotlzF+Goq
3TaNChW/A2HOekDO+d2oOx5EoJX4s0tgKSfI5yJVA5rw8QEXcOK+slyQWP8z6M3i4T6RL8vAxsj9
vtRq/1iqyKQ25peITBHrqsFdqigQ3RF84z0Jx9UP/XpCejXvAwVQ/eXdyA/LUVQXm/GlwYt2aNeN
SdQ6QmeoctYOaFjhZ3rbZWDOdSZIsnyNQJoGsWS/m3x54oJR97rW8uddi0wQkZSwtyGTcE5vlVqU
dtClZ0L8fbw+aWg2QRDMxogmKsAltUWBPZ5CENKewpi8gqckSdJc4+3frt9+5RZ/64IS0hYrwGol
Pxc9JCG2w+cSf3r8xsuQ0g5uCNsjmkm6GI38EJpKbmA6cXUtRA12cR94nHDDFI6n6eUP+KaZuXRA
Bv4eIYDaOULumswCF3Z2Mq8F9HRNiI2S1df9ed1PLLAvd/zlKLSiP97RDnyLHxG6U2ZJWoZGhzGU
EBBjeEIK038Tz42HCQsBr1k8nI5whwFk96Jq792W8hY4cC9fuUlBiuc6HgWEFFo2Ac6DicYFYU2x
WhxT7X31cHkyqwTh11Knr2Q8dv5NB0bpDyBbt87WbYb1NRSsvSmk+GbrEgvX+9WrQl0DbHDmRq1u
JmVzmbFsSK4gAMVExf+EQCfro92MWJ1CUfHcu/btUVMAM0Z6PalXCnEXtH1lA988bhkh7lSQWeDN
bR0GgidYBe7PfiuJA0UJYBYmHaUBpSLUfICYJem7t5G4cdRHvTfeJISrgZc5hT8R/zoCvu4H7spS
OP7SJZVLWknaXsw2kgYVKLAx4Wki365E7xDWV1GFpCFgksAgemRV6+TxUlnuvVgcx1z/XlXL7ls5
xj5XCD1zmGccX1HXOz0pOFbUCHKbgjcE8JMELL/88KE7EwRRzHFjeQHu/Kdh2oyvByIHr5GN7/S4
nrkFxFjkt8e7x280oTvBGxKNVq/WcQ/467LD7U0mjVfoi2NwjuYg02Yx/DvfL3zS2nhNh/f8yhzo
2Vxe1Ry009vVueuPSilABXyO7fLFVFw33UASwEGIoEgPTqNCw0xfLTIxtTSHEdP5d9y8Mq31AQ6y
huXUMvvTzbxyKi2IOWOc03g/Jt3kQlKw6Zc1Qmas+F11DUoqrwESCL/M8rHs7v88BlPXRF5RMlMJ
D2ol4bsqytnL0HGh+pHKRAXgsk74T+BlakOqxkfLuLciCelFcBPY6irbkeytfgif7urtnUjpvSbq
P0ANrry1UntqKTDFESR9XbOTli1qeKEZCX1UCFuDgCUYEwV5L9LwFg8xZ7fBtutdwIUfeR/CY1+L
Xq1/aJf2n0mLr1H/Ojs/wGLNhE7x+gRBC390U5zu92cLL/4Tw+ByvIz2Vj5OxtDCpRATE/bY5r8v
ixvUJ9D93cx7/2cg+fOMR1z864youk6UlGo4ZaZi7hDXV2lRNBPRt7oWZ1eY+5sZH+02fz0N8JGT
/sSBBpWgNjlTLWjlw+DxN8Nc+3Ocvm8kIQYJolX+veTK9AQorL7Ekx2Z4sbssrKAXzvuB6H9UdxY
go/GxVNNnQmhKdoDQ5DXmDXRq1pJ6ThLj+w0HrnkR7Ta/rgo9ryW6h/bMQuWC0khvGIejgoxM8bv
j1C3K92XerOErCAhpo7w4oQMZtUOuuCYihpxsuwks5uMvxd1HChZfObyjXxmf6GavsKAxca9SJ8x
US6lUiaHCV2N/jGtOhk2SlgRZ5JxUFTBlqiBEmTht91Oec/tdMfXel1FimCRqtAnZWDHIknj6pEG
stXVqvHavAVVG7+KcIszsCfIzGtkK+EqDyKsKLuD1B+luHhlNhybO7coVlmv0DGTsTYSBiE4a2TO
5C/cwvsTz0Ozan/MYyRRb5+A+CHnZNNh6xOMJR1nBG0CP/JHPW/zi/0MuBzGBBCwsHzaGz/bUJGF
VFBF/C6NOkTNHEKKVW0cjd2m0fTyuXy89L9HtDTVjFV9sWxc13PbI0XvVqF6ElKdgYS2XE2KZBWi
YbSNiahEi5LUo42+MUM/3AJvQgi+VUrLqQP9X7wnN2HZ1KQAJPDbB6oST7WS4oplg2L2Af5rgNR6
ypc27Q3UtDxI3vIFSbacDEg6nyP1gF/6DnisJOF8zRHd/iSD1GprijC28aj+3kBLIVFokLhy8UwB
tUdAmhv77SUP5678+w3+Hz6NeF555V/icOu0sUnKbTyJHj+gMokMjlPtqy3OKJ1DuNcJK47bVL35
7EtIV5yOf96EJ+HNUwpy/KM3kU6CmO9rgoiuev5J5Tn1XUCBnIo8HuG6k0JoeEyikcbO/vZsZzQS
ZJpwm1HMVGB/n/FgqiHWfFFowZHKOk2unstd3Si6tV+QZ/QySBegJL1KZbnCc2VhaEO3e6XrZtpT
IffO7rXKD8ZLI/TZeroHjUEsLBhLuqJdllM6Q0Os0JIDlTrQ5x4fkotTnSOImj6CKUzqo5dXiVMU
y5/iRbIA795w+U+BAzKWjZQzkU2tW+/s/t2Jt7tFyn44aeiXx9rLkXCFjj2evJweEneQaUasT38N
1HIXUvrx287HUt3jVzhM+svYDzIDZbdiiHJQ5+NT9h6etyRJbMaAzryXVitf/FNyIoV9RilZ16zs
h2Lyl41/diQRuPlFyS1at48rurPZjeyqkH756TPLFsSA1/JT9GxiI2yjSbPGOMoKv6lyhCmgHY2w
QU19tlLSgvQvT5MnknSGOTQpAImTkv9Q9ig8lgUQpJ+ppMbRSEfwdiyP82QBt+/IuviM36yubHc0
OqaNlNPImZj9AKqa42DwTHIb/YtMwoltgc2Ft2loFKw09dHRmkx4pXZezOITd38e85nc73vWztUj
vqxp58llmIV3CCqQ6ykm+INkp9e9WXJ0E0pzbUf+uIogdGriK9MA5K9Ce2DNepU5JQb2FSWWnMYR
DfX9vErzSIwGDAf3o4ehwuz6IfXCRCypAAsUbQzrhF6AkPFjctG3BVt0nUxkTepR+lgZHxgLs3cS
vweJGNJEl8Fj09ccHBUJOzhKZe1zcmaFeX5l1juf1DiKhdGpC07Rk2iTfHXa1logY9/7EdMF4L06
wjcWSqa0A6pCTg9d3U8bwWuM2T2aw/8UDitrZzRtb+e5C3EcMxsWdHdSK97EgUPhtZNEZXkv7zVU
ofYIGBs5Yf8vS58z5ThWP2qNJaXZZgWq/QTl81pPr+yUTdaa8N0d6zB2jr2OvMO5wOj7QbMaayRm
lliGM0CUmDT4UxiMUIFeAmutlCg2fp5jNSIT8L4+7YjEhmKgQKWkHzdYKxpGO8gb8raKOt/TYHoE
k7CVXK7x94fnsQqfq+MLoqv8OYK1lGJ3fDpNAXCBXfvMZzk91cwRlsk9ytVVmSfVXoPSkPqrG6nZ
FG8Ffx8SwGd8cydMaasyutT+ZWNz01ZaPHmFpA39O41gYMMkWIuerudC3kKVV7Zqmg3waSwz1w4/
nB/5cfXGNzC9q/TKvlS/vhAbFNsUZF01r5+JlePtc8Prqp96ImK5GtyQ8oa6s3p02Z0YiVVpvPPl
aGbZ94cAOs2G8xRw88BanT58BEr2ghJTQIpHqwlZ9CID/2AXJTOR3mh05dwpJ4Hnmoc4neD3wjZN
N3xyTvM45i3fpInIbGM+kKjCFIGYywD37k1iNj/hFIF+Pxx3riUvc2D0iz5JdQuZYohIprZTOLQD
SoeyWwjYpw07kbvxnFcuwkFle9B15ZS5IkPWYEXne1ou7K8CZ9g3uyPK+ncrgV17R8X0gZ+J2Gwl
bOO7Vmlgvmm0dBu5aVdxDXJUZ7yz+0Ju3fgZb1ihx2ywnNl0vMfcakbVDoF9jxe8j3wv6/yeD+AK
MB4Y8etNSIKHUTv9p2GRBbeSJZ+YQ3ynEHuopE8oaKPirOHxHBthcphgq+7a8skhkejFGtMHPyWh
FyUr4XBfWrQ99TKACZJIkaXJJQoP7WHfmJpW15tCrdXcxWBqFfrKACJR3l4O3rebxJ9egrnv5UYc
F4aB6OnipzmtstFXL5wpyxm7qa7J7pgA3hwxBLD4KtvWe4mWT7/WS7Lv9P/MQDcQ248MUrIwalb+
4DiAfRxDX5TPwXQF0uNg2u9waBIcoREWYntmJ+BFJIiYKc2HUTD/Jn9P0+W5n3m6aeYX86/aTAAd
6A//M8MHiM9qi/eXqS5CTHuDPOZmhnz8bPUig7y7s/Zu72akdamnPflMSMY2Dzym8LhBzH21g9tJ
HQ147q5sRwnB6yCspza8695U1Ts1gvFPWpqnQH9miYq5NXrP0fClPbva02ILtFeqQsZjOoyqeIy2
7JCJ8yxaSzsQthHoUJuT8blQcBA4m05tBNkmWrV3r1EzT7qioSu8Z+9hyCVz+Ol28TrXfktu2mZf
5d22VoS+ZY3dse9gvF/cU+s0MbcCVU3MuDyjSyQ225YsX3GffG6O0fRK4mH0xN2zdpTVxIj3lrcj
DZGnjvijxDoedMQX8DcPtvlfFhctxHlUUwNqlwkDm1oBRDZ2A29hCRX4W7ouIxBTtz8jbwmtWRDh
rpTSRzk5N1arPe3CRcNQ5zOA3jU9RDjvMVmsO4xRZMQ7HDjkArjVC6nQi9wMCydglQKrveUxA30w
sK8OD/1o4Io6P2GQH5wrSd9ejz8a5+n8g8KjoJcNlQltQ0+njkHTxow5+B5O58PoUmPUL0btB2Um
yKY9WWC3fAIRTzpWaMpZ0JH6GII3WK+FfnhS+5lPBteNgwNoLSzK06I5y/6ncogthJjftuyl7fhj
PXAY2frRTbwzX2ysBDvfmPITaMYho+cLSKGjUSAOTgVg9T8HkE4Ds9yMuuGMnUw3GFLgz0miHo3/
80creQqhevMZTDSQqf4FDEDy5rMGbtuco0pmnLuvwmjWnOx/HyH22k49UB6V8tIo5ni+7swzd/sq
r62IT3yz91W3wFK4hIEp+RAkLNVSQNCSaDyVGwh35W7JFT29BWViERS8Tgl8SE3EvYRP16hWgmpl
H9wEYhwZzLCFPOW8JU7L94OOpn2ENkrjBmaIahMEtSIB+zw8RTiVDpfPShdsyv1XWwvL9kPW6zDT
IBY+1gHJuxMrcbfyO6PoobTaPZCW2qi1g1RX2IuUsTBQnG7GdgM7cog4PsgUCqu4iTeLTux+gyHD
rGs2uC/zNKwX5K7jT0L8Y5L02LcdW2/wBTmpLxShDl2nXiQ4UXOInevARFPUl4X4PaZb5gbCn4Ii
rv1AcVBL4/mE2m3p8fhgK/sXCBtp6kyDBRPaSn2H1HiSm7RBJ/okTqhvtCxg3Sk3tbY3iuEv0W2e
4IDBJJAse4FlsjMl4+ooy04sE5sng22EyGeHA2nybJEEgOJ0E1peYgN6uOkdzPiPO5r4JbETMKLf
EFiKFSd/I9UqbDSoWsMWC+Kt6DCnWmvEzfRZOD0kC0wjQXHjHmunm2zWfNoyphhnS6snogGDcUvu
K8vz4ZRMj0ZnVYG/XhpPN1dirCzT7mbWz2oSlU3wL43it3QYHReCdTkJUBLNsMsxkdxYlZGziXO6
WdxxDeaKKe9KDoWIL5NEZTmNjeukIh7sji8xXrEus597u+tK2YU3L7uPE6cdDtoYNSdDF8YT9h0Z
9yNm15jxOc9G1+lnQiWJX7+kAoVyHb1mIumfQFr6SBgLFWUEjpdrtsQKubQEI2Qi5Qb65FEfC40B
3wqhSIBihv5eFoasTg+Jdq8CJp425uPBSv08Fy42almBjGGa/adnYFmml6RV6svrcVPcsbKojydh
RQbCB9XYxz7sKbvm41F0m4Tp9i7SobYInZG4mPC4FcEZQu8uZ/2NRIOei9AECe2SK4E6jfVnbY46
bRxHpq9b6jS4j1YAs9X9aL25u82iRxbQHDkvRUyE5ZA/v/3C+tZCsnKKOdubrUA62mAiEnpkQ1kt
EOIN0ObZRcS8otj2S+NOsh6QGXlRBjS49CHH79OUkslpG9wY38/2IqRop2NXvPg6XK276axIrk6z
bfFwms/FZt7ifcktfndRa65stq8Jj5OGe1zgpNh6p6kRZ/7boRN8dDNuXOtAkFCmfB8/Gzbnsw6i
W9mGiY6jSj8j6h2YQRbdcgTjceZP+oelA54H/GuOWIZ+5hmkOBFRWFrBjMiv6zsJ84CV8+TI8BxY
h4HUYsnP3sGEntmICv/Fgx41OE3L2HugDJ67a9wA9J5AQRuridXy0XreRpiAEA5lYxyBOWS6lMxL
5dJG05+6akN2/84J9iNehr02dqDmpor0aY7SsxvdLo0CWhHsl4N7THiWErmcJD2drCwcGzxJs4N7
ZSEcsVXXvcfIGzE1fCrZhWD249vTjDB5WxxuVDxyHaeTuIGftwIKqmw0UWlSnJMlli1fyVQlZsn3
c6mUj//cku4NqwmMqAiWhLlhUHCimDCkoN3NBRVCqmZLqYcKMSYEOrCgODMkoW4D8jIWmHEIWcKt
8BGrX9tZ9GYsYkzx2EfSC5GHA9eibX3cWtZ9rlrOm5kbKA9f6ici5Sc0/KA893cyu20W51BAIdKW
/oJ7Kk8AnjKGEIYqYK1ymwjPQ+5GiZ10nFR4gRp3xAfMyDkXWkQ3h9wz2Wodj8y8UhQEt11oD5Ty
bja9A52TfToC2oZiYnOzf5jokChiw4DHLvWtK77BTLQiO0YVfX4ZCTx6gAcJpi7IXSYmuNtrJ8zk
ZNWfbe+5AHFoUbX77afbayj4F4sbVKGSOPNukyznbr+7zo77VsWCDLOx70FVcIMyUGcCTIIpcb/q
CpMsPQpfn/GEPhiWcVYcYLOIOFc6oIMhVrAF00+0dIZW9HmHmwZ00PZOYa273dQMpdZtG8bH3iGq
wI6X0cG75zEIYQClPfRmJN9ZD0xQy77y0M4tkz7bxRa8P7B+osqdcutCNY0sOT322ML14RIMgtvP
+e6RQGn1btj6T6NZ5jidczucABkd2kd4dCdb26GBM/TIHwAggDjbwYlZXs1+1PYBxP3/GR3PAphL
p4vDQnx/c4h5i9s9D4rHbbHNhKE9M141+np36gTXSQ4x0aM686l0LUd7Zv+pzq5JYJz/nX7JU5nS
/2gFVpnBL+8VAdTxK2ZTO7kHR4GlGNPKsPdQ0eWQ+R7IUroY4U8ksvOWg2+D4odNeHBKdxhj/nYd
c04gbAkJ5M3Nw8axxlSlGWgA61wLdDfr8i2/OZZxSCroGcJ2QqVTMjmX3KI4VqvpvJq5C3ShfoLd
fCJ5FwTB5iUfimM9Sgjc8vOGJ/9jfhmAFz0iNFlfvfQ7RfcX7IfMRZDJuolelFO1obZf+4K+PIO5
VSEcgc/L9W1RuBPSS5NgnIMyCwU2rN+TLGZv2wVkrKdo9aIMz0uHrU2uN8sh0a0qcsF9k8wGLOCl
8/X+SAgQWpHKneQKhG8+oQOKApkryTEcQkCWFbmSLeRvc030H2nBl7xIawkTcnAm5BaC0JWNDMhr
eErQk1i3BrOP+tHLjKBW9WDlLD1kBtZuYVRvfTHG1T6fkTMOlhQr9FSgPftASlrd0aJ+L7WsUJnJ
D7qp+7ZIvgQ0ESepF+8rN2R7uDtNS4z/Br9EkhIJiDBykimYDZ1ACye/L4GIudaAGwIyLk3TKpqN
XfmyfYVG9T70b3FJLXj/vSCFS1be2dg9fHQCLUaNzNsI5A9nQMxZUyKzVFqUpcHA8jbDDuLNzDTc
ZLjxtpssTLpPo2uuU3mFUIYC5HlLFSgegLtE18ZQyBqLzS3AH10JKLpXe8y2CGXsYUDFgE6SiAAs
+ouWbXGf2/VcAcc+aEHcuezjkdUiuM+HeGxT39xChrD5emSk0kye5Sjpl+TTwTz0zrZ5dbtkWuHX
r01cZ7oiZoXJUpZs+Z57v5onmGpLGwFEmgG3J/wBgqBn6LpK7yXo3Z9h2E4h2swvMk303WKXtf2j
aA+frexJDq0m4qTWik4gNX4qd9hAhbP6uGkKVRGYJYk+aKRMIZLt3SS234S9fUc9LR/Qjcn4at/d
K+6F/1QOUA2t//2CjY0KkAjP5Vo8/hFE9hYhmjXADl2YuFD4HzmcySXU0x61wVnm1gwpHNpfODCE
7c4zysEJjm+r5jJhZwAetoMfJGrlGTUwGEcyr+f7FTL9eRyuCZre0pvSBtQzkuB0yDCQ0nwQ6Rmv
9zX+R2JT2jgbsk0asKqSb5bjlULtAnT48FG2V3B0TpIZUA5rljsKJ1yvHL+pFTD3N+2ep7+R/YlX
oqep8RCgbUyLkaHg8VF8Mue+i9+/nE1CEckK9ho1/nOx/RCpqJM5UoeFUZZiWfSx5+1QxRx6rhyY
qOUEGOUSYoPDp3yy5mCqbOkkPDDQmZHMcqJQnGseWnHwbyG0pDXW2LZAFneEJ7a4ZclWeJE1ZPMA
u5QGMCSp4hFK+FV/x4AUx5N/4JuHyW3PGWf/3QCh92aWjXU70aVJ0DlpC1gjvSYzxeJn46OAwJxT
DqaBwYSMsOEh6SO3jQlWS2452A8wHUh1oIrXd+WVLJ1KUq7FBJ5MZHa1LEJDNF2HCobZAxX9DqZA
9KWxthOUdkSxOAxUIZ/6Lquas7Z/9T/K9C49fy2mCoxC75j32OhGSjpPn41ZKS3T1ym0gq/jSoHr
6GfUWQDkUP5m+dotMJpPm37Ui0Gj9hpdQQVC7piWAEGMxaxb9x2HCurpkUi32agv/gtMUhCARfzI
xB+e4sgVOH+XA+TrB1kzFE86hhxcY2ZAyIcG7RIZVMzv90/tlSwmMgxyVshbH06846GPBiZGHvWT
hGqyGRqqB+wNk4gy+97lKm69UntZz+mo1FgQ7ln1oEG1t/jNuvSJckTczYYlKudHvFinvrIsARfQ
5G++h3eQW56SLFkYtGQ4LlD2aQVex64JCE4IlpJi8pJ7aO9Aea8Yzqmh9ZRGakKcgQNUrWyXExHR
IIPNOdrtZl1EmNDsg2qH2pZUcFUVTP6boB84PJWGEf952V4MZ9FS6tOIPKZ2KsmOUB5zREmBtbzU
LJCoZ5qREzjC2nriADvEOLj0LSWlOuP1I/btGv6fZR06xCmE933nbChG/sPh0Jwu7xI+VSEI3Rap
H35iZc7OduRCh1hVR351+8BfseGF1NfYYYlkNajVl2IOfBYf5aWNbA5TtJP0TRE55NFLJ3AzNtiL
R0qdRLMXUQPjhSWUMGZLZV+WibodPdtFKzjOipCzoYpAs3KODocjeSV3eIq39SaapRUUish8DOmK
3vvolHF+gq/xVnr3mUghggFdEOvI87BnYmJavcSVqiHCRYBjzP2Vsoa5StAHqGWt+lMJzYtsZ7cz
SuKhbkDKQxvizTHZKbuuxpSHAQa0ayvrdDqihx/QB1WrrK5DzYiIJne8KQnC5oLRhsdf8eq1KQPj
n0pWT2HVyz11aSreI0spJjB82RrDgq8WbmNEtdfO9yP0+v/i75rxd42XOxLPsgqgXE0OzBVmChyk
wExkoGVmdZf3W7xXygUaD4ABO0MHnrh/7BwjnkQjacC7UK4rYWOWcit0OO81R170Ulrl5eZQU2NL
awFatyqmWXhQG0FwtkT5+D8KQfKYA4tJSNRaNZQRgVEgF7GbmDWrdZV6WssskgyGYYddy942dMnQ
cyDP5i2Gca2oCZtlT3MBohlMcsn5QBYipzMF98EBcfWF4sWxB01DYkXguTunmrfep4xpYwTWc1f4
8qWImJhr8f2cSfOXvxWYDTs+E/uZB5+3eik3bsm0sPYWFaYY0DpIgGs86Y//jDMKhWZBbDASrIeU
WURPigBefYz8k2iIW164FKvgdW5IjYevaeOrTFoxFzNeYtZIkYiwh1/vqDXG5JLH37SRzn4YW9bZ
0y49gQ2YkKv8+bUsh2WYAfvmjcmN4ps40in8n+WaBwC76510PTM0wynyjq58Vohhxkg28/OoV0L/
T69lWCE/g6bpK/+ZzXzYtWODnMnF7Ke6mUN+Nci8X+klZl5XJnC9mZIL4s0RYxFGbZmy1iZQb8TB
QY82YtF81BksCtxkWwPVrEfmgNYBfbW3MSH6RlD++XBK/djJVjZw8HVR7j2L0ExQteaqmUto6rRX
3MeBGuqDnJrttwisMdmOOOtvbmkj0hae7Jch+1CX7tco5lBsatOO8MImqb0vBbLKhWaG6o+zzjrJ
pzFeTwCzDTRx8+aKrRQ1SJfpI2WA1hxtm/8SFZklnM3kyMqARtiI6IgDeMZu/zBWB9XEYGbxLlhQ
6kCCV9fp3XBzUHEy9jWXxIrwSg7G9BJe/qM/75SnqYZOYzdG1JN21DSR4jYOe6tzCpeKmml8U7bs
VjJjfsYzJr3PmVrvXfpDHvXiyhLy1qKZ12Rhepmwp0MenNQ5+SblVMio+kYPfl5CwKxUQgSRUOHJ
AhlPdokYjIYv0h9p4nESyN7IE4OyOXcird6I7hI7W1TekRkyCj1yinn5RZTrQuVAqDrviRQJrTs4
6Bqvi2vcpciZjdYgMu3Rg55aPwKrPOsxjJjISFkyee2wwaRWjF4PjbqUdGNMFv/kZowbBzox7l1E
fiBAmorj5YqzljxcXDOQngVN+Xv0UibGbXyEiLQlult7Yszqqjm7PkkD7MG0k3mXjfHKpJHJrLNK
2gxVmEMmOgEDjEUbsyHakzLA39J/Hou7PQ19fPjJEbWN3e+jDILXKj3ptTNLTGZGm7Jz5Z2HYUOk
WEVu6qp1OK8si7UZ8JEn1CG85bFpNNYIGKh6swiBJGZQpEpxUzZsMulnSWVqDLZfHgyaAW+fsOJz
4HrW3zBaz8xifs5WQ6AUKUGGeCScGRewz9iDd5ihcdb/yLAgzmmK1/0EimiV55ss7KAz7LHeyq6f
cfAK3QdH6XdGVJt+vJUDJk84OQvhiK7Jllav+ZBsqFGb3vYjdv2d6i7b2bH/IPpuGRhipJjNwZXY
ljxKtNT2QAwtTmZmhBPI+U+7swHQf/6x3JTQn7354LrQPT+83ld8iPen6EJKXZ4liF74QyOYO1V0
Vu06SvmRQOvw9Ze/wMqb3CO7jtGc3KbGOQsgxmzgI1jPXgo4yShRhd9S5Oqy+CjCc4Itcd3Z99Jv
UhcmcI9JE4wKbvTm3+xbO5wT+1lN1n+LCrxrz4ztTHVZ5yWUoZGnFh3HzaIIKZHqCSlrWvYQNp/+
/oHXJ/HF3dWE34C8Za1jwfBciJPnV5D+/sswSMoVKgxzIARLcLhsejgt7O1Q7zrOvPIGkPTX6vZn
4FKcYmsf0D3qQKHPiFDirkXL4905xeyz9m9WPb0dW3flKlLumz4QLw60f9HARQ8BYNDmf1Eo5qH3
qK4jGTKstYZ8FF7nbIfEMqPYw3JnrLXjatmsw6rdkdTz5moO31rzcxraCL/9F2Bio7Ur5ZRcmobI
Xa8BZX6y+zEjLedg7XjCeU93bSfIk+5UFP4se1/WijCYi1Q+4C9FlAd4+Kw0iTjrP/7pOhhtoNiM
MDi+AzG4b57MfkIMEONzz6n04LiPNwkgePAZS5P/yxYHa++exySmlf6n/+JQs89v+6FnK8iBhGOC
5zqKnZ/v/RyUZMLRvyNKGzTh4rn9Eg8foMbMcolJCEHFXa8GUzboNDFYhwkbaNM3vAhtdOGDLH4B
36NqvP/qiTC5hCKweoUjHOfqubQShWn39Xk2DrZvLKWa9kmq5z2HsSKhT/KemNFlOrfTWkAweoYK
wWr7AdAkn2V1ZaMiN2rfteP8w7tDLlgOTYUxfIhv4Kfl3VQr/kObJM6+ufJKeGkH/KVkvxTAgUuo
9wcCGHi8zJi8sKoepflA4r7FYQT2+79tRV8GvKBhvBwdp0M5arIe1ZjnOC9qaAW8VnDY6vgcNjz3
HoQ9Whb7mW3/VPcbmKH2AfnuNN1MHF7XIGHO7ZFW+SIewrXz504sPMlErtuLAf/0HBnqm/r3qZF9
FlDJr1C6YIMD0/djIKUHBBluK04iajR2hcebudeGBFOxa3k/f4yEk+U+dXWjl+1Jmx55AP+3HKA8
hZgcLCIOOX6iDTtEv0rmMOEoTnzYFR0Rvm2UB3Fec+hIi29qcQb6XFEwKBDcdLUrgE1GIGqnf2qt
dOh9gOxoWSKNlhSMcObSPA/efl7xaUrfaOzNu3iB4KycIwECtRid4RBmrYUV8rs5P8lmagpa6coq
CdBZgQEJ4CMnp1Rmx2JjJtnLRS902hIU3q3oFpBltleNRwDCIzP8gCvW7z9Dpnq/4an4jytBUYLO
0/oAzOTLcW00JWmJZciVPxBAu7I1CoSCPQ/tMmAg/GPziz/SXzcofjOi1smH5rMuaRcMDlYKV5D9
glqJA+VziG+/yapbpd1Pl9LRrJH5YBicxKjtXX/BfGCs0MFl1YNgJUL77J2W4OUN1pjUS6L7Qgds
ANklIDeFKXTswSCNse2oFdbVWE1SvkjoladDrEd8Fyo42xz1J8J55Lofdayb5f9TBam980NE0BkQ
ECXN4Yg/ZkRtLYDNZe4jUglxeEGqH4trleCJkibfOvjynv6QCeEFecUTY+/SjmMzTXjtIpr8kN+f
CepegBX43SvlP2rpX6JrXPnB5lYziV++X7EDIbhsg3vPoeAaO96a/hHhiX9s7txI6B8coY2EDZNG
eCAzSukCpmTnc/rqOI3Hv09ch5jUJfejzirwT6JeRPMtfeGfK10KjwnV4pzT6creCTC+kRjrazVl
igpwzpwEAZhz+ACC1Lks0VhX8zfLRQ3pZQf5n8jtnhFWZyssn4iir17RCnXNKJ4HbAqOySKGwfwj
dXpj/0aYbEoiM/MxRwMQFdvkUiBdb4iYkv3a39A4Beu/UHdatDDk0unUohJyRXoUH58cCjTJNkl/
NmcXiwlWBXtjfrBOqEGgd6qD0f/ch2IH7k6rcj2CUR95XTmTpGU2NTkgkca0F7mZw5ZNozWjRbn3
QYiBo+pVm9drOOJ43BCnyXx1FvwDrjUq9/huch2h0a4Jui+GPGCxpJIjxtnGZ5Xjfkl33Ujbstdv
r1pqq8mZ+jZrrfaRItkQlqE2sUW6WbQ75ALNilqHQuwsSOSovPCjbe+UFAjHpLfy7oY9v1OtVxuQ
P9hc4eFAGJdCDcl8fD/qNZStdqf6wcb4ZsPRdPBhQ4eHql7nfao1HL8XrTnsuNhNLegGmo4Xn/jq
7CcDJjQKZJf66Ni2R2fByL+3hCxwOAN3uIz8W14Ae38g3P0Uk5tgBk65jxT/f2kGneumc7a2wmbv
ouq2nhDgVZFk7BLSr2hSNCREMfxJeTOFLaQ98pSBrgiXITob1c2ygRTKIVY4LPUrSDjCHkAORFd4
LcAZq6s+bCWyCgbFNPOC92+ddvwYQtnTVLD60XXrEknCn8dQ+e2t5Nqh9ljDFd0dYjkzuKszaelN
OVUtigNoXE+m0Bjr1nKds1WcbyIDi9B03mYkgSycHbGxupYg79TF070Mp5zfRLovorTz+3UJ1kVy
//Pzu3B2sHEYhhZXd10zYfpR5jpbP29Jg/uBKRsbtUXlXg3BaKxM9XyN97CCwqaoyX0vEPyCvOot
IJ8pmrZ3g6cQo3KT955wfY/xr79jS0rGu2ZIaKKOGEBm1lTy/SnqDzyatDWmbGGXl0hhsU90BqQ6
1VSCL0Aztnomt/2GInQkJzHF833LDKvbdwZKfIGZhMhpjTcMKzSgUOVju3luwOADTLZxNA7T+UZJ
qgMfHjIRiSuTZ72yecnEs7Edtrrb6GDQeoRzNnQ1L8vZj0mrtmuOXSZmSbfDbS+PYRhysksm+P/W
16mCDIlRFKU5ZvpkyHOgjZpQMUKvGkFtVSgbAzeNpQel6qrTERvgcP2NI5FdOfI++tknVQDmp+Ua
SO/QJpCZBbgV47ezyw9t/JQiGLxCpl0NUOO69w0c45q5wSoC73POtWpB55skpyVrGI3mB3QI20jt
DoB5Cxd3YPO8xRagL13ZHdzrhP6Q3ZJkCAaJHbS8B1S8Rop/4twAEJajQYLJxAd3D8c/Nn6B3VMD
hnPZ75JK/hzc1PCScNH2xQuYEra1sqpqExj6ipzJRxLnEMmwV5L6vccvgaGBvk2hZP7dqWRxBHye
dHPYoCtx6G1iEQpx/VM7U64VgyQAmPaA2ffxGm35uZkxYxW1zbYtBzsR3wtbBDtOcpnkR4DppgXE
baIFlcFYmi2LK+rvrZtnhXccvUCZQmhEJYB9/ZFbv3H44M154I9xsUAEgRK7QhcRCHRXaWE3lJiV
od3g8Bq/BkCMsM1m81VhKH2eHnDfXBdDhDAsHvYTgDvtEP5s0qDpqRWhCxp6WChfmmwDWcM0M/sx
xOTrW3ffxcN98rM8zyasUcdPkrBGqoasdmGp87cfNx6TVjLhBl/jMfe8YEaPEQ8OP7kl87SqQtF/
rR6Y1896E9Ua3rN9YvwFbIoyju8l19GmI1aFX8S434/Ai0Y6XygAYE0Zqg1OKp/nPZen5TTBzmQE
YSKt8OIdF2FuInCYwLZ1XrjMjFWHsor7KP+SiBr5uQBIE//Lc+FttgcVyCNWEsf5LKvpVG+pjQTG
4MzxW5fd1r8mJFJh4QmH70GRT4P5My+n40hdU053VK9r/ViqdzReEMCtGWsCKDzeR/4wBPRae6ZE
fhboshUPnEpC+L5dPSsK4ux+IfvACcoQ6YeBJ6gNm4jdoWv1+5b804oaQmic3naNushG4CInfMEu
p0Eyvoi7R7k5d5GGg8iZypj26TiaC/T5fJjlQYpe/Jyea1Ij0j0lENcDeL1m1SYMOUak13K90hWB
JqvtdsLXNjKIm/ZucMfu3zqYOvTPhb4Gsn2cTyg4KQEP8hg8EAYtXVeEEuwUc29xc6Uv90fG6EzV
Zp12cYf8GbkrCI/x+yRrIhncVjG5acXQmLrwfbrH55RwXsOAnsfO11JA88hChhhLqFFhKKTG1UWN
xNs8dQDTC+y1kczLvHH75kyCuWwH6bPzln8Yn5SOZkjuO9724vPkemvW45Ez4Bx/l4n+X+/zDnNa
JiH05XnvexNLhIhJM7v2pfbHJ0VcPuKOKrV6R/ygts/gxGdZI0YU0M+vU8boPJjREL9ryqtuROHf
J/ElHV1FtYMVC1ZVbOVWBV3JajREkWNPam2/sGYlcPiMONmlqVI0YvjSvvz65/f98fpeRRqOrx9b
gFCQ1QLx256zAACTgV2shfzS6CY24NH+5gQADhykktkqfxJuJpNDGSiovGPQdGUUrcUUH/JLeFXz
CzuCW335YG70Bebk8HxilBjwCHEb4iekNr9jHxboBL/SYfa1FtYQrCJflWYcAG2H+yXGmsDhqZit
e82e67oRqkLSUid54KItxKOl+2KXknszhe9lt/oyctkZrMpBen9Tn9mZXHzyXp/tCJv2A0TFht6T
HuSqhwWO4bGHaVjc9qXaykGjXl2/ofQJFioK03XEqrZLZE1r4jjZ4Yd+mOYgBV8httb1F9W0Xxts
AKXL4/Z+2Rpi8o5MFwkPtkriVpQgGC1cMplkep1b0iPB9iuNJ9B2kJ37YLzStFIjEZcxIvalBQo7
Q/+d/SjO2U64v20R+rWAL/A5zculBHwo162/Nv5gJ/nOBAOWXLG/IdlJgOFgBSN3NFbq697iQSNe
a4Djn3ToWAJ151cHV2AADAzA5FWXkcUyTi5vn3Ts4UWDt1snD3mR8TrATNZWZ5h3KPey9w1Bq6kw
12aOzlemBI+X1WH0g4/mbtsvl7FC60ow8Za/umgEQQDmijN40u+O1zEpNaBPvv4/X02XWKDOgkOg
py+XSf/l2iLRmyBmSkiNifPN+ANPO/jbtc4XbnnTca0V7WCx3cW87bmqzJ4jLzK7asbn2T5203k5
1I8x359qnr55M4PqQBHJa8L/0tX7hH21XsXbWVgiQjS+BCE85VXv7/+/APXOVPLr5ix/nDzuMUpL
650FW+N362AZ/FqpwRZpesSrs+9F0bnZWFb28B2e3HjVN9OJnTLDHiTcPt4krvf0CG6wVh3UvCb6
AlZd96A2LFBJEWN3l7Hj7si0Z68oWQtKHsk+Nk6x07Oumsf+pnV4yjeEgPNE8JV61mFN2k0ppPak
YRLF6xXKX+KozVY7zKx9TziEa2+2kqo8SPz0NuRCTbRxUZAqO7deR9h2ZSVMq93XPGGupqH1y4hg
T+Ydyl3DgiJIlvDihEH6xbgzV9SBxdIONcJJ8bz+cQ1PDhyfHsTvq2hNI899uB83yaXZNceEiNF/
uuDubYrjI3xx3jpGTr40TWYO4OOW1he00Vg6hEFItu7Z/BrKISzF8xPIFPs08Dkgw6XvlXsFCFCc
/SiN4Dz0pTY4sAuJ7xUKx9x50O/P07LFqbvH3ngZrTmE4DHc5FJsDuiHM/yTe6y5dJgMfFA9CYb+
RuM/YP9xUz9eWeWoMRL+1bScEvXDUloojGL9SI4RRtWvQHBAxfdLFg8JlTVlYkExIf2L8yAVP+gK
ywP2pyh4LkMxZIbzSF3lvx7iTnJiv2mJXRqn4kXzkVQTdhFd01OdolUAtTexiuS9XhYAZK0/4XGu
B2oWFQBUgOQBpOBAtubzfeukKcSl09I663oX01q+NSaLXU1N7zGsybbwj9Qw9PZydm9H5Gv/h4cE
aPEFUVFEahLgfKmdXpIKQW8rAABXy5LbsTJZ75gWGl60To5gVD9ibVOt3Q0+nFRUk2msS+tjXYAa
JDrBJYSVwpUOYzHDBZrItsGcyHbMzcEGxj+m2U6IJTMEgk/uOtjLrSB0SP/j9jOlqScb4gOkGl1X
RnrFQ3sE5zyzTzzO18SjiTwWob0QTGosqAnnESUiY62LxoijH1rs1twUSzgfgIkSUNaIQDcYVhWX
sChIdsWZiDtsHqBImdbQ3EFpoz1ZVWH+SkVdza/F50qIfD8ZD2GUBPyDwn6jUUYMtWJwd9SH2YNb
LjwQbSMXjiT6+NMEPPt5y6Xjj66bdxf7N3SQwdhulETOhyzKepNbeuO+LqeiUtGrq3wKG+BrCDlo
qphyFFuS7Lr00yuBsz16569kL4PcWmDOWamXaLeCyySI++T7okbIUtdNHADSUIShyhtQcN+P4KTA
IS1BNsQuypFNwzox6YuN/Mw15eeeG5t5x07nEu7Hn1aVhP6jgNuhWkKwUiN7gJ7Okm2wLSckl328
DaxF6uagoTylN5At4WbvVfU0seXRlGTRfiUACGrNIdmHRmi+Jt/hmSQnWoisi+9VkqU4wWNhXF7d
IMDP989Ax7jjrRoUMxj7LC2iIXPU0Uv66ggD2BvWHb38pA3O+NBqJZiMKwIeQ0fKvSxU5sypco+Q
P1mNeKWHOucsf662hFqEfssIhTJLRCPkGSVsVQySxTJ2VzZmQ5aaVdhKmYEc7ABTXoOY3HEpUyZc
kQf3wJAUEKmqaHgqvmj+jy6lfVid43NQYNUP92wypzLstOeTh7a1cWhaRPysT1cQJ61FDLUBVtkx
ImOKrpY042IpH/WloFxRiv8r3q4eMChwY2O+h5067YdPJLo4Mv4EjNvM/wlZrH1o+55SY/1903M8
G6+MmW1cHykhY6OtaJui6E533qLFpp/Mf7UBbON+tvGKIg4Q+pZPKK0VOm8BqZzyBfZr/k3uDDZ8
PI7GjO8xAo2feomZLXq8f/y9AGiafsDP4bQtDKUC07pFTFar2ft/QhcsIKE5/5Ycen0HlrvIRuGk
/Fm96KQPrcr4Rt0pg6uG2DEV+H6CFechLaxbEIAnWZEGqODDn9rWb+GEYbm035FzrV9u6vMc6sX/
AK3jZ3dXiWfV3060YbnnL7BEqPNUiBRUWOpCF7ioc28o7K8BHEYlWbueHc9mh5GyoAlSsd4RLe1R
TrEdD4wv2It0NkfMUSrFM2aqdacSgkJhbgbZXvhPy7IkgUcuHl9jhJ/NuOmuVWWoWAfXgQWSw+UL
2EVOnW9z2KsseCpngtlEYaFQW2YLPqCx+6p+z7HNbkh2pUR0kCukGato6PmIWr0PTexBbYy4A98R
rDZ9LW41YrvhGsGHsb27bnVfOjrtooGPxnsDZjngxjn6JHZY9tU7DjLNEKi7lhdEe8cCy3k+hPDM
KUKA3XmFA2tT3TCjHQv2F3Vr//xCBUgEnSZeFhhbxJulm0qA1uahWO26QJCKSDafjBqTyIchQbtj
y4YOwXwXxLV649hLowV/w2iXm24IH/Pm2EhSful6hqSlxF5gdc3SvIvVTJtyKwIk8Ih99OHH7TgA
IbgI34MuvvYbK/QPk6SYHsTGoV9U/EuxqcLcUD19treCCM3YEHk+URW3yHcfAHUhD8RkRGO9Eiks
lDxDzfkLEzhks12JQeTiVuKGycZLmM7K/AkNOoEhiYnCKTB2K+xqQ1zaEdSJebzDSTchgiSbnYny
x9Y9UhGsGFtDpMNS8+AAmHenpaVEhfmMB8v0B65MyLE3xVzQAlhlZgrC8rp080UDsGaPYObZCqUw
hgJG7aUGZ6JNKWJKaXJdD3WSlnEpN66hZk7jceKEPQDypZ5qSVBPxnuo1ZveISFrtJJT5fsOsawo
4L+f/aXW/t1GBYrTEgFMkY03jh4dmGP4AiR81zWwUIJzPgHJ3Zr75U8C79/jsjdlwACvb3uv2mzE
0AOI2dqOvMLzB5CPH42mdIZCHozj8B5Q0mWjQ898O+LXk9V994i3WrlKFeAVqcch6acPwnqL8O/w
pWJwIvhM8jBJb6u7NujEHsWGEqKshD6lI9gzAnNK2MkrhKoLu4vTFnSQ9NmxaqW9aePdkxKcUsvS
9oxgSxtBxfQMnqc/Tzm3svJpkbOhUEGq6dfv/dN8AuG5HbzF1Ripz5aVw8kH/utIEbsUwzdJeAzL
4VRT6bJ6N46t+5XjGXttu/m6ZBAstEB+1St8/gUYtTQsQoN2UJIeGDVESVc5Z0kQ40ciXg6Efgkv
8WHv6iofylwFgARjwFW2ygju/5t5g0xX3oJhenWP/BhwCzKDc/kyRCOV3r5eGELm0KAyDoJAuDKU
lJslbSSI09xvAwsAqrEK9mFtChlNWsZmSiQq+TCuDo4rPtBenY47+r9BIxYlEQfUd98uJrnKb2jd
9j6GuyZ1HXvfqIACzUyT9//FCflWFGLhR7KZ4VMjniNtolbOHtkO4xNXOQd/kTrGB/y/UVeMYLRl
pmcQbsfe6WpMGZJ1kiG3QeUUrFIaD9Y6tEvojIjDrE8FWq8KsBA4Fp4I4efXU045xC99loTspHKn
/DREYsQQePp/VGi6p5R5bsaFB+T0jzaj3U69cbZg0BSyDGS+d3hdXDk6sXV+8FRsp2vRUYOOHeH6
/4gaaMptkq6EZRxuF0JYsrUxnU7SffSg9L63s66ednTrw5D63Bn12Eg22BpOcXkL1schymG66F4c
vYVHxxKwyp1QEupCqKf/gWn8SJe/OauwamEWxl6RWQb50FryRqfH+Pmk1I+5Cu9R93Magj/G9lmI
fOLbRt2HIzwrg8zBHEGgw1l6ZnoQQwEZiC/YTRdKkgV7Yabwnlz4ZAtDQY/AzgwO04yyZB1Bkxuk
PRDQ/L3MYdzTEL6StYRrMXRbVpEuCRrJlOpzbnsfqsyBmj1cr+MplIYelktKsER3RzmhVCv8mzh2
AHJ5VRLR5AD/KKW2oF5CehsUESRj3klOZw1XqYnUklfpwAt6FOQYF/OuQq1o+JjIY0G4CBf0jLhQ
O5+U2kpcj+hI0Vm6GbfXNwjCI0PHj/4lXgAbEc84c8NOguu15INlZonYl5ZE5VbnOrx4TpUS3RHs
BoiNR+Y3mzi+E0eh9esmBLNwj+q61v1hETV3UZISDUFwt6mYHBzZfetpRu8yVEy3g9GVUpxzjDd0
19+0/WSV9D/f0u5aIo8RFWk0RGX8hQ7RLGqKGLDFHpB1Tviw9d57S0vPU3kJgeEL5ex/oOjRXgUL
cNS/EaJ6h3Zq3Bv8QbmjKIgjK0Ri/99dauf8Z6yajSxWeEddFX6uGciPCyrgGVw2ivJM+WoKqe88
RsMIvNWe4/Z2mUVaO3aNaqIGTbsttRf20qR1McC9Yzvn8rJMwP3ZwsQrn4boN5lWGcFDSnlTEoRS
NZ+vTeSiViLypoX8giUYhcYDOiZClmqcFadsGp7zxzf/Qhdzk+HUuwhplrli0ZIlRVQUVtmYTy9c
qhW6TFbYe3Y3GNNh48FS39puCpgQqETQwOUh8mZD5zP0yqfJuknM85Ihs4oOIhNpjqma1CQ3MGQc
jKoKnK6csAPBNAycOg38IMsp1kjjq6UF5l3469haC5r6S90oo4nNcGin8znaqZ3VPpiDj/1y41HP
TNOTgyqtlH6f6ATsXwamx57yd3S8WUTgkyEYgrpaTh0cfPoL8Bs22CnM3o8OwKTi9pJeBQ2Ohmuq
NQZasKrrNBeKKIfhvJlgdaiaQWQXm7sMG9jowEfL/5IjOSh5iE0gjroqC5ZJLoMZg5D8EA+AyZew
6SEEfhmz5xfp76BZ+bA4h9xN8ho5ehS/AlxdoLzvhMVI1oGLFpqXDfEI2mJQGai5ERlhq8yTdNgH
BEETUdV+yfirb5YbWw+L9L9+auI3etjpbHMqgBSn3gZbnorBLUTHah/oinl+qNY9ZRqi+Oyh8QLj
O+5UOYySdQqIDGes3YsPOTojuXkbD71RIAiBFksDpWW9wtCMv9SJN+LGyDXOZ8IH8qDniXCCHCai
vONc8nU7805JclYEyO7zErCBc0+e1LVKIOEsb6JI4mlYhp9x7VeqZng4e2dQ2YV4bXjuhROWRDca
cypSN1G31ifK6/BFPt6X6A9lswMFyYXQUOHymN1od4EAcmrPNnre8503bbI3SrabZo34tB4IvVrX
nTR8HrEVyKZ+HwbEoYR39/Y4miFJR/3GoZBeuTnHHGJoHMpELBo5b+vdkPc8pXUmzoka5vYpeXw+
rApu2wGvGdULnwO9EjjmWiiyNuWZoQS5c+ZdzeTWKnbA/rJzo4iKUbzONsnjAzFffDPxo164Z+A6
caZJCK6HSvq4SfqIJhM540lZhNRGinUwlkxwUGrhkCYwMqzVYzKknurHjJTlcTtr0uw20+RGHs+j
my9zZU0KwyJT8xllaCtQJWG2gzD+cxB4ig+iVsxPO4cIAh/5ySnbwxyemSZsJRTcAHX6uutDxzKa
vIHnvM0y8Y2EDJaMxuT7fqluytecVIZYUqE1bapYHICIv4ETMqDqhriBpJw0/k5Dm7ChngvRwSY2
1RLtZjfId3Itj37xOOTVimXEwSvicrgbPexpbfbUDypq8d/VDwKfQmHS0TyMG3ypL1/fMOXx3Rzg
GDjoEqe2jcPx9pT/aD7Ty3O4f3sJfOB+Ew2XE6uZhIBOZn7VsR0qVoqU0TaFEc/YeJeCmE54zpLT
zOJAw9Pqo0UzJTkUons7ZiAB6E8mZiqUbUHa1MLz+I9Wrvh8+DY6NKttDUSrnV/SIpkyfKR5YvSI
fnbYCNtv/KWLsunbrQv29UUB9bTJZQJIUgPkWDwpp0uqBPJ3uLngj93DsW903iB9cxSbwv7RgosM
WZw1VKWrXd5FyYN9dS0wb+edFSdSe+9cYHV1D4m/vUKdJV0epHfrLQJVBmP6k9sv1t1EQ0dRB/Gx
AJ9JXKLSWzuJDTFzWbOImMMz4FC3DPo3vLdYixfDWc/buUXpYVmqgH9KpeOcoamSVg1D/X9fQFY2
qREroxDIBqHWzl+wZKERa28//LOlr9FCQhFt3U69aHwmGKVB4ZubNsXzVFb55ssJKX1b1SD2giam
vfvY2x35vIzTQ7avMERyaQuVIc0gYzIUyYq6MALnPH7J0IBxTqj0ddQc4wv7MyO511gxmUVemNAB
1mQNfBcpVEZFs67zoHjMrxb6M63bZyxz92urLVmIHHkSp1M3T/TQAsQE10t1IkYXzH7iIA9KIl+T
rBMVIcn3l96Igt5uP4WY9yBGfR9Rc1qAW5mEtmpY9Z0SfDQ5ODhm7YnXiO313ljoImvWHhDaa6Tw
YJWjOZa9ceGzKmnp9Qay7jvHYiI9yCGCucQCe9aRWLv4h8QwljSRnq7CTlki/TCVnYDV62svB+Ti
/In9Fv3I8sQSxYILq7/q05ZnRay5z1a47xBb+YgP1vsJBY70L0RR1GAOzLz+376xyawBTijXNZEF
nqyiPRy169kFoaa57CZNhdGiSGhEcol6zDvP4m9VaJVDTSlJ4d3ka2egln0QIFg9SPXarUBrqVJi
gWqN4d1PfDhxWQqj0ZuZTb0wiiqLy/cxnTfZRMm+63iF6W2Abn1GO+Hb1yZvJjO/nBfFAlEGNMbW
0yMnGTnHHucpbZCszd1Pgt2SBCBrrulhPfTaFtoTyF339VFZN6wm1dx73TrZzqjRZuTgTETMZmd0
Kv6AruIIR8+2vuKRGm/4ZR9nwXab0DDcy8OQJ3Iw+L11zrlvYAXqRDVrUdFpbmjlpKAzPe3L3ev2
xcCIL901R8D4b4y4tYyBJG9i9MsFm11nD03+cVb3QoH3K6D0bhoZfBdVlVxUefKONyF/nCctcZMH
xAzlunPcZ08lAszuURWVu87o5rCu8S0JY4USDZFIcsp92FOLhvtULxmMTHpQeRPn021a+tXO0p7y
fkd11abuMzWq9T5tw0m/PJlpIoTeUC1us5jej9vYFQmYdybZ3hY6QWe0tH+N2fv2mKMhNSaUAVfT
GLNLNL2I1XJ1qnsUKerREiNULA2yNsZ2JY4V5KLMAvbyfcRKje613FhAAPWKgHAw6fEJLX/Wyfdv
LDb2KqbzRroUeMuQq4iNqHsMa6PgaR+9tu2QQc9TR/ouE3eFP9c6Ngm0m/jHtm8nefSE6xuKNHfj
r93+gV7Irnbsf6Tz+4X3PlbUDAgTLul9buJmkJxVafB0EfdYhLxAoSoF+ZQFnlTporwJzTV8hgWN
hmHhV+qwePPQMqtNaZ/x/tze4yfphETNQ9yE6dluA3SSQMt2KZawjFhwZ2SfWEM1gYksExCFomfP
83fRAd6FW8T+wg+jMVRXxmImjt0KaieQqGDS5DbKSPAJjp5rKDbAID6KOddo2Morru2+4kPbghtt
vsxx4BrRhoTuIq8eEev4IyzHpNKUepLNhXjRJ8B5qfK2d/4E+FhyN4eT/1KmW+SGKI/uGe1yD68y
Zpeb1GiaCUU0Atj08fjyU609hDAHIEIZfqJj0xc5Uv9tTG3U0MkFVjYVGvdWxXti2WaeU5MIIJ+z
nMJFaiovNEZW18K4AsOmzmrUgH3LjhZqZkeHjLI83XFHmIBCmuShYMub074sh3J3o0TPqTCSG3L1
87AiMpF9BcgY3v5e2etr7EHUlowm3CLoah3NPE4EIgnQUKwrrU9lH3X+jMy3fYOuUm8EUy6yWDuy
q5cGBtoemUlA6OgVw2gBmPrE62ccZW/nyoicI8VTKw1u8ZotSjd7JngqaoDClB9Fc1GEOJmuhy9D
jAFHfu5XYL2cdb0DcCG61DDuYWqzEtrAXagVGqjixul0MKcs8XKmDA6TCxqY3bRJ587Y+DpSjinO
/szxc/i0LOtdSjQrp7nmp3wiOgR/LHgWy9GGZma17gXUSVQg2s+2ayKZuq53IUGfcVhMW/6fu5e3
2paB3q34D0FkxSaa9wQQkyH/kz9bTHl6/4Xs3+IfYUc40tTFrC1GCIjeOMT5d0kGuNOvahYcE5vV
FjihNSkANBckyUl3J3sjyJ1JpYKmN+dE7SYbjo9qkCtw7GEwt+2W3TpdhCd0ZGxql7WTe5pfXiHw
0VFhi9JA6m1XlAxiRruxxU/yfVLNjo0X/Rh0JkIs/Z2Iy5JmkS71czjcogemaEnuRy4x7DHMcEVK
CM2s5Q8zcQBEbhhoC0rRuxeXl0ElQIIArOcrjKnpzb9uD/8TXDuTmCvmwJSiRLkcewRGU7WUi/E8
vvq/3yhminEIn2jh6LHTMrSZFmf1dM0fU3GEWFXHwHT7Fq231M0ab3lnGfWt6/EormWqWa3fcFsG
JZV7gS5VamOxcE8I0xTQAbDLXOVVJ96sFT2Wi95/lfi+uG1SfBtGtyotAWk3BQm9MDeDqq/LDzqQ
OgBZHF/eJSWZgXH9uLSKjcF6CPmuHAyRx/YUpuiIlDLZVmNXU/cJsbXeTFdLBIjdN/EeM0FDb2O4
BodoFc6SQcvuL9BXqUClWwGOPnvlzWxUC7B7ToH6lkvkk0MBsGn2aSxP6nBdRGCbzF71fLlFASeu
Bd5yBxj2hDOarMP0dOOqdwc+R/S6j6uGub85i2r+YX1T/WdK/dN6M5EIzcMFk3rsyqAha9b0ElRW
VBB+SOxNDuFF/z3uwvz0D5GqDdxuNgCIfO+o8VK23x26COD1YdzS6vueUV6ONKKI9iJYQeWz9jXY
6gM4EyN7TLG7E6lReWKO/Naux7dJcHrfP2+KA+GK1INXkf6JUzrli0PRG9SWj9H5Gf9BJRSzuyGc
VrnGM+6wa7gTzKKb+oh0wjU60IcFr21pJLgM+ZbjXFHXnBbqnIOF3vtddVHF40GvQZ2Y9WUwe2OR
CoflVi8RNDI3gHH6uC2Y0Qs6y2zHGhFEp3qfPYqY9EUhPX2NKRuefz9D/CUZ0Kdg4QM6JEhYlY5b
1a2ZP3UCDppEiQSPsb7dxdzH1gkzJijPv4aPGuqhrSiKduH/MPVq2PNY7s5FGuCTYP1Oz0FeOCt2
X6smmoRcSAAe2R38TpzniPCwG8Nh5rlJR6OcrQPWc6KseKGMBcSky9JdvMn/wyYatIsVPWnQzcuf
jaJBhKc2XEujSsuLFpTGqwxpHETj8HTB3IZMo12vr0Nc8N8Qgg+yc+dUYQ8CPtxBGONcN7GtR6ri
N54D4oumeqpGZTj1Jjc81ruls2YOwOUHCA87LZLlaBfy7mkDnz9OzcRDqj93EINyjSGkhQqWzfal
kFzjQUgc88dA5RaB89Xrgq1D/6xOpzIHjCls9VEjkfZ4EemUWMAGxtaTTlJ2XntuJteOF25TN7j2
nc2ZWMAfX0FUlCg+ko45AVWNwtNiHChH2hw2z6i2UyzUJnuJpsIk2wHwqSz1og8W/rNgIiaM7PhK
8z6EBpLvrtBay/L7euoVEkytnM2xWZOAuWygMcp/+J28Fv3H5O3b4ZqREYp4VxHFnYjv0M4kdXFk
HscG5lUuRIsMril8HHL+CLY+qub4T3LrOv07vc1b3wLRA29aRg1Rd1WVgmkrDlCZSBzYxdOesK/Y
/7fh7dbw8PukZdG3jBh7SofUIyC1nFegK6HGW0HyMF50ve/H2nBfdpHo6szyeM7cC2r/OTLqUFV9
+bhuEQzpQ6Z+iMdeVxoNvIOO1jvkxE8YKqxUnlAiUNEjNZjAWQlng3Hsd3RtDLIS5fPeDhKqas8b
x92qFSt62sQwrA02mZMSIHgFuxw7DBa/yqhTZcqmtnGzayvF7WvrkVDgWtXjRJQpfvKjVbIEgNYq
Bp2MzZmTFcQHISPGGEZQFBGVTCTYPji1rQCXvtEG9srEAND+CgHttDlDOYVYuDjJEG7KObtEGUtc
F8C2cPYR2LWe0D8UM4EtWTFQArRHcD3rohjNKGJ+AfOwC2CuxE65lS9QSp0CIDQC0vGspZwnqDvC
HaAgTPxiFwcU86y4AXITUS5K2PZeakbFwhvrDbo6NwqFBwaV6XalaUeNy8xOnaFo3Q/pdlwrefDp
6S9aAGnKTPfY9NE34FgHxgeuDdQq00H7OeWGy6JO+yXuUr1CwZrImsLqMnoAhvQDlvwQTrFhBMs1
1E7392gM5cLLEBM/B7LmjlcUmQ1DhE7+vRgHSXhWA3Ir6o+P86VJP7++WJaxQ0kVOvrz5981JeJa
BpUomyT/Cqw0vus2MWx9VuFuxSiHqc0XzFKq/c3y03HOZus1e5MXcOvE2nfe1wqJauFc9Os6EW3V
bI1bWbG3rFFhLjmosawQJhTqr3TyLuu15x8YytFJJW7HmeHosIcYaxlNakbiRX8/gjc0fqlsPLNh
IHYt93WMWszKEQ62tFoE3zrYDxTEdCApt7dsiJILjPrhl/3C32UgmiSMdXQFrH1+tF2UTsyh4hpu
DfWDZ20m/OeC/bbuElnWvi8Woa2OlOdRa6yAvQnZSFc3Lh26To8o/U5Ne0YUU3wvHpbZ7iGcWuc1
+VktH7A1de2AVFMIjhpLHO1dQD36xikLjdii0FYBADcYXFwZkmJcB6wbazyhSWYMv7ILc1u1EbTF
00cO4EVwF55KjgHnJAmKWt7tUUoNVj1ZY73JVMwOvVf8HrEKc6NRdlgie3hLexz7y1OA5hlGTHlk
TcsZTIKsKP2+ToCR84qR86VZOyHFfV5kBKy+2kr7+twQHiB+lOtprYAL+ajkKjwIYKYBQnjh2CgR
WicZ0RelOgSbZQp3TAcVjC5UzE3R5fqq8Y5nJWibCOZQjl80LTqQDHx0CDsV0JAgnDPR2lJwTowK
U4QHiCkbndZ78d9jUd0yJlFA/+QmLJUgq6DvXpkOPAAlbHIMJCENfTkr0djOPT0BkXisDlNJ6PPJ
0RSZ3yv+kKDzlAdyVm9xlnXp5YxIt80ZH6nUI/Q1/QqxVrQzpZ0Skk2soPDqdlyDzgnboqv1t42H
HpldCXtK6F/yTupEFBijAvtAcOfNVqsSHbcZP2SJcDzEZV7RBPmK3ongaNZaIfihCt4RQlnNMXWe
bin7a05B+LQLgaGQkuuhqT/aHTJPx9UmoXvB8LL9W5huqpKio9uVBJcp8DqDf3ZYbZrvOk44jnYh
ygF6PVdjFj8FOWUZuw47E/9cMNMVrJpATfSAji1Lywy4d1Equwv30zgO5S0JY7bJL9fDpTWX+nC/
cq0UHBMoN8YAlUO7uzE8fIP0oy818eBfN2juZE8+Mo3kRu1OhaUAa7Zp2vnXVsRa720OaPXYW5OC
8BuxCIJMTlXgFx4I5Qy2jt2FYHUqgMjLWw9L4D5T5T55eQ2ywtEvyU+46RJbiPIzxtGr3WDwVB+M
NdSWpYAjJgoNPaHor7X0b6w6cDJOhwc1DWcDrwl/1ufRigqyzlInGLbRf+0D/4jbmU4ecqnsLd9I
oMTZCVa1BPHD0dPVl3AiQ6UuAUnQbfCD6S5QtGk6psG5rTo558v9ppGL7V6/9xgJuLprOUWfQvSC
8W8csUrLNbx4ghzpiubwrvENIjuasU2eSb9pOqTXDmlUsYgG+0+9zjydyb8T2ycXuLeci6GxqsMK
rw9GYKgHKAbB87Lp58JMv/bvC2TpDuTtRyv2dKUDWyPAFyWWPkeF5VDPCGDqSOqDzHfWjlYd9RAr
OhU6Ez93RbmjJUG2Y14SV7FNWX/+ASE7TDF2skyoa9YTMO7THkLIeHbdouSIrDwzdoxGSUv5ZtZs
MMzoJQCWj5hshqCyiXQte1+r9TVoH3aiY8ns3tEeyJozNIW7Q9gN1O+GGPJVTK7W6E8fBSvqd1R9
9CgBklLNPmqposmnvvroXKa14a/v6r+ChJCEiDXkP5+10b+2Z/BZORbgqOKJTcLso8t94AEt4BKL
OF4eQ0gnTqx4WFfns1KMZnzyEvUagwGzdRu+REajU+LRRo97j8jelf4P9zzyVvnKZzyifEko85qt
b/K4tN0rV6gTRoGhv7c3VqeeZvK0WZieV5k1vNXRDuATHs59I16+4odiGYQeNHz61m5usZ+oKiqR
I33fY1Xn1Z01vmG7KmmEwP8roAT/YEY8jf/v557C4FtlSjGZJcTkLNfCtWYxoLtvdxvvgsXAesqC
8omxtxHstFZrj43+uRQFv5XMLblHq6oBhg0DTakztEgWN20cGzFac0qnqT+YuEch9XdhKNC7ZH5p
18ZelA0pC3QHr71ZgF5lpqp4Ov+yFEcAuEbN3IaAFLiF5Ob2eYSeq0Ogte1CkhSBEop/+/8Dkjpd
cPOkvgdhl+qLiyv7vgsOYmIAfuMMK+BqQS/aZ6GZsP5WOGNzI6pGb+lKdVr3OjN0F38gmMTuxIJ2
KdfiqGd1Ad7FlgaHIUWAqpaDxosxkUzko6OxcMlh9maS7sTeKgN+Q08cOCrQzssn33ocFbayXvYR
tAH00aaXweLToLNPfmaH88srz5Nc2GM2yKgUa5YDedhGpkUzUtWlq9HSml2Z2AWUW/xvpis80iY9
86PfILXPQM5mzfKFc/RrOdBsmVqoReNy3tZjpcdHThdvz9QOwazh/wj2yEJZexzFcLIrFL799516
YydEY7lpmGXA2RIzDR/yJoqcF4fZyTWLFnqpvQZWWMsMWMs5b4YG20V+6/hCPxfa/snpqzzOGjaE
3kpAJZol64URRycOhkDo4bHhHz0EUUpKZcCAsOVBdxPKVUeBD23WB3iiTXmf8j+u8FR9zOo4W8XZ
MrfNeNO+/J6vRzJZA3/DMHh0WuADJUD9F0tk5n57Y6m99InYCPwY4g4E/RjkGk724XFT3zrxts4Y
87UN4jkWFIYWk8aiHAtl3FPojMNEVw8iQp6aefNl5oZHzu5dRxTJKfLBGMAUGnWAEZ8u28u/ynuq
Au5v/JlxaVIq4dkd5lHk8dBg2CMJsCwKc1VgozPNnOuB/ykEpOpaRLQ2jQVzFNMhoIfEKLS8PKBL
IM0d2f/NlOSj6YRO2m/0NqS3KjaAKjvEMrfzQkhGeFl9d1uWK0czysTni6ELzWpdGx3j6ltclz8N
3OEh21RDeIlw76fZp2f9kdbBKvyDJKqB8hQ14dpbyvl2+Y0yfg4E3/qh0CnaFB7cQFbBleHBUdFt
vRiMNfJ4pKkNgMnW/PqgkrciRjrT1dx1NjCoXrfnWB89Z5CeTL3D9OMK3ZGxAYX7ABat4IZP5zo1
bceuV5QPf/T6hUGFHKnyRWQAIm8MD4EjLgwJhzYfjz/OSYdGXCQb8iEch+Jl7rPhBAj8srdnGqxJ
RrfMkHH104QiTcmZHY5cjgKb8uaNIG+3lzyejaLNsdVHoV8OpMFeNiL2AP0mjlGyax1ikt/5c+Jp
CYHu+kh2k4tfbb9SEz0pw/t7pilIF66DyqH4TVS12zISOfWUmWVzU542WpRR80877YdQI9Oxhrrd
JgWr1KkEAfF559dKtqIoLE2behYGW33NFAw2qVVmzNANKVVwvkpan7XVTt+GyFzaRhvhQagOdQlF
VqisG93ZpUBnTcN+97OVP2UOBOJn11eLNtS+UPehhMnReK1M1ns16XmGAO0+9uf+fUL0MaEtOMYD
zLDP2zpvDkMZFfAJJ3FxTo7TrakhK+wZM5JGwDBoE+/bM8pZxxybC6N4KvaBQCcXuHdQdkez6Qu1
W6QYI2GahR/j+vqrU9cqzbkzZyZNeeO9GTjAo5xPxDNg1hSuImvL40cH9ucDHDMn9RmvakFXzEV7
3UXBRoEa49XMXTheyutpB/IdJ4HMZ2ChWBT3SpM78IAQ3yOmI2IFAcTeWd/beA3jx71pt0EmQ3/m
U7WrDDIb8lYU+PRoWnQmEWWzH66EbQGT+rnLW7NJbZCtCwmRXJa8hPrY09gxFd7Qa9xD8n8fnfpW
ZcHOKgcxpQuRBcZ5ewlbwz2izDvQq637jGoZ/oKii5EhHtqNamJh64oa7Ez0WsFgJG4GfH2iuwm/
Ds7TBMlu5GJ5gcRsoYUAW79zeAG13CwnOxmV9wdMKx8JhFbMtTXNLmMulmcFEU10PzPRc/7VM7tE
y7r42W1E2pEYFTd4VYs6bbHn2beJGrLutxtG/OXkS7ne3ZJk3/asamomSIvoXsKPJlqeXcU+L6X9
6t1QJxSmsBOU6g2mH2ieHN77u4iv1xzGC7H2kN2eMiIuGFWku20Rvpox5yZrhBjij2Cb7h+eExk6
hle/SiS8ojA+MrybUXixhhRdW6+UtzcTYj7etTL/L4qYUCoNKTE5Mb8fIpr40UbwhXhrF9sj9JDY
toiLe7+D3+xkOkCnA0gGC10uajxJotdnfUgOXp5swoVnToxeGY9t3PSEy47Qc3jIyXUWJB8cpVmD
x2stD9ACpho+VaAF9Q4IBwFGl3A/tQD8H95IANVd9AXe0lCF5i/0D0XKJwniwlcYLBaUneumNVuR
1bPtOdQeqhop8nGpMHNZ+XiT/2HZUjvbJgChTV81fwSZioLpxDrbTX0/Rl8/BlwCskKrg6v58E7B
Y1r6GYlwFf3vhAaT0SGPpkIh7v7AO6hwRr1J+NW/VRfp/GcuGwypRdqzHrlzbzIln68eRiM7kcwH
sTuj5Rk8l3/fWd4xcWvUMGPdAaHDpk4sAO7+D/abPJZXiAb17PsAHFOxZ8v1upAXYrtezqOlXk9F
FFmr7WqxKY0da/+vhuffBf0ggLjcWOf9MvUm4TilE+JwXVAeJbEpdb3ZUPNDzwu4vPtcHS35ahoW
xP/Oj0ep3qRbFe5mRDe89X0lj1etmXaVLrcQ2iNghrEU5yHmWTpS8D9h7wGxQiPQgMQM2yYdk4bR
/OC33/FnK77kF4O35ce1SAVhw11t0ZdTZM4ZnVaRJjEX92yLeivAfA2eQ8Zhk96351T0OVruSMsw
DPEXRM8/9jrBXwPBEn/Hx/Z0h1yw9+/BENAabxAUNqeypn2I2GmKYrmubj8CgG0AM7WmIwsJ0tte
wk6cr/hgdtBOnXtqfDVWzbm+Lp5DjlZp3t1CATKaYImJVOreX4Oc4XchZH6BunTeHoEuSIPmN3iW
sjpihDxxokT2E3zaWcTcbxLizopM0rzZAtulSgTW67CEIQ5x3aijkXdSrko2sAQAov0yAnvHGIEG
Y98VBn1/gRmCLM00jEgRAbMA/TuG1/v8o6htFNzseCMOBkhwEPFiPyRrwMzMRP3U7dkX5kZG5mIR
QtU7CmpLI7eSgH10nvxz7oi67+jsyzXjigNk4HYk0oDWGh29oqf+LAmiwMnc4P3Ne/fFw39UEd73
ZnGzFrrIEz2l52tFAWITx6B86RIpJ1HnN7Akmy2LVjHBeXIlUvBl3H4OqwSpm+5oS6Gn8Z+JmU+O
+knC8NrLMAhhhrpfTPZMQcibDkPqdjnon0eypHPfLl7v3pBU5/+TslPo6NKKXs0cKmC5PbwoY62t
+KV2kWk9aPIg+leOQWpFpuZJL+bxUjZTvtBrNv1bNwayGzRh7UJivv02JZeB+7xwIrxunQKnplSc
aiDF0Ct4omL8HOkBpJ09EBnlx5fSFxvSYa1vV/rhYV33Hm/DwhGLYi61UbuBTAlSv140H8qRatM2
CqmLdmJ6yJ9KcQ8RmRz++gJvESe9oRcjS3BuzqjxrjP4gOgT512OdtpvZ1ohUYdn9BEc6vX2E4sl
0VOoZY3ii3+cX1r072eiymEidxRnNEbA2OY2dqPJXhTdcwBW6P4YGYOszyKjnDrdrCk/1VA/88CX
XqIu/ba/06HGFdoV2a52s/5KSwqHiLl8RBiG3MYJG0tHm3x7kp5lIkAfs1IXv67ZmIqC5hoSPpMD
AlNyAQSvsmJ+qEBWuqdfIDDJKi89/HSOieo5E+SG/qau72TwA+Uqethyha9fa71EzlJzgm56Xcnh
svj0S7FoyzMbQvVHUQdFtl6d4hgBi0NKteJxG0lLauWRtxe/rWnj358v1KqB9KfRNv+FxD2lKe2Z
R8PwzeRM25c8uEWlAFz2JZgbivV7JlU46Fp3+1qHW8bj6j8BGzL2OhUgnm9aCnyVlOriBWf2lYOI
QoQs1XvN86a3987jtvXOoLV0NxMh+Nqzu/9dy/Hri9MgMeZeJ1IZrQfShUtiri+7Jmmhhe0MJAuI
9SpS1SxgBD/m174ngQB6nvKsRauXqC4q4V5SG1/wYh6mxAXYFozwEojcD8XTX+nSgogxfc+Olev8
7u9KS7rhVqS1F8rh3K4IeKngDdMinYYOCcpbzGjXd04VhOxBc3yH9ibDylOlPTsfl7u6ie1Qe3xb
im1boIj9Ghhi5XP3jFiWSlEmzMowTSkBp9uAabeILQLEzfAglE0K2tPFB9VQNO4VHwi9hHdMPzx8
6Mb4wgn5ngN5yVhK/QNU2/kSKajzokXEktc7FQg++DhmgucPZl6refrLzhdHA81+xN2oswFQ3PrO
OlzWFFgDxIvo/z/P2nSRH+q+YPxRe5HRPUpnpbAVr0GMEnDZKcA+2ditRbXR0KSJyAQIcVjFyBB3
CSvWuOpx87SRZaM9qWXc17b3cPohlZydFCkY7YIdag+WjHZy1LKu5/XZuM8lBZB5bzca2WJokYHU
Axkv2pDpDyqIm/Em4IWjYyS9zvOwQUvFmF+aKjHP3aNsJi+MVqopx8eDiZakZ+Ux6KIgiEf6uSe+
kiUItvgWFO851zQFjJPvQqT4Vfro+R4r5u3HsfrJDiIDsbsHCP6XGii7p6Ivr+U1PavO5AuQeY7V
P8PuFd5BL2V1esjYJxV+uOybpcjMcTAi/fDgtwzzTHZpUH/zlazsRefK0JLQNza2iWPLyr8nQp5w
BXSPEx1Zeo8Teflejoqu/QvW5uq6KQvCdpzhga+aiZPA+BMtLzScguoxOy1ul7sJtAC+VemRekHJ
RuYoWpoJlpt+CtlPp70F6OkRnwnznPP+92j/8FgwzTmG3el3vdbE0i9H9+cjGKyMGolyRsG0DLjP
6PvI7ZtaAGEHMRNDrsDUdavuaK0U3srwWopq5oCCI0WWtSU+ZaUSWeurjeDqmlxI2YnQJO8oH1P9
k0JF8WBzlGYkuwUeKs+B5MaRE+m6F92Q768feFVcpjqT7S7/LKQwKDiGROdwNcxHRQAABfgUEbQN
BRIHcSsWgcRWTgIj4Ju3j8+3AcQRU9yxFZEivhEoRG3pYR8vXCT2iFeVTHzU8SRzCGVAyUHOio1j
TMaEVRyiKyvMSOjb+gvjah+BxDzubvy7WYaTtVRL2J/WIzthBN8ldPfisQcULRgxZ24DuCweoYYR
zmLy7PLjR0YKc47NPy7yrgRdnmdnm+iXVLpQtxVU/VT+HtYMcGPzpucW5HLiiZbJx9zh7ePeHQva
/L5Opxi5WrfTMUViR9bfcdXbw1+RD5KW/23zuwpPcVi7SqCNdKMD4iENVwOLseuCx+QRTs7hK9SB
BcBwtgeZBvEEMXq0/IxXmHTwS9abtr3IJnk0qzcwC/XU/tQuIdMxbHYjfod6pjlJPi/mu4FphVVo
4lpGx64ixTvFMsJer2Gf9TjtM7uXYeSJ5FcCa1yRfrFWHR5Z9xK9p80/fJIMHjVIcVSYS/i+Y+nw
NNTMquBDjhlWXiA9zXLPiimRVyiinZfRZOQXUZ3kc9T7LNajyLfNItrL/6NWJglJz6u7y9W7Jo1t
PLA2zCQta37tEg64uA0GLDLYToVenZ/W6KI6zq9/axfpTsE+fhk4ooxxCAhc9pfR1yccSzUDofK0
KvTeKLECsn+ZTQ4+veii21vtaPOIeGs/qvOldFrUQ+Ki1dH7UKRCSROyov2cztXy+qPreCL3yXHj
DodoxK5JdFWE2JeV802V0znqwITZHEDWMo1w714pox+LPVxlwPX2TRIwpqRqb4TLUcErDv9MHkLH
gHT7m5valsmMZNVazldpUfe4yM3y5h2N5l+TkHj9SDQwbHS2WX/8ABn7hagXpWLm2ib3bcG/edvX
y8JInD7kzT7hH55VPMTP0nNTEXt2cXX9WkuEJsi4JXDDAEv2omv6eDHube3KzwQjfGk0q1vOGcTH
c1MKSt5FC01gG4jNRmdReuH+VmgCO8JS/FpWHEa94BkMdTszdtj28TskDQjznB9maCAr2HUdZO5q
mFoaCaxcqWx9Oetws+eYKgVYi7CnS84cBc/C4ASZRkXJl7a3OC30NOfmE8ABJ3GRWKQVGnPbFayj
LGaRLhtj6OwChy1FIIptBejSB4a8IKPGrIrrwBRzkpGR3IIcdKRq+PZ1dRqdaxtwvUoyavE/cZcA
GfZvqtT6Y454HH2SC2sVhe4yIWyjlNIhWS/K1nu/V9Wuj+fOuTHOEtMVnVQj8uAaVLhJF/9ch6dm
Jl19aDyJu7mtHiDlyu1JNWEGfJfF9U/l0Om2dWUpSfiha9QlUFnYPEofxJtvxBoLz/qRem+hCwFe
25Ru/ebxGwOleQ97AbWqV6ZQ4XhEWW37v1tACH4p9f5x81KV5mVfABuSR1Oh8gvkctzB0gLdqa+9
YQcwdNCcyLY2h4mKt9dWTyY2ZbXRG5EQPq5zsY3BNjrrXCG1mIAb8prsdFHW7jx+3FapEJH3HXAe
aPyJwDxFL2HMf/DMZnZc2sx7ETE/GWGb9FEsxdv4y0lahEeBMx+zdPsBwoCGSWcF8NxUI7zMIkIs
y0OvbHx5i2vYlQ0YTW6q1Lk4gSqIgfz6fYvFoFaeSQfJ7vuSYgd5QH5qQZFV0dgmbXIevevVOKxo
8h1wFBETaAT5i66ycJkzdsXNaLgws15jcYa/8jiDlKkqAnDw6wtBQvAop4m12iGkN+QlpWrm8Iv9
ugV/uO3SAOEcWtFvlw3TdhdU2shFF0AFcWS5YiSPY4w5o6ylGM2KciV9C71YvqcWvoQObSCkBuGq
tpdYP3iTLmJDmjy6dUG0pjWezsTPB3CqOrJRt9nmyKgN8BaNzpXlITG1kU2EuEbrSx07GE9MCo9c
2jp8uyJT8RtHeYIbkX5Oc9DOigRtkfn9PBQqeaRsSZ2MKMA3hU+F25Bg7fHczzISKRW9YRawzZNv
FjQbP8og35mKLJWG135poAwEGZ4JQSlpCECGV5n8rMSnbJibn5NMx56FMpLt8cmmp2CzD6VcXGQn
ZjjpFUZwwCUkqLbbhevhqZtpBV2RtN4WxYKdUIIBqalALGSNvd23Wzx1V22wy5Hgvooz61jDSKva
LFm2u9I0VU5T6AiJ+0hQcmZYhphrUhLx4qnh1MS2ATNR1CJ3PtbqT79v6S8KGHeLu3B/75mzhFOh
81FGYYDO6TAtv7a2ew5OfCdtAEHWLk2NiUUtYBUf/IWwKtAD3ZVDHvSQ8jjuTebCa8SKAaJUBKBi
NE0vGVZqGkRLP7+5xKV9y91tgAvTAAlHjwNurfW3LMtBxlIF4eYayoa4xeS1VDji8/f5FScDUxFr
KCo6kcxbB5oYyIM7ohClsVOi7gVxs54VGzRRu2hBIqR46q4mIIhoqDcgaEmvBg4JkLi2cMvaA+tr
5emCdKCqiYTjPzv3IFN8tw6qM/2CQNv+R5Xjhkx+NDFjCIYMWRPXgFVYOxyOH2HeDKkWS/36kx8Z
ifpbMuY9XiSsNx3a1p8FZblnPWqPHdJTmVs6bz8t4E2KcBfTl1wDebze9edoBO2OewJPUD2CgM5Q
diR5RY/imSa0n7TEAs6QDkQLFTWgl9HxHjPSmaPYHYRwDqTFzo2LcQZs8qD8oumwzvanqMKXa0CM
hQvxz6eYfDUb/aPEnBUeP7OxyLMrMxvHEP3jk1kbliNVSmnM7OQSaGaGgRHPV9yliVfHhP/4KBnj
Mv5bE3RA+lg6zmdh2F8ZQO6oUYCBhOUpD+r/1rL2LTahSbcQvioNpBwgg+T4nvcbOPzIu6wPkSie
gtlnsD3nixBdB1fBO5/t5YnYRPHxZXtYdSPLY7awikfyz0uLNPk0rrEFLk6wBtROGNhauroWd+VS
W2YUK9D08OD9d9pB4dLrbLp8TOHdrM8WMe5idBkTYT+FdkupWBUl+Eh9vCWTHVwU7FUn0qwt0vyP
RpYkeGVuBtxZ1NoDWcJWTZjP8FIWB3ewjH0d4HlnWEjJrRgcAZHmsLnxQBeqLZ0p4BqL2NoV0ELK
aMpzS8bBpzEijRO/JBhGELApUgQ3wmyQQ94M2iIPCzMHw6CLyuOCZhGiWmlhrp9qI9McWItkVOrk
+8Ywb9kFYBBaahWUxYdaqEWP8EO8pMJi8AdOs+dwa+vN2SrTwVG79KvNkoEQDk/YuvtesALJG1+/
vqVbfNQCF1+hz/ygSA41+vMEMAwiT29BMeZaXm478R9vO4fVo62VdBY/NIlf64au4qHi7M1XkjqA
53N755ZYM9loKwBskLs5mQ+xvCaUfLIhAkRYytU2nZK2THVSCY+cnzvxFdJvlYtDCtjAdKxF6ch7
gyJ94jT7k5CsvKzbLeMtE0wGCPBJqNAvk1WfSyv6uZ+y7JFxeZGXG+wfFmeibORiJW+3snBN16e9
pyyoLcEUhC+DRstouDp5/F/ypipb/yKM49l6HUUrikz+CTelrx/QPe1MLBMu2EDUl8bsZtnjAzq5
JTs95zPe2xd03FkfYEAGqm0xZqRRoly/PGEZlEVRHyKV/Qsz3IMBHmpBGAX28D4yLWvQ42Ki16VS
s8aFJxKmmGyeD8U1yfm67tU16i52/muC9pMbtdrQz7kgfw1inLqH9swZUV5zNuXIa/Nek9VuOhdW
u7uVAxv0eu1KkuA4jdPGiLsREhkUR9aedmb/VqgCTIzc6tMPufzGuYqH1xSQCE/YZthzqb//ERvU
GkZJDXOErcMnp9QtrEBG2DT9V6xJOW6HUb1HnTrF14O/CX/rdzUE+W71vUaICyBJKhpYXE9hfYtY
guMuqXqpy1YdPFlK8ymDxzC5LQRZ1XQHamwdd2C1ILSRNhOaYO3WnxJskxpcxW9BxzGmZtwZQJEk
SMIKIXOsX0yczHBwGRglX6HpCqb1eFJ4TDcW3CK1BhYweo0o01NYAyrvk40ZvYwsEvURs8/KR7oR
Ao5OR9gE6oWeNkTqvE7Jkb+bx6fROkt70Aex5g1p+Cf4kDzZvAT3WKkE5SwFWOhTtjuuoLL1hJde
MnSkgNDVRCLrpN4D2/Hzj2cJYXt5c5Rb/phGoW7pJcBH3iuHJl2BMXE94dbCDMh50dIpKbSVJ7ex
bJ20ggsTrfD2MR2gOK/1qtK/kZRYf7T2l3kRmwxzCLQABkXnjgHvLL8JNwFiEt7976Q8lxMEQuCz
onwQmBajBqSQaJrRrAYwNIjy9YwMQMX4hwJigsNpgvUQdkgLvimTNfHtmxegD6SS6UTQmLxarOCc
lSC/DHSQ4rDm6BZW/iiZ2xlrFyM8PPK800QT2jK4u2OPW6Ovn9Cfkon6U5xblw3a+XE7KCCsXnI2
jTYFsz8L2IyIg8jyW4ghmwzZuquE0amxhbGe84s3m4yeCqxN5Uon6bsUir0uCvmSVzna1J/OPy+W
ZSaRveAnbKvr2jFm5ncKtOlMHhW0sGdeJe8e6cc2dGLy0BOJoG1S+Il/SFggTWz+qVUpNE7PUUAC
I2XxzzWEdT7IiGZS+GpB3hetPAwwxFpmE+7A6ZDa5w91qoqsbc9B9u4zgmRleCfNwPozUZDer0+O
/xH8f7YMwkugMVBYRsECJLzKbf8lNuhNQ2p4/9MeDhnKz3QmyC02oyHxChFLS7wgcblOphgke4xE
XIxfISN31xmyMo4pekG6FqKUJBFeq/IqJkFzfHTvgnkOuytqzB5i71AGABCw1BMpuONh10ZnMC+J
WbP7c6tLw7pbmqWn2c+jZ51HXLqTW0O6ktEW82PeLjiEmcWb8QZB5KRRZl+g/gAYSMXNkZ4+L1nL
isOrWlDg7LrOmzGMMi8CbB2oB1p8l/TS7lXuOojl81L7JJpdGuUR/KMOdo0teZK6mVE24Y6FZkTX
12nrd3mo6EvijJBcZrRDrSj+8UD9vyCp2F/QaUwZpJmTzC99anPL7KSfRlg+1DqV/ggDnK3uOP5V
dXQ0rWGBqXA83uluF7YQKR8vh3FvxAvzHHPFXfaMAbgVEQ5N41wODe7Dsvd+T9wxHbKofvNaJk5m
ZYMAzvGgmZu1K8OrdZwqqmbVs4rsgtE8kgLE3vHSSKJ0hocc4uN94f7GwygFw2PTVBuKhtfeT07g
guwnRIC4TCFKnVTpzT42h7Py9y3y7/cKgHkdjFj0Qh85nMmxJDSaQDRfu8fD0Hkf7Rd3e/C+c2rL
OFHH3D8mwzVi/vooQi9pem8TuxNLXPexUeYyXElyvWokRMF9hXyBrzwTmbd9WR7/zdnv1Z+HrpVj
TA8pRCxb9+A9TdrdWD67XpMAakGi+fCCp4IXm2RbMUg9iGiMOwnuSfhrQm43C30Zc25LCJ9czU4F
Yth0ounbOYnHByX7gVsj2CGW1Aouzgr/ddl5MnB7CusKQY3DixWoU3Ws7grDbmBc2Q/2BiE8Z3yZ
slaOr1TEKziFetLdTRnx57XzitNRwziydPX1+ajoymjMkQ7IlDcBzyMnpy3/yzNxgWW5x8Pdq0rX
zDy27bu/fGF5HTc+1r1/2r2nz4IGu8xe0Q5rVkNA7ZLGTcmJd9VK08Tle7f7Qq0ptCneGjy/tyT8
kQwPqgpbXS5Nsgv3LYJck7G9b7Ew3e1S0o29L1ke5MbwUfrxqCIXbpXrh0oZos2V+hM1irwXg6zz
23cH/s75Om/557fPNjpUBMulvNTz4U+6iRoUN3lST1eM7gpfOFcKLL0xpt5+KX+uIAqGri7H3cvF
vTiDUPA2rsFj+kQ2g3wT9HUyfnVKcGbFa8Lc52pq8CywWj1MNhwojQciU6bOjVI0okUTjKKwLNCy
ZQaH5wzZ2166d0cno5pc6fsUJDUzRbVwycyPgldadwJRoXi78QxYQyRaASjkgEmjiyrZXkzxsPmo
KXsMdUunk0bwEgegUYuBVbeS8x+Bh57Z2X0E6miBGLIxnl8OovQYOSTzazN30HMbiQWl5Tg6z/xO
3kasW3sM6JBUy9CqtcFqv6uxFZBO1LEjN3VQ/blBi4bWQgD6bY5n4mZwX3zjDngx8KKxd5QOnXVs
g3TFx4pFDxGVkmtkJdISv2QkWmV7cn/hoqlIn/zSfgL2BJd9kUA/ykFOa9NiN1U6r5mNq45II4Pl
pvKvbiAvfgC87PO1n8S7i/vvKhA585Nx8YqRf9hbtEnT98EKHm2kuqHQxmBh2Hjxa3/zexucdU74
yucZeuEPe5GwFWnphBDpr5+vHqLRW8vdJ8BbT8bcvQ6SyFo3y3rzARi9asi3XQMHl4SXonhihRbJ
ETu3n/ZsEQfXBZgwgcEcfXLy5x64POrWwAsxanRZUQcCZAwK1jJcKORNIsw0p5KLUx/FQNEjCBoU
WWaIckscwcZCSoCglWTqc8/rCg36AZ5oQQC2AbDRhbtd3J8K3OcaAwVCs+LwZWIIYR70F7whWeHi
CZnoFgWoNnTa1p+ejP442hqV8tOl5ydxUDSOdySu6N7GO+tsNUfzFKPxJyOQsVRUgQoVmqgu7AKX
R69U2gmkuHjB1MpDdI1I9WrPFTMVXlEZN724fSINqhsQpQ6/9WtfXEO55nBxVYs4YZp+TnuXIdQh
sg6BgNSImabSNEjtIjwBWTFUVRuBNThQy53k/iJVq+8HOcWWzyAhu0UM7ylm4n0GWicfaJ3PPgCh
lij4XKlTvVSOLdj/qm7NgFJz7JKkO1fgisv4ZMCcavbQgJ7420+EQdtyIvjTAKnpl/zpAUqYfhbS
3tlnzX5GwKKXVJheJ2Kgyis7rnyitY1UcBrYPuxeq7gJhFCeFfvEdvqStmF8Gy4XZRRJHz0yeb50
A5Pt1g4Mq1NAaqaAK7tOV47vh+MtP4fZwPZuMO9jsc90Dm0LCuVUkuBNDrv9pysZ6qPrK6YEsmJp
5Pf/fy3qOkdkDdWnmXSAldFfz47YCb9h+sh7+/rCSDOhzBK/aihqTQp/nBMNmbsLbugkct3ODh6s
MAqME+3l05x6UZ941/vvq+7YrLRVnSYaK0UKTfIuEv83TriSGcHcXazJYHWBk1X6ZjEOW+cEiVhK
WWcexS8sLtOV/wodyTu2RsMgOjGEB+VJZFy8Tp8jitwoRJuaiBMDdrBtR3YN0m6GLErdIBR7EYQP
Z8JEI+eyrcNZ5ceJSr7u3np2dIjXqet5xYIryabQMms9xYOIaudvx/mKZF4p0I36aEprwkHeNf96
mb276ZrtCkKsa6FMozK//8nkWFUfoOL+yBakWGgGx67Oc4aBLdXRYUms5zkSAw+Nwjgjvv/OeeZM
iNArQc4/jzKAhAjf0qTR3O8JFOrbsQa+BBizQEXnW+2DpHjRztYU/OOf7svrSikhWUEVip0bQrtn
aTZyW6xbmEgodRr9pJ7Pb0GHwTNtadKXjbcaPwrJ81qr1iDg3vGfYumluK8xlA1VxWOjFcJbLMnT
YOlU8p1DPg1Sd6X+AZPoL2e0zcTkw9wZktTj+Lb9sfwWnJeU+KTJDcfD6E45z5uYOZSPUO0pqXn3
9MiNylWxcTft4JkPRv0sFqNMf4KmRCjdKGF+Vo92FOI1iIObjxmUyFBxr6Aks7885wyxJ5FZSbuf
9OTR9Bfv6tMMyKToW7bsk89UU7i3Zt2E92+qLCn021nr0H97ldNyNd1sV6mLXrr/xi3RFgNUizDf
CaBJs0X+EmSw1hCtpcQOrQAzapQ2125nKIcAJXHZFMNdq7V3RFQSpvShAwh4liqDOfF3MQ/vq+Lx
aEj5AiyWd4FBHRefkrb/hZOyQhM9WS9igNhUZf9xf/saDwoSfVc4atZJt920VETvG/UXGQicj+fO
nT7gbdZHWcDHTVPIVWEUXXw6D1eoiXjAHTW516rCaI0SSXCu9sbCuG8sGGtr9h0DFu6r+nEg9gf1
/ehzhdtulldpGwea7e55/IWoiaKxXeDaaZx8rKgODYmhQa5PGgjMTbAvh4oudlM/jgaSepDhBCeO
FqWCpiPDX73AxghVs4NUVZxousv2tdQBB5p5IfDX2Y5wI34hMBDyFxMAxV1RHBG3E3eVmgkIASxv
t2VqnrsEmjnzrsgxVOfFQNMaN9z6tpwyA/VsziI/oaBDAookfLJrO3nNX+9GxQDvuGQIPOQEXrAl
sv6x2UR+Rb1FBl9uKtBqOAlt5prcgdv1/zwmqiDK217CyTsaqzuMjubuhPmNxcZk7IJxaw9gsPwS
fVvfgRFXMPymQWGc1IF3Sfe8CCY+l+al5ctEtPD9sX9bwFrGJ2Za7glSPjuv13raPvwva0i8sUy9
3tMAMPIiR5tq8sqy6AsDIQICSdhdIcnoPpYzBzmekWqj5Em2ZEmLd2JnOMnLZFFDddWjhr2URTF7
luFC968iNh5UA8O5GBy3rMF04LveM+CWr/2j4s93E/D83TRlbS1mPDfC76GAdwYnFh9IaiqOk8MV
jJeQdaDw2OJhnYyt+Kfm7ChrNsTdhVWZOEizpIrR06APZM4wEftuDJiIujbePWB+TcmPrNZ/UjLU
SyVnf59ZIGOKtY8ZuL8arGgJ8oyvjuYCChGYnnHI9RHku+QoiSh7aAE4Lf+64NXlQIOTCNaDmbN3
E3Yaofkx8R37LmvonJvyhVzisn4HFXHenmTyUciOH8VFw0jezfHP9SbKkZNqV1q1b06ZLE5St/Ir
fhtdygupBx82RXrpb3zJM3cZKxvldpdJ0ZDnw2qHP6v4yp81mKLS9rNqioQJpTWsoWsgDey6MMkd
E0MUF3i9NH1TMDOQjQDy42Bqnf0p7L4oRP7Tp/XwsZJYBBwqS2j6isIVfAZbIJSP+cuSmEk4W0rK
ct0TmXSIJAyWmvOO/ACPBJwxmLD+fqEJ4WddH5YHlC89/yNfETTVaOMb4KH/aAf3RbFeCIkop87o
vqR/q3mbIPf1HulVl5sNXDjtodA/xt4SpDykApPNuaBWSfqGxQNwoln1DqGsXLBzowst11PCIomH
mdefqxCtbyiJB2S7k/LFLdTpZRRxkBP1zwYhHi7s+/MkvamAWvG2+vFx3izSHi+n4MCJH4EYaC5V
0P9fK6ELTdsKagIcz1x3bLeISDdYBla2dPLqrJ4y/SyrMCVuREui78DiY43J4KV6+qMC/6mz4Oq5
tWakvtVZ4FYVylZ3DPYH9YiAfbr9mRxPgtWks+uMX1S+P7ojL4YJNyb36nHd/TeqYtrQmrkQ0tQD
JiFcVsN8wsrNnrChE1OXRL81DWUUYklJXaTz6b1jZF2TviaYdD32XM/KyGjSEqotFspaNCm1whyd
a3W0Z8t8T3MwKM8ZvLW09PnWTiKxDtaxpFdyQlZFvwQQzOGQ2GQ/Yq6YMjnnf3TkaCWnld/mZcEj
uWidTPZ2QK4BFhYdx/WoRRLuYtH/GFnD3s3OjYHazIJx9BPq0mEPk9xXf/XEYz7ERaFSWNJyBzjQ
SgoCg/fy6HroX59Euv4iXfDhaOr+TcYzSoOGGFL17hdTrSkBLzxQieIYnagiD0Y9XDS/ksIaUcex
Dy28NJO8tFoUYHZLjJL1C9uuXW7vPZ1j4COhph6pl/DyZARDoJRRFvXyi/LyP1hUenqk/8PvgPoZ
pGw0eEauNw4NRF/RdlQrgdgAA30mBNTwOQrChTOH9765ogpn81UFQloBqJK0a51kGZtzDrPA9pG/
kXvVR+xGGfPtjQuw+yZADNeNWhEvtAsTbzwFKc0DoU9KKK8kwfxomhF2NujSa5g3Y92+xxDz8tMV
3LYLBjETRa9dnAcZnu2uuMlkyPCE5ElLrXvhyHQbzJMX/yk4d44ZYwQ2EN1KaRDGbLf1zpiZtUcX
RorvFkkkkaOvLJx4FzWJwpqOgo8cywMWIzlJrR2rlGolzRWtaQAzmFX9kysBMTuwOPIJ0TZhuP11
h077WF+jZNibsZ6YgUOeWt9AijL9gzAM3y22UVKE3FKMJF+cwbQP+78FCtv502RG/ONO87eZTUI9
v/iv53gskttbXMadB77fkVH6ALlVISv8/B2ZWk5fw3qbaCUZXpHm16RDbeiqvdMX3wwLDTeXQiZJ
5T8qVWCpLgZ8dJkDyNDujVAd8ZO7l/K4u9fCZZDjgnUlzt/HOduCv/eyZCxJiiLHg7C7lVEzXNN0
B8YrUIjXiJ4lP6Yf6XUsVejnLayGzf8kxOv41ZDMNmQv2qh7VSZuIpHA27IOgMJnraQc4n/qsUCj
MiTVtcso38u0A2GAew2YItsS1/YZ8gW66MzE8CAXqKD5fBshcpPkqJUDcblineoxZHvYjpsTG+dc
YgNH69xjMQJ3b+qQxYy/3fMHLODCleG/EFOAga+vuqwqL66IBJTEFLjR0KkeGce1qreTK7a5jE3p
W3j53KeWqkTp9qm68LkvZYxjFp0arPX1Hk3b7b14swfU+pG6Y+yyvD/Yr/EK+Kv3YYMQgmHSfT8J
zO1exQWcepCit0YNyF4t4EmqhGZJ3JBNk/QitejTA/DIvMSOePd9+O/WOw6WQSLa7jrdxMqP0u/l
kPJkgU1ZZKOVtUBREGSN2GpgL9+wv0l3qk6h0VubBnHgd6C/gLUrbiY9A5ZiLmvDcdRANk7K2Alm
h5xP8rPnxAbxHeuKM7RI2h76cf6qT0T2nmQ4oGdrwcPxZGkvZ832210W18xL5ZM3O9FwMsg278lr
K2odxhkTFtWSYa7lg0k3aij/NzbjGqS5QEFlH/oizw4BvxL4HrxSi2jmOyJhG8lJ24HQu+Me+89Y
FMHSr02h2Eu5wDKSFXQ0LI7jKN1UaoJi0bJv2BMvmc/rQaOsIEBo1dUGd5DfDam8ArmOHUCqCwrK
PpTSvOcQqlqDg3bGNb4vF/cItKKN8FAGGsnLTjz7ipUmlFXfegQnJ77icXFw2ypluV2jWcNL8Jxf
QdpopT/bx8vdWg1C2CQgvAqfJCj1i0XmM73NRDkiyoA3Od6eNp4uhDMMI5NMZMjfp38RNWpbuQJj
j+zdksuXUH4CQHhR7Ol0hTpaY4X8vfIHLzNiL6AurjEurqOv90Vh1CYmBgk5SbiivfvkHU77E43o
Oq6nPIrMeJHnAmsx02E3Tia7GyEMMPNLwOSTtYGGVqIUquY4hLD6PyCqvr7alvsQoQ2hq8BbKobL
WaJ2i6O5x1VUWfDl3ldAk/2knwCzItKn7fhB2ZaPDRurj6je2rZ8OxAOz0ZK2ggW2S09H/Wri/6b
toxB588DGwXi2WXTbFC3XqzUsn2+xpk68DYw/Olxhc0z/wkI2YyIX1YwPrk977hIFgjPCzbCISHG
Z/ffoJX6Y9Byzv4qqpqqzlcvOHPmDVOHMDI0AB7rZqX+wponTRZDQZoYKau6LgqsSMCl5WUijvRx
UpJEwjTksMIQkJ5E1j0AY1Ri9X9Pk5FgG9NvsqWZOXxWrp5dA4iHNnov55n26IXb245kMBdBE/wn
lhImhcs0z86WGiKHocb28aeiOyiATKUWusI25YEMvnKmuN1rx5yrAu+HeVtNHqKsEIYo2yL1FWtB
oKeDw7qGwhY0kNkbJixzmaSiD3nZCmmZbQdQ2avjnmAhdtF0LVFfpoqPokag0oUpY3j2MFyaQFsl
66EGY80AKopD42dlcXBpaCm9wxDRcjHJlzNlmM33/tzextHGyypeWIsv1GLybRFyFzU3ddBSJmYO
tce+JSZpo01CCNavhr6RmxKZdpJy4384Gox3R2pAvXCkC/dkzmngrR6T20iqDC7JAKf9h6HagDcW
tVv2jCMhh2/1jn3kqacEHxikYU3GPNWOI/lXrfNsL3l82f+qB6to/f26YwRMBYrVUO3DQqlWPfMa
+Bd1J36kqKg2AdLRDiDyFasKVBJsqizba6ZNB9zOZZHxGp8s8fYCgDVgjbKd0+HyXN2/xqHS8eS8
77CFiWp3LbH25etjnKHF708FYqGCTSMm+PZUm8VypgvYWbsUU6j4+MM+iSwPVhZZQuH3UmZIRXd6
7lxVOedF6Iubxyrsao6DPLhkszeKf6jE6YGVHyM2citEZakB849tumWewd6V69C9OM0T9pvlnX5C
jkvXWbpwLDQx3KSx84wjQnly5QERx7WJN8x6o7Lr/PZbGarAsbVpK37dcU/MNc7f78bu3dUvHBDO
JZ77M64JpxxCv7YtWiGWAVrvJQbsZ/1WbtcxPXtrFjKcXUtEcHA6MenTWLDNu02HD0O4GvQ9WIfZ
JNf/6kpVxA2D6W6W7t9FEAAn5Pb4F204QL7RoT0xCFUADQJVPzRta5bq2TDKI8Mg9oaAW0Z1u7Ba
KvDusQR8kjHZfGud/FTK8qa2dXkcAqmGwZie1y4E/9vT5nrPzFS/JtUdbTZHtc99onTO+FWD2OTZ
wkY3WLze7VgVTOqLfEZ1o47QWp8mmXkoIZXFmfMcLM6E1WPCjpxg9uQKzjApLTIKP1gcyPb9LaZm
O6LsCoEuc+3sv/fe7GZdV6cXQ+PejURC9+e6yxi0PzhtELRqyQgPysUBG3XfjM4RHgXvk8HHxMfw
SHj4aOXhXGEnFB/X+xkAdV5pCEMqX5XjRT7iiGtLa2kp7QgDLG8AMCx67gcSrv9VLDQhCjdSm/rI
e/qP01x+ZqjqfgFb2lxMmNrAX6c/nuLVD+ejOTt6ok8weh7+Njb6xfpCfgvqANkckUvsd9Ufe8q8
GRI33c9Aqq8zVC+5ihnppLNvkzmHWw+q1fFfZtc2iLSVGa71PcH4Zr1mTBJMUaZeh1T8bXjQDzqy
t02ff504OSP9Ezk9YuJOkt3VbsUT76iLo05akzOdDQ/RsQjXzNvyr/wQ4/wqsz3bScUfGhrMHObW
Dx1IR4VCmXm8FSCuRTdzbbfP5hGRjR4V6MwbT0iT3OpO0nuliRv26wJy8D3kWch1PzhlBPJ5hS1n
+Ffw3Ul4G1IIaDh3W0oG+Uvn2dVUF//rSFEoNg/UMjvlG2enlVfkDzgICGGriGspkp9dZqW9lg2c
hnhi6d4B3VcAdk1CssAToepjn7dc/PM9RztV3p4M/BshjF61+VeY/wBVv6a+g+Rxn4hPrCNUH3mi
dN9xy+3VCfYdy+LXc2u6DP/+vZvXaV1lwemSwlyXgPZ8bJTvqtDA/Wsi2+8WUreKsjVRrcq7JZ81
5uAiWzeNWb18AnyRxxM7Z+BFPGkeuufdojTharUk1A8bYRvqd0w2pPQ6+LXI+58Ryu4x9MMhZ5+3
KV8lv98YHbKk4TrmApatCj8ddI+JV8JPv5fOppZ9x+YVEtKkpgmlGsSriCka49DlCo2VRh3xcw6V
BMdMBeyR++syXUUzrME/krUbTXMJkYw3Hjfm3PTl0tFDqh/yiD591bplSo/tij4eCWaI6c/t0PVD
c2db5xl7xmrxB7+W8dm0EaQN+1C2YBP13adCC9MghFtmYphFvErJA8KLgtz+HaoOkhbVBk5dSanI
F9mopU90szXgZvFEtlu/0bbxOcRu/laLAptQaz0cn2tqrri8VSBh5ev80GEXhl0RePmAth01ma3Y
A6XI2Yf8GlR0yj9j+XDVIRHUYr4pN9xSehTYanHFBd/CCzIPjq3FhnDcURyQvcW3VcjG07t5m230
gNXx1TvTkIGdvtIvxaUVMykNDQgzkqL9B735ljYyKfLNKrS/7RXgIL3m4BPdUFxx+V+Dz1lz5m7s
aJIu8NcDubs1LVMRfbnWWEMYaxq9ZPvGPOdW1Tg+xg0EOAdOs/S9KdFKl9iUDtuVCnXqGlimwqdT
D+StNL1DLrmMDWvV7CjbgmO5GMep6n0vkLHTXot2UrvDcvmOPnV7MskVYhuGYOdUFbF6CcPXUs8O
HI4z1e5iw+Lf+Xr/iecq854r2f/EPt8xfdjsMjthMF6n1fTV1N9SoPM3iHXuHI6R2K99bj/cOw3a
rPCyV4l26bbZurA+9lG9L2U+QqCoWJRnWeYnJyBub6AerXHhNwqKq4DUvdn5UdjUlS7YfAPMS/Kj
wA+nc70rjwiBnhAP+AIQfklBvST0LCg0NHMZD3b1GUxTfec8BgWLVL22/UnuMzmz29nExPanTxWb
xKDFFe/s8laabzxqS3PQSif4Y2UhJfPpXmjS0bJt3Sps9nM0767dG9xjRN/7SKkaHuftJA+ek2X6
rCDuIaHLeUy/FfUw+9a43Q7kvmwAL6Oa1wWOdVz3QQPgcglNihj8PBtszjw9+q4+kLJP1b+HfvFl
cPpVZiGX+83RXNfe6rr9cLDgVCno55fixjSA3jSmTsOMzndxrm2NwoX3r8IykODSy1SrZrEkfFxT
7LnIeoazDEoFjzUPNgHxa+J2F26hKhDKgTl48U35WAwCed5yNXYtSA5oBAMlxuW94pIxhO97uxT0
YAJOKok9Owhfrx4jr/M3q6bzUW23kuqNapt5R5R8xL8AUIPUxXMYvJ2mfAoxwHMDE5W3X0Tsp3cl
PrwyQ0hkh4ZlTrnP7/xQr9SxKDlFkWzHnALC3S6/ntaBapC5XNpjY3Yefaaq3edjOwYCStQEynu2
uVFAYCBLcgOCqGKmBuLhSeMhdvMqcry/rJ7K8qSndIqnNZRCLK+fzceq3Q0IkD1z+NkuSuzo0Y81
rLOx0+Jo8qUDN155ehnySo2rWbI7o1d+RASa92hNZoQZcUQIuvjrrbSYhgSgI2qvqzHxgIBRzJCV
AgBRdyHpTFbfQmxIelznstUBD2cuPfAMPhIiWm5eBXelmRCn2TIhGWcEEQghiCGZdHVZ7vmyonJg
rnZU1+360rpfiguhT1z5l+zF5IwVAk2OEuURVOyVirxPBsIUE92oPJFQTCqpzPDyFnRauc9eubK8
48lxd49Vp3Vgbs0ifZf0JsaDmIPwZgc949BA1oCmBwTmwoV1Z22pREehyUDkExTDnR9HHbzBlrrc
dZHeuWl1TgSuHJ6/BDWipYf800o5MESg+tsPMtYpJbsH4oJxrEnI9YClC8377VkUUXch8Jn4V/Tc
pSSjWKAN7v8Jm+cdS9bBR6eyFK/ZXygO74W7CGKHJUnIqi5F6zEt8iRCePE3LoHulFBLy/pNu/HF
MaGxuGK8oPqqqmdvoIV45FVfN8qCNYdFFFZa4ocSN3ezESn/+v+c2n03c58+8UtmWSm1X4z2K/++
b2W+K0o33ZsunCXWvLvMparhjCE38JhiEn9ET68ehyqZKMF53ZzVaXJigNj4VNhl73Na4RF/m3f0
38X5id1ep1jFCN4fO/wYJJEy9NIKxGm1SZPk4jb+nWd4ixp8/YklVIYzzzeVFbCmbclDI3u2DRH0
q046vkzcCTb4l0KjyMwHQrOpvu3JfMeW7dOHaUyqbGfFh6V2i8te4uvRuCVV9yygLIttbpdV6ZoO
HcMsoq+7AKt5BS3lYD/ifxMqmH0qf4wtrxD46KeWYM+LFbkjqyWiDV0zAMtEz14YBXQiKBU0fTlS
/qR+hGkVVvb90Yv7vMSCcOl4OZxWMhvAKjCpsGzgyfzt9yUyYEJwWiOZcTYFSBl3BBpqd8o8cToS
vBwnDWpM40kSTcV5iUwKi3sf2jcTO/p5VAFI1zeTre+5cgwVH3bpM76LFkvlNsNju29d9yEYRWuW
nlq1t9/ef8oLNHNy4Fg+5l6iB5lhJ4Qwkhi3yveBWuWg7xpjhUPQgwGMOEP8BU3/C5eS/mtEoHrA
2FOT70jVi7LzedGkeqx883hdhq3FV5zaD/e/L7KkMLoReuK94sQwlOwfoWlRjlq022Xup6PV9q84
Mnet0f89bbynH9pErcfvzWvqz4DJVbqOMn+4J5asnU/2fDwSDtprUu79CnRJwf+O74TWFy1f8kw3
gyQyl+BvgRYQsL/uHFI4iRpn3EkwML839O5y10klafHBx1GyWjQz0ZNTeuD4vkzv3qwS+ltnIRFR
1ksPjpndNzs8osocaY1bsEiPLBQHA2oivkq7nOqv6KXFYia00VrkjL4+X+JkmZGplJ4W9tSkeDmp
ECvf0k47uPQma+1SHPCzryG3JX+kikikUHdKWOrOCgVmKrkKCkc0VW6oaPZRUIjka6u8LsULNQUc
m7y8soKyQLtHBO5ZTOCCMaZCfDECOiI07sDo5VvYhINgfTMsdf9sqZ4p74dN3hrVxmnp8nt7u3kI
LnVhk4S+yHxMvehfCPcWAylxm3DxPOvjnQeC0Tv7xsNm0A3ei+Ft0r7yIQ/qnHnvIg/G1YbzFTmB
EP5Tngeb1O2NnplU+evpJwO5aup6aKROLGbGqLK9wTL+C4MEnFp5JwzS6KxMkX3WB2SHnQy0XosL
gY5+qJawQIBN08zORcArKT4xA35T5jGmvdDESLfzIj/e3dl2gLLroa3+uFVXFW0yN3fXxe7Pnh5h
a1mN0GLjxiGaYbB4DeAjMS8OiwX2JFaXvz8Xn6HBYfUXoYNSm0mj5DCCtiBY8kK7RIsczhWTTHCu
pg1XgFuM8Me+ezzNKeKHowJbqD81f6DRM+x6vQJPGi9GQDgrA1Ki9WPBuCUNzMMeXGKHyZrOYYwW
8DBreHBakd+b3atNiu/ncXya9ItdgmEvWinu/N4wIQI7rprHw2ceIw92QUGxO5D1/GOT4qUg5Sz5
7jfJt5nOHM8lmNAB0fNHSV3gh5xHdzk1Nq3XPv3fn2wGZ2c6awMXtDG0AbiPuHX2RfCb9vNdc+ji
fEFwolNX1FiI+tHkr3swN6cxXplRH7UBg/Pt5xXg+el8Gf0WrmZ4Xxb3aIkQjtG2lL2s48yiwx9H
zGYZlCh+0vUGvYUG1kY0k4qckf+yf4DdAnsqpwtboap+92F1oHaif3vTui4fFK7idErTyGTy6uJv
Wkzcp/G7nMvOphtRkeyhtWJggIBYLqZRAqOT+K1ZeqhX4Fr8/ZPlNjX+KJRp+RdADy25hwyY2NNp
h5PPJrDJE70BnzmE+RXzUFkPEdBaAkRTwl3LaHMjSXOuPLBpQPYdi13Qas/1XMa0Cy6mR8frqvia
IxmML5LxgdzNQcy48Oqtp4jbcFDyOxMfvAlIxk+WpFuCy12ztApjLisC+bTfgG7vn7gFVIonmj6V
/yL7q8eOJTuXxnrJrbKXYsPJNkU7naQOndAsodlb5Ude9CTG6NIJfNkB/dPikIeMQmGhqxV2P5RB
NWAYqe0Bb6PXuWdtbnXNZW4i/vXjNr2EfN7yHjhTebWEC99MeA7kjqPDod2AX/zsIzIoO6npkiFK
Hr5TAPysgPN5BWvs63LG5g9a9/Qe+aQ9oupEUSDDpMb9GL+/kw2RFAHDCwM8MlQQnoJhy/L3CaTq
esP+JahobpXLX6vp0EJUNpTCEQuaaGbkuwEpl+qJW1HDG7wTDVdH9fZwGss6l4vB9Wz/UxwPndRm
B13VdDRrxuc4EMyZSUcU7IammSQw1w7UTNC6EzcMjptqUfF3C1Vloy6Zz1mW/vmFcoEk1yFV+XM0
aameVukdg/ynTtJOE4WiPxaD6dI8XMJz2U4QIu4WIh1DYXj7VoQkwwj22a/dUGHEzZFa7hmLKsii
ttTCPj9Cui2MFjSIu9X0Oqoixqm0VEVQmxmDEZit9128rKSOpv4hNYCxllNsZXEQqcG85inaoBMl
2k8xeU7O6fDiFeomM5SalsEy0ZOAeEkX1Dn7eH6mqAUvIQZuR9ZqhkYFsU9AuiqTwqFGGvfZl/ec
nis1Mnhg/kWdsWUvhd+r+injnRozqhrsGIdNsqSn04Uh1+gPGFFQ3PYhLHPqoYpyeb+6Tn2trPN2
ZJToF+lVRA3oYnrV3oT+AXM846zBiigWWNkbj6hcCZZ1lsN3PV11Sek1g9nK034UWtS+qe2UNLI2
i+/4lrHEmq+sweEsRLgWfJSrbPMDcgboYSHM226xaIw61yl4VjpcNCULMerB3XikSxa9tjpZLy9s
ZWh2XFSSXyPPW6apcNLG+gXwk2hG01vcusm2ZArbnz7vNKPv8UVtZg6lvLCe1isCAqb17I/K9o3D
CuBjnb+FCev8BWxzMVdfetqg2Dv7Eb12+AF+Qp5QsUl5e6kpImq40w8wSugSQoXU0BrmDswwGPq0
og4mE6FQGkngAcDo6xgadlMPo56ctYihyj6u9iEtaw5m4IOlUbBoI5x6FtdF2y0j//XqDYFkplqC
/rQstaSFIVSwWn8GKn/ahDiF3yTfsFc6PHlNySuvHuI6pCkRbRkEbKcOQyuK089fXIEOha8DTLN2
mwZ6uyhN1ZeZ+t6TtHhZbuVi+cRX2rfLZGxqh0ravkqXz/2inyJzuUr57Er2I0VXhqvT2C/FQRfl
jrgrkI4tn99mV6vPG0jigFDmr6Nb0T6qkMAiVFY4fGJWHLTMp80R/SpD2ula9/MK+akUz9PP0w3R
82plRy4KXuvypatBLaxssS82MKGXWw3Dfh+XKs+4ZdcQl1rIgpGB0kGbnYvQTgUw9YXMRzXwG+3o
s7KkRN7oBgRd9BDYiDqlISwzaylyJHUyUIEQQ+4AnFFaKDoCeT7BPpHi3robW4j3CJ1EB9ZqYbZe
M9uemJnJOH40XJbk2RdoTp4EPXWHWgq8sGIy9ulH2QFgYPav9oZZt562W1AKF+vQHn7NR3j0tBnE
Yc/ySjwFbIkr/daVjJhz62iDruKrWqcF1+cR4ADfqEHWVFQr1z8qS/F0+LeYt8uo4/dP5icmAtar
eyJQ/Ck6xIASf4F/TrQi4eXz2ZmF9V0guJ1bzH+s8KZaW8dcapDhR2SQgiGbPi1MIJavdXdbi1IH
giBFIRknFqd/Rh52csnrB0GJnsJ2G9R8ZSSvMVJ/czIx3r8fdEAYW/BlwhVDsUSVgQQN6xFn82QI
XYMAXN3j1xqH6aBzUet+hpGadFdfK2uMjScMXmviUPfO1sF0b+msumo7QiGV0A77R9QiD4muARwZ
qnmK3AD4Q2K9u8HwvWQCIJQNuQAgEFzJiRbV5fR9YAN/SBbvwDRjFyWu28Fg33HtE6dBJEFtlEMb
rNkIdOoENaKUoE7NlxmIxSRYI77z5GMTGqykFTjIkcYziKsYyDmGebVKGmKNYZPnNTfSK5GRF+J/
C1JBsaXh2vcYV4EV1lXaGMJne0zxfAWI69B3ircECYlw4vskWBUNGI1kyZYWQ72ZoToshf2m1LIw
SKAWfq6vL44ZWer343T5IZP5vbzfGLli1dWe2Orj1vDo7ISDQhhPz5H+ztnB7U8AHTVjjdrACaOa
p0vDhbJE81Ny8X1Rg/m7dATr5VqEuIE+XHClV4eEHuLxN/DLJq0w2Y7SPvWpg255Fj6T9mm/Q7VQ
hafDtiIjcTWdxVeq93/qUSpyECNmSotS4WzXyiurd6CLvtu6wT7a7JP0RIV+fZ/WY8W2rc5VpVqy
7rEKtyZ2HD3DmWCymtsdHbuYFFcKJxiTtK4Fsz4EwPsEaBr9kY0uPXbIXO0Swr6M/re00mmQq0tH
wh62x78V2bBFQvQJOP0J29ss08Lr5F1hK2+IYKwyCXs+e7ziCwriZvsF2CburIBQvu7snEmQ2M+D
gJvHmU1pdrXtGVMLe8+pjZSPF8fbTLubTVhTvHh4FJi2PtdHvU9+bvILGelB5tWKBFJzW/g7sOJV
mnh7zs6JO7sArwgFlbSOIByr5jQn/iSIcx6WGMK8bbD25NYma/ej8t5HNg+yywcgE2x/wj68ihzB
g0J3BjJ6oU6H6wur3VbjQjKdr8iHEg6NejYzM9v9sTHO5TZvI0t1mQPg8pwbztjKQ+aOgMKipiIy
wKGL+8vq4qdVZXGhHGErWJryGTHKLmL1It0ltnenXH9gYWpRdihdEPx8IGXm07KacHa9w0nh3DQV
rS9vyD2/5KoLjSYtwnpfNsCoitjS+DZ2IHMpdUkNwbi4rukMiweaGQpi+SDtdt3tl5LeEkRxN82t
yz40WFzcx6EADNEmEr39QESbOzq0JTfDkvkT0UBVD5bny7wNmoXRaOyjbpZfSFmFfsHktITXxwHn
sPCqh32rOKMsEXm/e8oaF4Zj1sTBz2v/a3sQuFZ/FclzGxLP172w6fDS0RJj/Wb4fR+gMpotDhRa
JZNRMD6Mq03mXJwJMJTA4zpPValonfBJIAPu1q0sSnMGc5A+aluiZG+DLnD7SL8JzHVBTeolXKa5
2iv5PMaw80XUyCjjfsn/RCjxAQlnuNz4SAY13gkytupGjhExSaXQ8dRhq6ggd/oT4JDquOaODqjO
wm1RmbDAC5TY3DWoxiI9B9fVSvUZpoJOvQFrBl/Ca2uzF1AVFw6vwX56+jdJj72cdwF3iunEjhsL
cXMy6eKezxte2t2Ez0LGPDKqvF5samfdTCLIHF2cvKTK2IftcxotSEbPEN7OT3ktldKAEC+Oul3s
T9p8ryKMQo2fjayXLYZeetmDqvciuTsERFd31jvxmi5Y3UuaMnXJA/K7rCV3Kufl0rgC9fHjrjCe
bv48vwdRC5xmwQ2zo3uAzhJppTutrIpMNgf4v3e5Dw39miU+fO2aA+8vVLpbgaDk3aG2u9T0pag/
wfvI5SEgeT3hGcsCi/FixJkiiURN+4ixBfH/sEcWjNs+ShgVi+2+HulbzNv0jucg4selv4COxkJE
KH5WNLvJ3CoHmyfB6eIkCOWJL3+c/jIzDy5Fb7XJDSqb2ykcHTsB1nIrY2QIICk6CCA9cGPBr2Sh
ftmupr9yqcy9B/0rIY1erGLzOnDJbCKMrLvhrJs4ZUcrPNxnktbb/a/HIqeJXqZBnnJzWI3XnDkf
4/gLN8mZ1pzIGeVYrBJELs+Lp/OzlKshqWn36tQxyLZFcvPebQLnUqXG+fZQqhpT4107nnVqo+5I
E0dNsOWC4o9o40xpManriPD8vtczi41+lOEp4qVKIagUlZZCPyipdHqAqtb+VaibVMlmav6JIMXp
iN5vOvcxc92Riiq/zTZRZ++EyX67GSScZWiKqqa2kM8Dh4/PMeOjOmcYK/S6ONymLqrwqnNoYhli
RGTL/8i1vQse1S/Md1hVxeFFCKQfawv26wTi7Hp+Na4tuB4lWEIasrSENDvxCgn8gyFuDLeIZKrc
SkW6+WxPO5Mq3PF9Di0J1ONy96bmbg06db8A0/sHjXbq7QcvgjR5PN00NiNNQhstjEcc/A7hw4jf
8cIsdPOdIOhbQLEj/cPuPMWkwjKdg8+ne5b2Thg7SeSxoJWgHAxgMjXAUi4/QToWc/wCsfVBcx6f
g03WS2TjMe4OqhHvdYqTbqFTH/5WsPvkUMIA5/cFe2+vqCdE73k8AyIjo8Cp/fkfyk9Cm//+gFR8
Mm4uDsHhgE+rDFkYIYYA7LXnV/v+Of0+yReweKKlboNI/fuIz0v0yCD7uOQG2r+JzEQVBAnbL5kv
aIPUGPtWJm1iPcStowj12mgZYkLtWUxI/aPcrDtk2BKSwBZPIppcUwij3L+kwh4rKPBKbiLnx0FG
lOF1D8kM7In0UPu9jp9kddhx94t5wQpNb7qzN154LZat2jKz6bzHBfwEnXwHqdNyQUlMo3xroR5o
d/9CEySvDQ6SjIbDTneEm2PAoCeujs3CCaDIKnI10EaukTRZTAieBvBn8yDxsEavYm7yH1+s9egi
uZYyG6oxIG/o4bVZ5fTk/oG6Jqz9d5AtRr20flF3BYJ7mCHhjNabGwWnQC442Q/8PESRpjpgX17u
YTpT5cdet73BhwvOrAlTsz/vvpqjuS0WmPhqxNCUcf1Vk3L8/G2LmFtu6+daeDxbrt9w2sdmiQ4o
gHNRzY+Lli+P0qWIOc8DcRoLg1KEjP3qLWRCArKs0m/RHX+L8v5v/M66Vu/rVTz7KqB8SMyjhkyB
icHSlDkqKvGD/1Ko2FzNm6NtV9F+hQmP7XHFwYVXRozIoXDD4XWCb1Pg1tGXjhQGs9gz3X5NhJY9
3FzvKuLhFq92CgZbVSbp9snBoZizfmQB8TVpBcX4zHZda/WyfNbV+hJW/NIa4zyXwO3dTEDrkheY
FnsUMx7sLVRNM6dvL5FKzILcyat4CfJogHBO5NM15h8pOSI5HmygOqnKkjDqeX2N5hla0r0AQYIw
SaaLMy3ouPnsXIpbYxUndc8fGiiu+FhsOHA9OsxRcG/wlSjYDjWV/ptPsuYEiRfFLL0DyjzaIX81
Xi7tfU1iEgs+whOy6957pJHsabYceJarwHxdqPgRV3I+9/hm00/7C+m9MykWKzGtM0fsM038ZIvS
m3cUG8nHvnoV6PODU9dma8DJzBYzUsjYD6ZxzxeVnqwfUYnhvxr2uN14pm0SYQN6lPxYJHm/A8ac
xJFpwgqRJkzeOnpN7zg/8PBfxNoW1nYhvlYEYw9RAtztZXHzwiYtnG2c8IG7uqrIviZdgy2prqQs
MiEjwqcRsaP4UfWinXj68QckcJiYTXWplMnxBscGdqlEYKnGRTrpZ0tecS8G/+EfyX3ZU2b28xz/
PfCF9g7PJpJ1cuPQkWTUpgGu71E/uOOZ/U7cFT3fSTy2E4OcrxzUQKR4qgf5q8JSmZwIHHp/7Peg
t2vN7cuqS6KHXRlpOyQKs35msaMdJKWkk5FgaINz6FPlR1hqpfGOBgJyB1zzFgBVScrlsKBIXfhO
yWMtCDocaNzHnhtCsOXaH8lczZSCevxEP9dx/l8xRPaQywYd7eeEBlJju5lbTdPxLiNlc81s/Ui9
GCYAUeKxuLLML71Ypw+iM808lZ/BwgDS3/iUfpwQEy39rOb5qk2g+UWkendyDtstTzD2CcbZMffd
kAg3ThQvV0HFlpKMhkI/R8dAzbdkfpBMkb4R8gwZRN4QDlnAXZb0zHOxSRcAXjWVqh7lAuQPt509
l22wfgcmkhIm+hTWRtdRxqwJPwTylMTebZwa4WO2hIytvJ7S7tLRWHKFwYtGicrwcg/IS+KsfaQC
F8DzasNuS17LSaU3QgPWgbvcA0NnCsL3HVv/4oW2v1YHgPqSGQQC6Ex0xhoza52JmQrLPKEyN00H
vsRdauXdzqOf/XsSbJgwpQwrhOW/za0awKnbXJ/kc0Yo8SgeCRGFpV1C4xFGtLG2/2qa6dNU4Y/A
J6Y35/SjcyT3fauz6kTM0gxNEF/x4hxaEd75oNCrth2t8Gjjc0hT9QWNFLH2FuJHdxlM57qmcond
zLlJprF1UOxd9DL1j7Px1Q0orP721fFsv6vB7SIGMZoFcR9jzE7TeV19LMtW1W3keWc/QKoiUR0c
1VEC6MdJrqViUrpPv2tQMxxSLBmRwfjVABgmsPyXKQD/Goh18urKzBWPE7SUQ7VFDgxaz18rUebS
MaeCh1GJEElaGneVQ8rXPdtkAGknt6O0MgH3thcWlDFhwm4hHKmq10YMqmamDBAhbV4NZVFyLHlA
KoUWwF8H/C2V5FIsxmMyp6FJ2fFEj701U2KxtMP/yfAZ+ahi4cNzM1N+RGR2oayalndHTPJvuNGw
rGzOw5M45McyLIhgSoE+zV1vBwsG4f5XRkdhCilJdP16++Koo23azE1dTZazoiovIUx2zcp4Vs9f
4ZG0ZeVM+Cq4xz/0Me57e35DDVSOa7j1c8UwV0Fomb2HReNV7L8MMWxYz3cI8leN1JXGLjXeq+ip
PK4e9l4TdaWncrQtxvmosFg+eXaSi/5H13QD0KmcClOjgzpcW6B/ePIF49H5sGZXe2a0NUnbIgGC
XDxOAwZx4Gl9ko0SKJxKbQoDvhDOJNVyoWXSV/+Stx5UjuRV5bT59H7CmWBO5SZyEExJgPMDqOc5
a0PougktnrHwM1HKIlhT31sEHamLK/vPsul8eUtZ7LcbMImUDcKGnwqPpGha0dEK5JOwAP15ZhmG
5QzeyFSaZ/dOqxbPZLYMIU0ioTR0c3gOmBqRmfZ9RSgqJMIeNAG0HU/sG1pbvNlECHQFMgaTSAqs
jDna2BVcgH9cdvdPpeud0H+FBICemMCo3ArxW/VMoPLu0uGg3JlsXYaT6YLsUMfTs8/B/Vq3LJbG
aSjiSQerWASROnlp6DmtnBgu/c6kTvH/9A/P1OUGlWeRUFgU0cvC4F5JooljJcZA1i4+NvC9z7fV
mTfEm+Tpci8E+Z+y4RWE6KHOmOS8SXHGO5QR3Wjgk2QvFw5a5br5v4noJ0TwD2Xa6L3+Py7L898i
17o9z8OOuXybq4ezHMOmeKnW3VF+lMNp1repOQyUbRap0nCTrhXLuhEEVLIEShLe1oWmbuVVj6KQ
m5tcvuWDOMKYgTgapINnZ/ttsr6NPC/Moh7jRS4PqHWJq7iJhocdHRymKwBAHy6oQOovfLorcXB+
GnjFqGdg1GZ8ud3+Rw5jjCkc1YuafzB95FWrYc7yiiQNTrxx06oafG/w093rgmHT/gSn0RCZUtHZ
9ujAFF40jG27tw/pTjHKhnNsJc2BE/CXCFLEmfIzDkO1uR/bmOgQqB36O0AnBldAkHTqhnA/Gj/h
YW2iZdl1mc9w6Z2oquAhaGSOLXZ1UWJu27Z8yspA5omXQ1FU87TIdApnvkMW4p5GaTrFiHqTxLfX
FdcCnb+fZg8RxE36yPZFRFpHSk7bxz81m/YgcM07NosHULP9p/bGVPdYe4BORQcZt4SRQZ/ITdfr
SgYrUj3u7+9HQa6QUz9b5LVF8vdZcOCIo9bcyJmylFaoCDO+jJXzCV9g6veN+ke9UVP1pU/MdZ1B
O8Hpgb+3wvx1ps6lNffoiXBbJUSQvJuhRFoM8euiBVTBwtreU5VUU7METI6ErYfuKAwN5izmxZKe
NLxSjS8uG1Go1tX1o6x1xMnCS6xQFzBi7gY2hGfOqaCJ1UgyfvfRmR92ObgsDxb+Pc67FQjV1LJK
4TFGqwMQ4KMc35W3CwlxeQGF5wth3YyO5Dkc85CzfBq4tC77qzmsmdQpCUiuszQ4imNRKJo0Rwcc
9koUzIXzwaDxgpgQZE2Up8Aas790BIXU5Ldhto6kBusIZ5zfjU6yGPhSHudlZdaRsl0CGh/cuaa1
xR0uafcaEe+yQXlHOissTp46oi3Doh76jCNcb4zNooXVqUyxSnDcYdJpvHdTnvLsW1aAdp353MwZ
MEjgvR20c/miBCOnTWYr8DWu1OPbp2MtNBbwt4L0YNsZWulX7lOjYXmX3vZX03LU3wdLEOKodQbP
b8d2+IxTMk4Eq1W4f9ThbnaiBXWVMuv9tPZEfEnXrLIwp6IrZ2/LKnAbwXXcDiUhb9f1tnffXKSt
hc2TB9hGswGxLITrtiuEq6/h9KVA0M10RZnPRLh10FcWbkpCzRjWWQenCN/AX0iK9MG9JnoyvKHF
k7aiqGgn7yEeyKWncr+TiCCOAiFlu+L90zZ9x4ftWPlQtQyVZz7EFaOimfz660kwQfqfc4Fnab4C
t2E9jxFaYYlkp6CH+gFzIEgbfoPr16Dr8l9lmp2YMgRimCu/6IZawk58jvtSZl0BdVYnEtoNFO38
vuqxGomlisDRCOR2QC0gsQMKPfX/86Tu7XyDx24ZIp1OUAAR37YPds2lMpi067NDHyg+7bSJltdh
jAyyc5t7iSFZR6VCHe9g4BJck8qpMlgYZJ1GcgQ1R7Z7HVmQwvYzlFfZ0eII2ChYRFDYZVmPUBrZ
sQ8YnOH3zGPhhE1/vBmqse7XDMBPEe8mNbt+Tr609munyWa/+v7KcJffHxf1UOZtS+AZLfNjW8Zc
YFr7VRvxlPy79AGZGQ+V8YQ1YnofB8D3qhwxmPTNUp3WjqY5uSF7goFk3c6FARTjvKrpBSVmsYHf
1IJ2IFLteKS1W8aadWjq7fo3AORwKnrKAXyuVVyB0uX1HboY1mHwP8lf5TZp9UY1B2pcO/kgqGds
jxpZqsZutEwnhDB7yVusodZVi6DSMi8gHQ7BN1FV30Ij1drfEaWQbQv7hgyW25SIdp0JTmQ+xCim
tg+ToK1ZsLyn8yedu+1UO9IFHkvFtGdgI4ueXB21+6gbPDBG0iGqDBe9cApal2Mu/LuHMaQxZrKi
tl/07TPSK0Je8qGPjvRH4YYPhZ/WY4oZM5WcxDlC5j1i9/VQtQ5Bk86B8y81cwscgXmspJD44i9h
HbXoTGL8YR2r4ApT5s2t9oHHYKGzKefDz4O38rLxh3yOoqAOqDhrZFN2Pe+0uqK2T+ecC+uceBHe
eUj856HJeFR/gER37Pmy2gJV7r76vAIW3HrskilyGoHWOJk34p3ct2LJm+kMuFOVReSCZ+IRSI9V
pUcNnb65ZgQW3VeVWDhdKPWYOFz5MALykeOqImodafsYhC1hPBxqd5XXJUxREIScoyq6KOQdcj+E
Ji74YJRGhqjr0+WBhy6Xowr4TSqdVMpkMLOOTycHDG2WSN7NzgDvm53bYt8cNW56SSJvtlzCJyUu
TW7z+fSXKcFh/BtNnhBH24qJvgccRAsF6jI1nE0nAJ4hFJoXzsh08z6Cpi1c2ocwLKswhp7uQIZv
Bnfq+kyD5UljFuOTf5yTf62DAipe4hun21hR2pWpkfQhN8B/G6tWZtZ8KKVrYhtyx0pFuw2CG/PC
0/kzsHlIT9qaMdN0OrJENSMVBRWXysapPMhkr0CgmrL3H2dRXSydQh5hlVy6re7PrnwUevaxXNNu
cBofbr+LSTjw3rMRE3vvaFLf+QlRDVZOWGDcZLP/advsS1LE1he1oJDOLn+hFAPj/SphyJTjWdip
LJ+1nUeAOoy1GobgJJ5p8RpVRFJVv1WM2GDUNBMeOTRR9XVCOhFIxGNTqmV/KhbsvLWZYrEZjial
Er4BmDmLSF7NlCKa4HBQICMtU8gfySGH+Ypo5Znn1caUjptDb/WXTnuhhteEJBOH0febjEJg4IJ9
64yyD88SOJdoBBCOTCXSxLTPLcBxf/vAknEDJuUTCR0J4PEJ4lziEe9DcaKKhUv4fcAUDV9SL4WC
OfApuiCRnky6HnCylRi1a772trZSH3O/xdCYBR+LvQ3HK14a3gHCXBYIEQNvmHC1SqLRsnr7WmKK
wwE7Kn6BrFHXQufZz6lju7pqYz0THYgRDuGu2IdV9tW7ID6pPK1Lo7VImEMKSGSQVqCILpnBeqGe
Jf9obYqmYfDdTttP9osrd0JqFZGfUHY+ArYgLr4Rd/yrApWobYLUzebBZMugEiBO0aFnBQn2zhFO
fas9guWuYZ/ges5JrS2or5dEYgJg5iZb7WNfrcmgyoXCocAJkEfcr9wNM7r0vA+MGHnGSrHPDBhC
FucOSsgSHQUSottP3LNlKBlE/m85hnVX2PYKwxihCQ/hBnYtaNs00RC0YetW+SoczYEYxG2E+xSa
FpTjn9cG/D7BX7yF9Gr4xWoxBqcskYjLGeFI4ttd2Hj053NmYChGIZEjudGK+s1bVbJqlcx2zjDj
1/jCvGgKvxj9ifSMKOarbgagBD+KuD1VJPCl8F2DEWWT3u+ZkfH9KLJ78MsGEjMz02ahD+nPr9Gv
/kmvlKRuAsxdAMSQPUOUceCB6mcWCVfWOXeE5Hd10Cgoi6C39b/ngJVTRoyVA8lqDlg15BSfC/lo
1LbCuIK6jTvpdKA77YauPJdWaBp6cGxQM3LY9OCmQaXPNA1vYfQuutKImL/MN/1Q9VtrWJlHTUaJ
uVzxJUHzdnAR4tBJOutw++B0PDrcK9A+sIQph54dC91VUcNrRk5IsgNzTSmsUUdy4X53tVHxSlgR
pnyzKwKaonZ4T2h7C1j6and2nFzJMrstK0whze4tZl2DW9IzJDcYylz9iqTIbnLzlGDllaBxVh3u
cpqSAkAvjmy5y8JyJSq3BT4XgUbtflb9yrEHYsWPad80ogjf1LK2T87ym1wWxyGZYmvq8hRXeIgh
LIHtlR+2AcRXVVn7dg1mNjWDQ5rVp5+ocuWpwZtVOwJyJmnQfUdynvXWX9Lo6tcgnyRLJ9F8XmxE
Gb2O2Ve49ozpHLZftQb9k+5wLbE/ogPJx9+VuFRlyhogE3GsF2TtWiNxMIqC7X1uDReXACuEHmiG
ie5C9kZuc2GiaQ8AK7IZM12wk4j0rhRUe5RkW52TSk2dFKs8pnNAIXBOMosnSsTk7+Zvn3lIb1X2
sG2oSMc9gIZVgfuY+kKMdfqJyed/HDCq2ity0oATQ5FLitRzW8kJFGDjZD3MqimaSz8gb5dSvzYT
yDxpQhhrQ1l6cQnwwTZNAa4JtjV5sOijkJdJqo7QsxUKULKVJTGmmu9Wpc9I2QlI231mv+D6ar4E
3mcmyeld0owopcMbyZXZyEzWUzyzD5F6R0fa5U4rReur1BkWgOhZwzwBALkZg65kO2refT5JQKhg
VBaSsOVPUtdebWxPktWPuAznFHN1SqknKIh8YjFYtXMe64QB/EO2t7JhkH9deNe7pK/OjIdFme6M
vDDzaoTz+sibow5mPfcLQgrMpYezaDTcfy0ywh+AX6WITuD4WKHttEU2tsf3MJ+tPsqaQRzszeCd
vMpk4mzp5aWJiCfOypZSpDXz/Kyq+2NJj/L1hVxXH2yKL6Vyn5SzXKQv0zY3xeQ9LhysaaZm0569
my324YzhjVALlr4x1w+Qs1V+PmBZ2KxK1O6F6LBGu+iotdyInoKr73xwoDxfaUhYytpIB+4RI2QC
PgW2kyutsBItqaWQnDWOk0RGPpoQEXEzMEFDZvDxKbsX8miaKZId+5iuJjToPWyz5uuwRYzo6s4T
eLQpHdMEfqtPhsLPz0lh8eNjwo8i0zPkJ0zkzixYHYSpOB1CpqqTg021ifOfmsXJTgsItaNbPKyQ
ve3PZDPUnHwHfAbS0W5Ij5HyzRAaK5olJR+dtU7TDkv1XqTsci+FToC2iPsl3IDqVu4DTbfvxwy6
YYv6FuRza4fABhWL/FJ/R+ku6t8WakUzjHsAVpbyHThLPOd4E539mYimgTWVtRoa1er0pCMUTmP5
kVeyeoqRMHfIJ6f6xOOXayeQuoF/9nk+tPm/Gi5PC1RNeSFuup3OY8Z93xXuhoAgJrsrdAD9P/kZ
CjvdxAztrUlC30voI9pFehlce73yqEQk2a7uXoTAUIDpA60ieKxsdQ9mWdlHgazpnoVRftw8GNcw
/Vm1S+yWuMeAUnWnXs8K/2qS1EwsrTHZQciUzra5Ml5/ReTSHZFqZiZCXhtDhA0KNLZC/90KDN2g
wXMGVO3RuSbRueiy60CF1RcFu84TVDEZ5n9JCEZnMlPee3a40ert3pD/XBkyNKETPek3N7hX9QuB
fItxhv/Hynwg6qtr1LxbOTtGQ+8vZiyV7RKKXprBZ9CVZn6DjzX2HPXzu1eSBDYKZ2z/KcMxw6XP
uDH5pG3d7T+d+5bzPJktHCjiwqHxLy6b/YQFP4NOEYxBeI86TiNv0FAg/09vH2kon13D0rXqwm5Y
VW+jgB6ZZ4AcJATQSNBu3h+RcWJSSx/CDyoHvX8i9UFTYLxcRJgvXO9oCaaDCkuxbddHjXvdPPsb
lyiWnYhUBhKpIBG93Y2UTBGy/mu5hp5rQKNWjiI7hMQkLUjp4vb5uf1IHJruw7kD4sXbUwCjnzZP
d4mZC9GF0DcD807gcW2T4FtyuRa4VcvYELM65KDCNajViz5e2KdHLREyLGzm4FqRVUdYGQEQHtzD
da8/WAzC4QYPKRM3NCbb8qTUgY1CF+ngAOtS3be5nf2dBPOsTRfHgOo90IqD+9vUpxDwKZmfIhsf
M7K9sBHn2ybRXqPrHNNyNR/Yjik34uSVkaQtBgTrRmC6mPoYiuiJvBz2YY2vpKVwtA0KDG2YX5Cy
e7sWS41bwIdWJjU9qD8HCrclJsWpbenIsDxytC9lGYAr1xAGyNBvfHoCypriv2BVr/gjSGs145uP
So+iyRNRqTprkumOLltvzEYnsms7snBIEN2kSdb5vc1Eh6L82ZK5lJcluffMk2p7OHjyee1JzQBo
BTyRw45soOOOizMW+KTHkcDY4wYawWBd7WtfeVWHd83cf+6OIzCHT5Jvdq0JbuMOGjnKZ42RTzsW
oKWmBz07fJOL2BfJAVGiwBPgmD3baetC+1p+Q1WloTlZtD2H7ah9ZEn7IBasZzyg/JDQxaqVnlhC
n0AZVLrizOxlZEhCbqKEBqoBNq78v0emrpf8FbXZS4qbm+GRdIWzxJGnTAEgKyuBsKEuZ7VuFhqn
9NeegmsWAmWUwQMP2FfL1q0OuTw3hcKS8YBDwpRJi98N4kbHo3csKeBRTv9KNhuXiI62FVuy3V8X
sgLR09/rBDGpb7072SJu9TDou7uWA6Z+afyJZTRjmvL04Ur9us0P7/oSwSFygp6asB1i8FecOQHc
OY8aJzUa5384E7I9G86tztxxgQoxaQH1m1c+gE+skmioY5Yv8VLJEjI1AyTTqwWcLfXXpxrd/stz
AgS7pdqfgjwXPuFP85SJQxRD6Jy1vMF6b0aRHfq0S005HXqdN1FrqXtG3BFAcfu+wl5GjCzwZxFQ
kZ0VblK0vo3JC0NvmXKpIQaCBVzYbICY214Y/AJL27PGReeuOOKcVYaHYxsveC+CFADCV+6lq7Jt
kj1BI8jQ0Z4e3UXlTcDYUJPfa9HnDIjb5Pbbz7OzedLhT8FFl0u45FzNFYj+XuS4MkIqqoH6hi06
C+ePXqfwW0VhAv6R//EPvwyxG9iXek1XP4GcOJmTwUgtpZJqjS1JzyCbwIRFIWpFoKl4E+wUh8FC
56hhVtN7Apok72JhDcWV1EMqjy4G8NpHcKLyBxlfEgETKvs5Wbe751sChKohb4s6tDqIHuMOp9Rm
uWsJsU14ofPNMX12uJMzZPEa7sH7yWg7oEkLBBDA87LjS3Fw+cpw88EBEDZZeP7SeLJhaYSKEG93
eFElVlETV2rKId2YfVlSlcy/Xj8wOLk+lrIKEd3+iFO5T3PeZP0YEEwYalxqMkAJZsHrraUlp02j
fuWvfsyHZA0pDDgQeU5yUJRvVOdHV0KlIVEKvr4UUsDlplal1+tmQmmK5OSzyUEPqDo6QbssrH3j
uVwyD+vvK8g0XYQD5tHbX/sgBnHc45h4aHp3pG+kPU4cM6M/TOT1eGnLXDgooWASOU/rAznGVK3K
uOGb7g2z6RljT9bTTirs/qKj+mKuRdyCjkXIZWD+LGz1y7UIqty9Y+vbUIMgmhAwNAaIiySDRVSL
oQgwQiGPg8k0OP5fztF3Zw4xinVyqlcGKHA7o5NUHM9cz+7ef4bygDSoRHbYaqCmWBGsOf+EWZNr
XcU9K+gTld4A2R9w7Ir52IVW6Ge7U+8fPAtTZdPekkAEb7xKKNCIqnQ1kvJMw6hU6MHgz+DHZxmF
0ElbIqcRshvo9/Oofo6qtwJRyGK0Sct+BCa2aAuQ0YWAuLpUcO5/dZYYn51Aln+70CsiJ3RdHqyp
4ocBN+7Q0sczZZ0n812M7WGC4Cn7w+vP0itEq0k/XWR2x3110W3xJ90dQ0hAtZl43+bbIUekNLXG
TeYVolQsaD9oLnc0NRJh9FdseVWSiAZRitmVycT5ovGCWCChanvokrwO7bjBnXLNil5uy7RStweN
q/sBr7K5X2PNUt8IUsBWcZXvVRHKoXYbs1v/j6lkMNqHjZyyvqRLIaYp4bjDMjYKnFYIED7xAHaF
ylPMSjHVgi8bvgi/0VbGL+ikAcvH/X8z7IeFToT30VVmeeHCUQ4nDpNVDTvrJuVIfwYw5bGsZAnr
iqimjXI2jS+nkSNE9nvx0FUH34hisLALBSzBDPF0RSd7h/CAjJWflUNf4UP7zNW7+Zi2kPTxFl8d
MaKUJikmIEBXFh/kd9JE6Z3c9afAaUsmB024QVnxCHDBt3gyX0PksNnScIW7OGp4pnlXmkojoD1Y
lRgRRal0uHv3FGa8FfFkl45ubeKcGkXKuRgZmGVjPWIYNkW50JP6RcTrgX/c+SmMnqVzd2VkUCn5
RtyG6nF2wbaM15iEZ1sLBpn55j2y9Mz632uW5WYZkvGEgCKhawAVxS5qqEZZ3WNV0J+tNqAmErEv
vJa2PZELMBi/ledhB3xmA9esyXmjXLYNo3JyGmj30P0IXQpMBR9P1rFMq8GLHCIGX45dLG26fear
/DORTzjzSwKayjhIA98AF9wX7d3HR47xQdqNyxETl8jB1vS6GGOZKPbw3CJX82AknOTyjEKF74uR
hTHGkjyA1rA2qg9NULg+CYT7J09VZkzwqLlD1nrhTiRqGmlaIyP5R0yU4GJNmAH6S/hlju9K5j+u
fHNBfJg7f9is2iBaPF7mhYkUXSaUTvAB+SpFUtO/wpi+JpUvjL3Th/YDtyGcIdPhZsdcKn8zop/W
CTXHtNZbaJUvHCy2tUK6JsZHKhinTLg46VBq8C3exbMWXLnHXl73PGcyrsa7pdCTucYoh32cQiwi
HjJBr1xIHYoaASg52gUYqBrectWoicgLfHXi8l3qHD9MstANZXv7UPPJYmEw2YvQ3OXLXWu8Toxm
no5U9v8ndpNA7T5ad36ZfYpVeDzP2GQ3JYnkqWnA6FqwDrCqUD1kcxRMxYWJOUKmozIyPPEfjBxr
ND2jJfI8qBRFqdySzizVeHLenvOEURUu2Po/vMwzU956trlf3fvl7g5ZlDSCLtyYujz5JzgE/WJ3
Z04HJdu9w1oWclHJoEgO8YwqKi/XTEpmrJiL+y1+E9NuaE08T+R8kzNNowdpcl+SCvdjBcKumtV2
xjNJkIAjjv8jH5jxMJMcYKSRP2qXi4PRPOkdPUAAawHgcg1BjuzEli+97mCBLlAWe7gLDEj0/Mua
WoapTBWUggcW+pFhLh5XkLDeQTj4SodgfP4uYuJKC0XmV4j4woh5eapt/DxqQo63OEOFkhlL6tUF
dVzCzQ+z00Oo9EOavS65ZvxDwSFwHwP1lrMJe7ClV+P2bjm5V9K2GrdkKUIhQx3IwIQUxmKZkPX/
r8qj8nAN5kJk505wcJ2x6wBdXnR4/IThNptZQKQjICVZgANsQ7zXJ0oCT9xBlb4sgY/Un/RKvSlL
dv7dKl/DrK10Lc84aFAI96ktnytknGT6HAMBfcLpQoua4/pofDBzoYPV6gsCqCK2pJ6nqQGBSxFB
DSGPjV3wUKRgQMF2qlMXT9bdPzDRShkaobwf8fP6HoGvtZCcZnCIoCfrk/nGo9WJsO/ZzqUASx33
Fs0InLzu0TBnXNE5y5pH8NsJCvHa2fI+h4eZiicewgx3+KNvmNKoWmr6TkURX7s2F+hx12GtFK7u
wsF1iPrFS6SKcdXLQwZ1W30AGv5N8jRpQaHCHJ3eqfmqgiAy7YLBCZ75/mlKjb0zenXdL4/y1d8F
1FiPQeDiCAQDo4Hgr9OuFIVm8CFi63RD2LRSePAL2m6WhVKy18NxbfFeRZdSwKYBlpM2mTbx+OxO
xQzlFfYSe6BLQjOaYC91+PEgQdvOOE6mMbuP8F9qHRRcPEQWhnY/8qrBRyFopjN5Gwg2NtOLAMyw
0exRwgeyQfLed42ehHUuKTXvm2ZtYt+Ny0OEYmbmCXuAjQBarKYISfNY/0Rl/gsJO9kTt9Ytp7Y9
Ojjk4dPNe4w3FI9Z/c8Din8H3Rh21h0zYk1AJKywclrOgUT9U1QUWi6CbS9ASll6MH6nIEGnq95r
USSxOn66X6INGRlmS/L63Run1Uz37+sM6ME4XccXRpBlzTiEcQSLn/ql/CNNRqXj/fN50H8rYop3
hUldeyXU9k6/hOMw1dQsNbCyMdHEUXJvm9BJ98ZyHCt2ZeCw0tiaZDLCrFtLSL/uNuz0nTHpYB5G
eLvrVmFmlbWIrTl/e8JYPhGpdeNS6RK5c2q1NTPpvTGBR3ZjgoEG3h1nUDHchiL/w+9xRrNBLyiZ
stbKsNij97faJYhm1dOmKppn0f7UO31MbjhQ5XkO8ZsrOizgj5WhlMBj9s81GBDmXX8I7ul5FPwm
1DBD/sjBA1FdfD53ORf94quWejg6Lwx0anpYJCIma0rKFzpjbCLJbfcpcieoJWjiH7uWdz2D8jld
HpSW0tTR1KyEopssCkaIVJJNw12k/4xwGprxclFjvSFEkB7deukdf3VVXzYVryLjXIW2AmHcH3D2
V4ublgIIwiXLcxsqvoN5oxvGCWjF4b13YS7CHfQfQdZQeJZO8NMzVr82+VXxEg4AIjqcghGNZMCW
7Rj8tYpFaxiDh+sr/B0Wg12s3UPq6b7QaEHul7xRuCex4F0BTKe75oDw9DysqGIuETEraQf7XxYY
a3ggQv+bDy7tImcOJqa0mu626q38b5MF5VUA5gOK/+qzZJKMOSQmSCowaeyWsdmT2pymQe0ZHPqs
BMm3ZHW/JTKPZo6cRc2TIaucdqh15gjGpf1W6d6Z+J/xN+LJ52eTgeL+q9L31nowFc9RqdP1hKpP
4MTMyjsZJW43BzBdjXDQTWMPcshpqt93WbCU6rFR33OHtIy814cxg93iALFOZmHXPuqKb6uRzIpN
gFTy11wGUBRhAIwGgBOQFr2husQ8SYphDiDKP3B5Qa74Ml+Cz5mnPHeoJb9Ct0W9oNLz9bIWOs73
YnRPgETNBOlSnW1cojSPpc0Pe0PT/Ly7u/wbsfIlAk9EYa/618y5lVVhRlTHTVb1CJyQTazBbPzC
JqQ4Tjwd2mOiVh6nj9HcWkSjiIRba5BqCH0aHFkDw9ig2jnEICz7SxhwpB1jZoHApvVcWN1lDX+s
qkOoKzU4hbTRuwMmfzUpfWdoPKuV1Ge6iOPD4fiKjIWxwKYXBXNMaynGh38pOZgyquHOodBWxBZS
mnX2aWIOSz1Kufn4x9kqx2Nrt46E7ZaOs4B7+1ZUDoHEmIXI8P1uhzDYDEit9mRyX0Pfp3nv67ZS
hTHSzH09RcPHrRBi8nnn5wA+6zONjkDlEi7Rgj4+MF5cwbO4nLnQlSeiNMGLtkqDr+zgpREPoJQ0
bgMvRDfO1ye1JBc8Wkz9U8iUsMrZP1zLi3XRiakpVRnYL0Ii/zFgMW4l3nZ6vq3hAfS9Wsb2c8IE
5V3cA45mmDeazc8dZF8YlIpzgSt8a2YpuDknke6MU6R3F9xsxGypN2aHWWHAVY3EEtLiJWB4d6jt
heCrn6Jae0frZ0j7Sksmr0n1+7uitViZl4FCkojNnIUwasZyib4AEf89tfu5o1fy4l7TxzH5Gf8J
Ol7+WDRgiR/J4f+MiObQrpK8VtrCl2/zxMBDwYrlztS48abmzvX1yF+zHm9KwJSy90DfKCSo76/7
5PSWIaVNpHnQPp1LzSQeRHsQRZ+T9wLydfSu5ShWGozZEdVzFdyIJRxarDjC3f9nhpbVWMUd2JMM
cdQyGSYyI39wr2pqS1eHB8D/Er/62jnIPCRQpHoAPfGnUdPJZ/O7gTy+KJyMA4Rl+E9cBip+onLH
TfAxVDuE3Ce+DTlB4Lf0V7ZMKktqpGY/in795orh2m4Ch4yQGJ+yWk7dE0sSvr81H+WdRUlg6MEp
zBlBn614fN7sOw7bTMUafv0FxGpj+coW/Vz0LX0oyHfOWg+DbAwvPP4e5NWZJ4Uj/SDR7AquBWI5
9FGhtn/uGmNJhz5oogfQk3Kl+R9ksHaYRBxYWqwqBvpRyPCLuI3KXgbDRlhaGFS4NPFddXmgdWMT
yu5w2jo1ad1YX1r0FeUenyd7ntuDuFpRhmAEvmRdUMo8LYQWwwmpoh5HWoXNkJnrVqIiDqyuxk/3
o9Wvq801tRPuzZbXLXvy1AqONefKpi4Pk9hSmemdR8wWiwnTUBfHXVgIKpZmwyP7PSZEqhWVJltF
/XHK/AX6sDo9XOExoh1KH+Gsmg4+AfbZ2seCCEzhUYMqCvCRzJFwnaNl+guTDOKkECDWcKvhcWHm
tJaOhKmK2ntWMZoZHs/lUUYZ4oU/7h+65dh9R/yzVauKnD8UPxItai9aVhQE387ePRk8Kh1WA+zX
xIJ1PSCxQWK5E8X8Yo46Dl/QL5tnzbi71Gc+aMReMwgvtT5cGmqJbGvKe47/fwoxj3/H+T1zKa16
nakj8Jms83cZetw+AfqAt3WtKlWVqR/RXHwD9cXMeLJBthSuXC8UFa/RHBMtBy62gKFVDsngFBt5
zX9XMWYQ5Y8Br3y5NuT+KBOpesFuGJlTT6eMijtGKLIV0CsZcu9thjpEk4FZjVQ19lVxnlel9KQq
S9lJ8Kfft0o/pX6IlYyzP4kdN0h58WcdpFZNSXO0jt20OSvg2O7bHSNwcHXJ/ndGNj3B/HDlfCeb
c0GnRYM2e4IkVhOZkAdxBUVDfSMtE2LSQ+hCDhneXLexLdnkhtG3QqhkfgIQIQJvZQdMnNAN8qxz
kvVnRpqy8z+u4PSmrVsGsfNAdZ2ulk6SrD/ncpqRcKrN7urgddyspX8U0SP3JSSEaoaPleEAb1sc
vJLgK8pcLST5UciYgVshuhKW9M67/vj24xomPyExnnTwfEz0vErLYA5JQ9GT67uvUW/H/DqcwY4b
soKmutvuVNkp3a6immyx30H/fWhELfKmqz7AvYIzWH8ONzznGu5G918Y42wEiacN3Lt7GqTKjZGT
4msXln5iyVC8y9F2+Q6XtcoPJRxJjrBni0IOHm8ua/pqI1rJHDAdRcqX6grfSoTOlxZPISps27Mu
XJ8bJYgi/VRgEFAC/iiy5RusRQeJh/J1u8KqcCwVmQvOIXz8qWalG6Q9jHuw5LqY06ANaQkWL0nS
DqmN5OnrUq+G2GDrm1Xgy9OVocoG5STyDijTkoUIsn/KmMku3lbcwzoqhMfdVupc49JkfDXvRBo1
gIzF1NWqZa5t5F6PCkA6MrW9U3ZISuGiOhfHf1ZFjG4cne4vASZhcaW8J/BoL+5rD5WyMxer8jCe
6ksxgGM09DO7r+DAnc2ItD/sur5PwngO6nkq9N0Imii94HUhRLDJwBaD6o+uLb9FkWb6wFadf6Ra
Lwtye2HPe5hzE28b0+pEvL5BMvHuoShwn2jspeFfHdSx0eNOkjmhQHU0IlcOdkO+W7sgxKsvJLai
m2qFMRtbH2keCWPCZ9nEykFVxCY8bxbtyQB0yUaFCV2q/qocmbBMtGBYzEQraEcgMbM8Zzw1yiV8
siF9haoiOOX8gF8ApywHAmZNSLmEz7Ze8sN/ayj+QFa/zYLCEU+dMYxtD4PBk5w9lHVloJ7pjIjc
YgUIdnOH5qEym4BS4XH/KtV2tXwmhRlqeWmKKT1YvQa9MWoZqfLtKZhGp3hbwkPphrRI5o1WEJum
+teC0swfc521tvDCTTiHHDMeF4S+lhW5W/JmRnSHOMmljjvsBpb92nWnm/N2QzutlmpNg9J0BD8A
93PIHgEK5v2nzmtuLbuecJGeNzE0z36LFG5KTJbvIZNBbeAaXR/39/mRvibUe/FxGpCNcr+ARzoe
KEw+5SPMCb5ndOpYKppnvC5BfPf1C3xSvA8q/RQs/xQdOGZIL4yd8xZgOh/6bCE5U1pwODskPWcJ
pOJ7ZvINl5ljHmAF36HOWvv2DtBlRMXufLgPaaOPSqRK8ZUXd1AoqMJesNXoGhU0S1TyEBhIg/7f
b/9rLztEOvJflHg0kvSw2dubVsM6W99XdqqjH+MavUdRibNDN+Qi7PYSaUuHJ/eXoTZT3VfNVd1V
my4I2nL8+KBYS7AQYobQB/kd45IGtxtdRqj30bXVru2M2c9hjXRUYqFEHGCPnPbpIhJ5HrZPTGxB
OGuYuFSK6sd1y3eVVl0VtT8yjhHfk3wmBOXpZi6WAL97f9ztMDONP4N3Preo/OFm/x7sANGU438N
VOGcKMWdt9F88T/MgwMRWvp+TemzpfsEh6SCKtgOPA4dnHAbdqGVx2G7xXM1+R7qrwPEhS+L05gH
J+9aYqeNUBCl6gXre/N1YGJT0gdEDr3soACPqXWPKVfX2rWceIpz2bm27AXTk7kiZIwVKFoaEngw
lPYTECZq3BrvifLdGuHyCK6VR6G83bU06XSBpsNnfr0ONu/6DbxKbChn1zmGFCKk85vqMAG4ON32
u3yg3lNqTcibUmBOIYqFBB4070+vsPX0JL6D4NCUsvVG85pufMy0df8v0iIy7D66DWtPjqXbulYu
g7+5SV3jcrtCiN3beWD+gaA+dlv6k1OK/07RGK3KHoQNacmUrn6JacBP/LH3wnR1Bx0PoX4CqF1v
7ES6EeBcXyDzhA49goYHgPK98TOPuH8IA8/x+IGE++12xxPJRZk1Q31q2nxkwCTlBPkAEmGtKIGW
kULLkwlQtvAMeG8qW1bfWCJYdrB0jJoD4sEiDHjQ5OVM0nYCIK+ZR/yxtS1J5fYn+58u010NrE7F
4i4ZRFOSQcp3l4lwsjq71PpXEp3sYpciraR0132YHLQ9iyjYYF9m+gfRMojqw9m7u/yX0DK77klN
uNxq7tiF6N43q6LsIJNgF6wk72JFGrcNj68QU6kJT3wrgZC6Iu69FU6y20SuN/CV70LHf9JFUGpY
V+A2QN7rYCVAS/pmqYubNgw/ncbVeTNLKHuCudaW0j3sS+C4odviHOUXzbn1jCeQnouuDgxXEJbr
Ngn3MSVsjVOKHpuBSbTK5VR0uNzFJLp5AbbeOda0oxGkQUqc3FA3zvNukxSEesUinQUCkDQR9mS3
upE/c6xJ/9qyTt9keMAwleU+BX4LeF0pPGJqruNi1Bc8BBtu3t2+qND8EDHOqb0p4oW43Zi/Fr4q
jK93sIu5EO+4r4eFlJmxX3uTCNJu+1FYf/RkxCCanPbhgEqSdO48KdUSDkdt42bPNMMx6IbwwSWP
kP6DVOByPCQq+AwWRTmI6gtVEtfaUU1qfZB8MM68AmhtBKRNqNtjteQLu8tafVaX610bBjRPu3lU
Hdv3uUh2jPJvt5NqrpRye1UNsuYoQwLAp8EasXfJ6pqdb+onsFwiw5K+xLqU8dpDY4f3Ikm9o3+Y
H2FwYHqEU6oSnEyPJ/xysRKzObNhKNqwYATAosOnnuMutqclfb9xCMdDI8L9nMjAhuIZDCd36iND
KUH2o0HHi5mbLLcW5Ay1QlPswDhtLHq+QgYCMly5qfcVfXLnYuvwcsMR0UcaEEjm5+tM0qSknGZB
ZcVS/vCEWzRx+zO0lvw7IL5UJZlo65TgWQB4eMAD/NIQtYxsHfcMkdAUPOzzYUZBi4iI6eM+h5E9
2pXkzdQAJ8dkX+OprZ+9jRWGSNJwMSiSfreuYByQ4gyky6e2LyInsQDRrT4gETGCpyVZbY2NjqSB
9RRCgt+gCd8+Q/vHr+fRKR7hjJcKUdEZcz+FHBaum8TG6jBJhxm1dE5LbN7ecMoXeNsphDCqNAJ1
WBIJebsnXMS51qiFYHK7/QAKJ+9WQes7diRzr64vykC/4Eyuamh0WhYTmWEjJufo6iav4qNO3nVP
OPTTKUDG2JdhyE5OkxQVK8HSFw1sIgeMA51eIucFpWKV9nVf6vyCXQp9XvBEolbZRpNodsMV4iUR
M1v0P/e4L+tcgBAh8R+LAvDhf1XUtva9lLrF3VdpmrQjRkOoMD4uhbYeObBK2IYjaZBLptQexUk7
0RU3wD2nzXScTf+TvwF3evwbjaq6BvtoJLFcsaBvLhMKI5LQKXyFVjIOQqoga3dM7mx0+rX1O0Qj
xKGoMaskhAox0J78SnU9mU6aL91GM2b7ck0HaqwZemlLxdpXNUEQ2vmoXSZLc38t4kFz7A61HzL1
U5LJRydnLwyAm0qXYiTJU4+OpzBxo66KAIkn3P1mr/CQQ4pc+5sIT3Ba4kqQyw2meWY232oQdzxI
e4O/NdouJ28nqfaeB+i/q2nZt38Mogv+DA7L5k4MwOjtsaqjOoRQysMyvKisjKxopmfvlQloThXr
knGvL1nS26VMMPJ1lsDx7YQ4KGH8GLomz7gDAo8EpqrXn8To4+yrtob9TQeVM+qvq0MdUGcNCVhp
OwmIdP5Cp0RHy5oLS6dJX1wAjmhk4/pUatsy1MBRhNCkCx4fTsyuFCIIyZ9yhozaI3p82KkBaAWP
xJMUohdUpet7I3nbIty3zC6X0d5c3++gFaSxt/LmZmiXFzIgRbzKPXah4PYhKRVQn+2TQWGtLI/E
mFceg91ntzVJBuYCpu5ZEHaL0dgpoecw+TjV8nVhXNRh6I7LIgxTwZWWtzUhkFauwRhvZOPSH67I
V2iWVJTGKuYZcDQ4qrfOD1cIolZ/KRXKAQwrKULtmOzVgmgMEfT4ogxZMv7fxy3iIpV+4BNEQssw
kbLlukhE9bq4AxfgxszPRRRkmmEomrwtUGt2R4t7GwZXnP+YC99Jgqu1wazChZRCvBEwj4Ueentq
i3ECsOEx2aGyHlI2dgK36ADAjRNCNyMY9thvNodOuG29habJE0vJq8YlqVVw25WAt+kKCQ2Hgyrk
rdByeqKLtv25CvgHzHCTwe64R/Ia16bud+9mDA1vweP/RAoShfbqAZ6LUSrZiS2X5yKHY9YlAtwQ
F5XYP74hbEeFp8VPT58bZCg27FcMStAJqOMoFd+vvNUoQgJ3KEgMeWVLl1UFRWdrfbhh9xYCoxM6
e54gyGX8JwqmryE4kVYKXtI7EVO6Ke7O3PtYHJ1PwezbmF7XZuwd5NxY2htdAt4L7hxeLatiJ2Kq
eEYBdfA0YM53MvtA9IhTQIqfS+b1157Dkj30x2LlzeL1ShyVh7FRPfLNspn3jSPvOjsAvqmugsAP
Dc6DCNO9CNGyRLscRF4pmDEH7Et05NG+mmiQ9vQ103biRT5aUPKjQ8yQLyshODzT+mrt2B41dtJ5
4Q8hBA+lwEVXzGF7I11QhzW/2O936wWV16zwB4nTD1Q7P8NCdlKt2ri02NjKp/sVyoZHmNJx7K8d
0EZIH3JHL3BQVCs7y6IQEmQBhivQouMRlmPE+7TSx4JyOkllV2t/bF6u1rhFfnKYe6AKZoD9QwwC
XHwMdWCRxV11W1vbdGkuz8tDEXrY6BGc367UNuf6pGsyYu3JzhhTj7ONdt+j/zw6GKbPV8kxM3DG
4I8OpXXhCFieP4fwV+Mtsgji4Ndi/3534aINX0EVQAjVEkE+xMafr+NSjkdJ1uwNFo+KFZNmE2Ia
6MwGmgbdHvu9Z/b2Ej5vzsfXAmYS1+CUg/40tDtdn0044V866Bjeob/Me9fGNrE07B5BIo4HnL/V
4Ycg/7isZLrv0ABY3zKT9IjRCWsFVyxK4CFjgbxUeQxTaWrZXof2SZb7mE9pP533sCV9+Otcq5ZV
gMGFtu8i53h45ZdFiDqtTJJxmw08C+vkOkTI7MkL+V3wmTikE7vDsU2PJxEWelTKSJqQPCVzFiWF
Vyw98cYpIZhdUUvb7u6HFQxnY9JMBo0StGUkausGqA7K/0Ah6/4dEKOIdcKiAyoNImEptVzs5Lkg
kJmDPMomqCfwJMcXIgYHsruoKRk+ERJ0OIFN5gtonL+fz3lWdxXYx72j5iFe2srqSAnbYmsPBAQ8
/GYrJMJR9+U5kBIRSjyFNRHXqltAX6iwffvhhrreXc44rLwN0gNn4z7vtNdGlv4dcJELmfMiozcS
kJYgXnDFC0yW9o4ZitqgoKPayB5yiYPaW6/AC7HIeJu5xJVN2t6elQRGuFQU58gko6GwuLC0D8Lu
Qds2PMKTS6j+XMtzYCbRIsF27+Lmy/UViI62wKLt8bDZd8ONQaUNvofyAWGJbS11uOIfMsmc9Skp
zfLVrfqt7fHLi73VsWj5N40KsrT+5CDJE01XxAnJloUDoYf0cxBfyrOkoMxB1ofbn1cgqm0WJ1UQ
6vP0LiaFYCoopMk+/fedCxjxyP9Tr+1NmxWKp4KOs7p7GhRT/HZ7c/TDAoKViPyfSMKZITK2FmQy
krki113mPE7m1ofAzovXVqvXx07rrMAZcxRWxuCNYnVaUV0aSzE15oisJZX3MuS5m6DveZohOQop
VWXq+Rs9e1wwvu+G302BYr/1x4Rw6AEsjwPWMQZZ0hilUHlcDi9rMGxNW4jo59AOotxcJO6pUTwL
aDsitRo5RTSd2ZP6xVUMQQPpEdp8Jq+IeE3sk8NOweMx0tqqTPMUPlY/D29Mi5XbzmULwESwehoK
pGi6PW0Rqi5vk1jaibA9vnA7JTohZl+DZfICEokEdfR/i6dukN1IvyZ/UMPqCdErxdYY0BbqgNMC
EzesOK65R8nTtryMbxvaEiTLTfo36C64tyoO/RpKPIeU8YdbCpnOqyI1TA2LERdQ3zG8vOz/XMeF
EhLh+Q8D4ugv21eMLIL56T58kwbHvGP26Jqbe1dQq8KGj/6/jilgJE4tKZzY2rjIaLAUUanawqS9
cTIumo6Vz2Mk5nkt9fAnboYdQwYsbt1HY1+V25s4uB609L/LmuY1M1dsqSTCbxpDM/RThTxzFuWE
rw2TsX0wE2hPrmTht/TS65NxwClWwsqGKn0/r3cV4ToVe30Lut+zfWTGLEoDHy6qC8MqCkbYxiCK
oXC2wKGLIuSLctbWVx4frkMpTi+B0TaCPtlLQuD1GYa4SKWWShOzTOHXB4M+dCmTs0CDP5tzEbbB
gdo8+KmGzugXI0VoPiXuB58FaNjxYC6MRE8b+NRgxVcq3ALjs/0WmQXpL/fxE7Y+eU/bq4mztyR/
Mf6bwLDK7rcj64lSwqDu1G8ypH3L8MRHirthXSDWOTTLcybbyucedpB0ld52Uu8K8cCRu9+ZXzjg
6aaXp4Wic4r6iLmfaGwyu/EKu1U2ILIBs0Z2wadRi53dlMDkdcFYvcBQk+aQnElhe/dp4hmmLhoM
jHW8FVMitfMHDsJlDfbNddfZKG9Ym1dm7c+q5mmxgDJhzZ2X9lzO6s2aDyV32xI6lCkbBiP8CRbe
7FNnWFsiSS+THfx9/UjDF7P2WYOYSmzHvK0B1YLHnT0pTh4WMtjAFu7BbCnR2d600ZPmpbJ6ruPZ
c5/TqhXKxNVWILbZTn9YrdDlbtLOsaE7z/k1SLTLM0TtkQZGbBZnPq8Ex8vBmmetMpujQcJkDccu
4tEyDLYJ3G66fXuTPkhROWFqFaJAzIUUOXlbobYVd845pi6HGloz590jnpWIeGIouGxcGX55+knz
AW4aHSqvrO860fAurJiDWGFHSecKAyCIunZO/cU2JWqBvC5vLhHVsVo2rkZ2mZjzP/LGviBTWPCD
pIFZxnakprT5x31ed8GFc8/AUVCIbXQXQAv2QZucamSZbmnBo8OVphq54VGWWYyhpgKx9dk/PD9H
1kzhjT8P4iB2QrEtMpcvFS5wqDtCLQrWRkwsWexujw3CuwV/i3NrTqchIhYG6py6l4B3Jon2lrfi
Ukxhr71exc6ysrNh9EWXbvoiQqHrAjEkdDD7vkJHG07OlrmMMys0DuRwLPkupsgTjwSgC8vq+lCA
xDZ4/O6tZW4R6bUbY1JmNvUYolYu5sQB9yZDnvXVxWnfIOYCRC2XNN4H8WmpIB9EpGs7Uu6Q67cT
mfAhv90PQvH2NT4bSwdK/bCqDkJhp8ymyLkjg+SaS6zvLCAeCsSCOYZjmWSMSkSdmE6e/U3/21/l
r4t+X71NaRBjNPXA34AVSnbfVnMq5CE5w3O0+eRjntd7WqWaskxUNnyGVCyI4G27UEWZNJuslIJa
V/wunAhPzvhWLjudiuJIAw8loQNaQpVC/IqJ1ofdFrzUwF90idWqmK0EIsORJMc+pg9tzm7EXBW+
2v/wSekZwFNOt34qleU4fUUcOz5ei3uaR7frX2UscFkgeFY20YA9mjEmQigjE3jkhFH4boZ5/9c8
0uzyRX4uYYb2I5WUn+66Fe4EonNDQh5S7awRcGnKntLEeLmh+goer4ScSOx/UqQsFQ97Ka/pPFB7
2NeL8kbARDgoSs8wI1CXDV8/Sf/B9o/moq/5GyrpMXt7wtVcl/Cgr9mTGARBoAEPEqPO+d2qOyMG
7/zoLnDf6RMjcWfGJkRBz7OKkN54rgtDt8clW+1oTuwpytuSh95Q3lax2dpchzePynnv1GIOT+Az
bbwzBRQ4PIcOOV9NfYA5wN6A5cxjoeZbOu3qjqjKrI/Fqqt84za3hRZbjeyFrMDXm5vvOW4Owiq5
6zjx3eOGx3FXF/IPVPpGEEZKUKNOilUZP3i1fDZUhNcf9UpXxmqGd9/pb+L8INcR7UdrQxmz9VWc
aUVP0C/hZnPE4aczW6WNDDVarrV6m2Vyw4d23LMfWe7vXPk+wMXkqYwrwne9Y08UKwAufiTHUvy7
r2qe6QrmjIzcPIsZQwosf1BJMl7SwcekBnDFso6HnVUENAliUEyek13iSQ7YvHhLRg6G1Up3O7GX
hk8nXb/ujb4rj09HVTPfxas4bB2ciQutDSNEZKkmQXgqhkoyLx+1JLInx+IWiMGmtLCz9qlOi8Ot
8X3pcMx+KCoBpmykIzAaHO6HWcGUEYFWJYT8ysAnji4MQwJ8n+vKx2AdR4QfZ9ixn9nooIMWa6mP
duGg6ica3A+lZ+Vc+bFCncDEsG4Gjgp0Vi8Flfu593g9MDe6Qw4GBkfvB2zZ/nHR/BU65XQ2ktrM
mufIuYUaMh/9rZo6UzNeLP1qxyrtGVhpKZP6HYFJFTUNl3gyMsMOB1ayUsdKsUfoe0EKpl1DbJQr
Y1PoD76yh9Pngf6syphhR80HzXQPFyar00RDJZQasbEBu2VAiVojWQ5jwHvRC5aS7TUGrksVw/YS
Z90SwAGAlvPM4Y2csIKqqT1DTt9jbTBRHiHY2T99JQ5OddVUA3jC7C2+Sac2x6kMxuXDg7fQA3GQ
jdl+YUqW0HjKZjSHcieuFDrUhp/sE6JoeDlabopTRtfeHBYz05EqPlfUk4u8LW2ghBVDxZ8QaLlK
NgVVRh5T6QT32S3ADJh6gHSBh2huVR/qIIueyyPXSFm4YGtqPAeWn9tEOZyIkJzBnJHxzumLRuht
EA7ZScRltbe54YrfkapSJbG5sneUiUbnIWrZRm4+am82muQpFn1jvjFPy7QkdLIiiDm8lYKJrysJ
0Iqj3pIK90jWbz7DCqd+3gVu+dt+4I1ulb91w3pkM4e7TyvWP2iWeEA+VDSvpnmN2mRI/T4nmTaW
xk0a74z7U/T8oEwCSCxa8QEWr0QY09t5BPMgtEThltKwiSi8bfWp5idgJaeKxcmN7vpL9jhakRFH
Ej2NB8cDPgCg3ZMsRG6ipgakiJlu+dIkp3RsU/jMt+EYk/Hts7p2nQ3Yk/Mfl/PJCol6ZCIkJJIy
WMbZm4OnpmEKwtSnEB7z2fE86nwksylqcDMTatZmARNjiy4HHK0JgZTuvW1x4vG9HON8M9rThFkK
LaFUJYgs9xkuPjwohg8PDCfRSzWhvM5Esqfh279TJPDBfPxy8DdRC7dk7E72QkRPTiNh8DrLLMVL
fWSuAxl7lZi3tXCbo5zZBXzv4URy1BhAxDdib7vsbs3YAm5BuUssPEm5AuE/6mivFi2+6QqdSiyq
W4+N7NnHq6ZQsOD1U3qHgZiD9I0p3PGOahGOYU7SNzoSkkEuQjhTt773Bh3mC3D15W98qkUQgClO
CAX1gCvwZ4mFmLRxWj1Q9MnKDqf7U6WyNA9v1c8QzJODqDQhwHI5Fq7xZugiRlwb6Pt5vJM6CJiv
b7wozQhHA4mXVCqTrtwBWUIkJZHuEuASCdNZ366n7tK4J3UeL/+1OAMBKwimDJ/BlM3HhPoINlDq
hmFGkbNHAeDYXxao8R9PuI/7j5cHw0OuNNMPM6sCemr+A1E3ZO2xhrscMUGqvEsGYZdSr6IMT4K4
taUh5ovsdXO5Eb/w07HYqpvLzdrD0REW/pZNoGMsCWG2ROhWA1zAcpRW6rHgkhVLV65Z0YWpUNIO
zSZO9XIDP+DTz6GapNCa1CVnuQrwVFGv5uXjzslxlCgU5IflN8tBob02D9l+avfQ5vjsabVzrJ9a
ZEzv7kj+ANXnJ7nkvVzCgPgCBxy+iJLGGgbcm1slf++UAfl0Q+5hxPUMf4niuydH37u295Zg19YW
kQgxpjA1yyfMlmli7oJaD96HoF4bgbWGmV4vZz69Xym8ONajm87kwlIIn1jFRjKjmUV4qtxeGixu
JFBNT3NcQg09zSWZQROUdekdc1lUOtIEFOmdsZebhY1yAJa53b71HE+677jdk4uZY3QPls1GcIG3
Aq7+RXM4p/hpn5deb+jGKjOM5UvWTXqxaRL3f65QhpjquObKnrbZKz0RGGNMcAMawoYdgCKnh3kr
+xWpZiLABn4ljk0lwIC/PFPn1o8kV0cmxBFV744X/QML5Tcl4JXHUIl7wTla4VliEUb3IcIOS0yQ
y5WkF3U1N6c1D/ul6woGJenD9PhzOFhV6dkbqPwvdw9FYf7F1TFRyZsOzADFXdGlU7qm1AUz6Hl/
J6vLsY6NxCVRAacfOBNMYEWrnRiV5Cm1xKYnjRRF/RjKUR5eoZ85lzEhK2X1sHYBJ+sxMX5D9ldO
8KuMPyNSKn6qS9zJGZB+fgVmvfGfoMW4UmrHx4ctQ1lBBJdRnKgdIAoz5CwKNdke2sPREyr6wZ7U
IZQhPqNP6I3G3zTM8os08wBFvHT01HrPbuIFeYZq4uoi+zXTEyy5bD5Xl2lqXur1sgInT9RFzb7h
W8vbKi0UZhtJo8w61+vchqRTHy4WZW6E0CbSPB0NA6crpLU9EJs61KUqH5u0OZzNpoRFJmyTn+Xq
YKrftVD3d2ABMj8e9tt8rZW4WTFkI+bc2d27smm+AFR882bSLADA49/ZphdnFbY4ORlqH0WJbG2d
zYCHdtWUzyKNzR6gKREZkxMe9Ut3z8xJfO/WofF4VX1mHrMb+zUKeQRI+N6Ctr4gSKcPExlAALnQ
RVkqF6HYYw5XcxIHmYkpuazCTHFqd017Gme7l2fTSgeGezTCF3QqZCfclsHfoGZE3u0x9cNsI+Fd
oidqcXnyx6WgVcAuepaXJbikDAv9mJ/u9I/sdxka9C/rHDlYuJ2dQzUv5A7JP60XcUHFB55ikOKo
Hy8Nm7kJFWWo/g7r2qku3EIjFi+2RfKwyEJLgMawJ1v8QRbUTyY9ASAp3W7DAX0nLYhqLMzgqfbj
rF0KNUMU+drQFgY+uLO3W+63iHBK/ccbemcil77/NMsQdHYpe5KejHTlAl6f/Lj2MNEu2JoAvJyQ
N7Ux6F9jWvyKMJoDllUr14wYJVRBiG8rBT9iuhoB87hlKFDyIL/XlM3Lzm00PI/I5eEh4WHG139j
4ZVpxmdw0HhcVhl4hiTHmwEFRxNVTU+MZwCmrEG+CfxhypKS/nGvSsp6wBWevb6uF9HyESwYcmxJ
fO5fJLHoZV/V2qGE7q+K9V++bSzP1/Q3uB0Q13U4qV39XrboRfctVpzhWmEIdXjIZ+fUBI38Cm8x
rlZRzcbaTHfve0b/MySLDI67AD1PG4/yMvldvDZKcih2GaBpI1/BNwF+QxhAUvnZcfLew0hJtRny
HiLwNMS3o8JR4XZBY+hmOcDL2XrgkhnaoN2ub/vUrgLXzkMtgOn6/8rUhyymvPbOgAQD0bbPcYmG
/SPUkVAC9r6FTwD/NBQcqzFwoF5qz0+nJI1veLOVnso3SmzedOQhfZ9JaFLGgkbkZ+7szOdDhm7G
AqLLAIzrWw27OlSz0rSb4uDr7yq/0SzMGfpVmiG1uqCvSTrXA2kgcvwKZ4lG4c9JwxnsXbRfD5EI
bFGwV7YaFTHOdTUXPiNHWlPZKP0DoX74L6glDP6JCEZIwJLif/rXpWh8BUqea7vCBYBbH1ayjGT1
SjKNAeVZ4BL0+dfelhH7OrzID00vCUayARkwKoSPrm+cfyF655/HMJt5EzaPEuNMHZyHiBKv7Vog
kIeNMrWLLVIbbmsRbqv5kH6ZkWPGvJdRaNqfS2bwAWYstSzp4MNEgzIOcBygo5r3BF0XEnawWE9S
25YnxgKB7qPH1uM3LoGDsw7dXrg67khA/he8HhBIEqH4NsyhHUje16WvRpAysNVacFn1k7sZRJEA
Tpt0IKrQjSDF7XeerUbAbLMrDUBBMHhJdEzPFkR0mjn4JWH70/WOhonnJZASKZmC32LWzmdM5PQ+
QweUgHYedig2StSDBbGcunhCD1X7WYXjzLSzEkpKzDYrzbvbfTBliv8z8ILj/JirGhKu/BVXdQLG
4uOwfZkPyfw8qhlE5VylvYu+uoRfJHxLVsYN4ICzblviWg1/9mRohTq8fsR0V6IQNrG/JRDDljh2
I2EERe/kzHv+twn1gKDGOTXh+471brdG8Z2Vo1gXgzMjBDrXMFdxl51QDVsf3LELcKbfUCdC5dgC
NqwsgLxV5+fuUpP2ek5OdZauFntZH6UNii8lr0SGcNcB2WRYxwRzzTequt3MDDnofrXOO+w5U0qw
pH73xtdTggBvN13FnoFshhYmnCvkWh1iMZ6bnZwxAh8k8kb8l6ni3MZqmEEq6gi41ahFFq8LxMJU
e37a+EomEBESLZKnhr5EX7qqRlPA0TlUSBKGVbYpGA2wkwQOHQG5VyFM/vyAUeduLYIlEG9xc0nO
W5HtW6oDw2pEIn+63f1Kc/BPi7TnJVJwWeFjmrEsyGZIVtzvavtvZC/m2XALqZbpyhGpNzqaDsUu
SCr9nms852x8/m5Pn+9zl1TJkOBXxyvkJFofpO5jYqclfV779ZQbF+DzVXWM3BHisUgq0xCoAT/l
gvp77lPSlmwM9D0WWG84NQ/B5s5qkmHb7otOmjMDEL9eqHdYse6wNuiYg2bT/D744k6eUReoi+RT
D389Z2dW6b7fWdSY5ZvyttgiwU0Z7sRglrgeawblDF+jVg0/JNIAlcV+wjYZ5cZ5sArrS/aMEdim
AoCswzmrID5EbggmpG/+ZNmrw4UFvgSzjPQ9v2D5sRBB+X/5x9gOhoYaJqM2w08wiBIJHC3FhyRR
OUeqL2UGZMkn+DX86zOkHD5WITUM9S6VwTB2iig53arzF43YeqPEM2vHQZgfD7feX7/baQ8r4xhB
nOig39OYYozkOYpwpSfar6ABL6KKkIadSbQ3ff33f/6yzzDa7/xZALbTGfQrWHNgMzeW7nShIbiJ
+Aw/LqjAouhKiNhzl1IqckdIbGmaxq3OB0JE9UlvzVYvYVH3S9NCVvZB1W1qR9HrkNCNNdShxf87
2TJ26oKIUMXOabFKaq8r1pdT2OZJetG1DSXu4FXEuBjYyeMOUTqQzp195ENh7B2TWKSf7O7LmKNH
98xJUOBCoY0UTrGdUFXoayQRPixWSDdedyBvaW8kTNApJ1qq/13kUvbNCeBVtvq4hGAY0vBRJekM
iDKV9MRDsGM0tOPVefxJ+mzLqv9+mPWcOTjcJ1cb3qvNLbJ1bZh0/ULOeI4J3ysBGlCz2AxbZ/OY
DEvCuwejZagG9OMyQeou1eLLUU1FB4emWHw/z9pJ6zfryT3srnBS0nEBBgkFl1vg8GIVjxTfnw1c
F0tcNaxyIYhe8lmvea6g8yMbsz9SOZhKCA7qAXZjclop/qWzSq99kB1TBOr4TkIqilEoksoUCHJ4
DPMCKuCRg9wta/CoqLS2g/KczkALIbRZlunjD6DUGyF0P8avhhM8YacZae81B/29LqdIk/0AhjNw
ZzqSnqbgkm3MhwGqzR6PnyNyViqobJWl8cS680NyGMEmSwR/AkRBhT07lvHkr1yqxlFNuUpO+yMt
NGMmGWH3jYyZzlzby29WhlT5JQ4VQkEwDF+8PnUBlqeea+6A7xPAQSMrJ/g4p6mTwVzAE/i7y3Y2
i6Inqx65EfvNXb/Rd7MVshUMceSoyfE1x2mH6X4ZhhDCU04LLA3BkinX5zRXHGT/fIfbdJXYnxKQ
jrqIH+UeeVyVK37uDBY0tklmM986E2oygKbFo5RXE/npSd5GnhkqDNg/46MgyNoD/74SKvS6lwWu
4xxf8NEiAA29YuISXNBDkW1BjlQwm+Qw56sJXksh7oayAm5Zp/Oz69bzhpTImnpQmycWa3MXf+pI
3ZIEc6kIDYixlg93cp5sUzzfceh48h1vYVWMCEx2sdL3bEGB5Hu+ew3o/XDRUc/fguS8MLk/TslM
ICkP+mLcXLycSACGtgjBA31JOKjOowyjeapxRF2hm8IJ9i5BW9vvqtAve7tMytGQNjm5JIBd8WTd
RcD1xlshJwGBYoteKzxEIFelx056X6rl/7+gcKfJa4RYRmdZ0AYjT4q5J7CUPLrADQnkHQ5tErty
zppDU7gycGd/vjWIM2wyDrkSJnvVlcF8RIdZqcNl8VnUbePrSi26+Fsj6rFO/ECjjlUMoa2Aq55U
GphtxkflluH5oYjREi6ldacD/6dpF1fmBK8bMHV5ynPKFm3lZd0PeLGQtYVHW8buwzRjbSR5JLLi
4GLtczB822zVZ1YXPuwFEr4B01441kJjOwnCXA263Akvs16A7r4rVY7CfQ1Wf+bXUqvH9eMwVVqq
DXDkeMpq80AU0viOGPNWCCiZxDLJZq8596EeYe9gGWEiTlv0929VqMCJu4D9PTjD+kor+r2aVTOe
91axz7pH/okAyn+axLjTfB7jUBuVjpqURYcZovnicBXhRagTJALFnISW/tT3MYtSPgT7294xzDr7
/mFHLYWfEHUNyc/4E8zptb5jTL+RVa9Z1hwjcmJRkMzmh40IZWhhS0oy0BLhPaAL7NnpPXxjILBm
qhqZVG7h+LYLnFlyb/eRvDgAYft8xOXXK/gms4FRQ08e5Mz5oqlj5kXHCVXEQNFan8aOZOh/OChy
yxod4rXfcN/jZVSO2dkuVgPW6sECSlQ6UQjqVzpWFeH/My/aNnxoD1vPtyWjxz7CW+Ofa4t/yS2X
t6jRAZ9ybH/TDQNHP4Bv1Smlj1lg5YYrHpCyCxB7q1w91Rfyzl7Qb4ZLEZoMRVSPuNOG+1212FlJ
0lO1tOxa2qP+L+Ycz+0ckoWjRHA6rlatOHXy4+tdMA1cFwEl7ecUiHgd7WuWmBR6MAR5kZ+HccT+
4nNqEw5W/SOVuPBOnMjWqzmt3UpSljhDI0mkqIm1m6Rtsg4TtPXAAfFG270KWSW8KaXeNW9FQ8zC
O1QkvFO0BZklVxh5rV+vpmFxhsznZ1rvuyHBYMEJ7QM2sTvQWXzwaP7hRq5I0eMgaszj1NqUXpDd
tTuMeVCy4jSbM4rVmiO7UTUfemVQ79HYr5zChihhmxzdMGcVDP7xlgQ+D4hAwLNknX51YILlKC6Q
FOuBdi+jPHQqP3DUbb8D7JCJ8B/YdFTjNizBHOe0nR1K7OAfBBqc0CFCy5zJi/FoW6h7LxPGTWFe
y9SKnDCU345CUDCCkrh1OwHkahSJj9TRQJH33Khndvn9PezH5d5Dk6Sq3hnMiYhha/JCpungFyuR
KLBoTYH4iUacpwd/9/i40T2glw69XZYKx5w1LbzhQtRZWuzvl0iFvAgVO0ExbtzI0wmR3v9YYp8p
2oz+09TmuJYLGydegVXzkBGpL61VilNahZWF2r/bKqIINSXM8y+pmBVkgydlYLXt4dZkbGMtfevC
6y6YqdMgFNgOgsXwe6NLG2sAxhSB8DAJXvlPUgcl5Z5aAnkEKeLYvv4vFRzcQoa/KEM0OT+ku6Q9
2l+F7K6xOxCbreYp3g48V+paRahMsDRv42eG+mbTt34Sp1khIVmnXtKlDkEllS/atzedrVSILlZu
UYSTNnRhoinLo5Ga4JvAJ5fYF4pybzZSD2WVCabufGbac5VK6p7QgIPDBuINfjlR/jusTxNtyJkz
JMbMNiDL3pO9XeRb+i25IoFic0Iar0zdiSKzDOi0l+vrG8VOjW/W4QEI4o1rtxbeMzJOr8+htnIc
adTdPoaBAF/rGPy5drcfG9Aza5haVNFNFCdw/OULr1i3YyWv3Wg1iJ2nX3L1gQlqfJ/eK+kli0/e
YFBk4Qna6PbcMvC5f/RfQkYyCrkrhgCJOZ1HQBr+old01kWpPdnffdvSa8p+7OEMhCGU2OtmZKVh
BExyNREyj+aVpl5xUE6PD9lfdR5gH3MJ7f4o0nyKZdq3zvsuDEfUQ9nAL/qTKWm0gO3kPU3RIQLu
dMJjtdBMt0HQQxDkQ7kxrws+Kp9wLd5Cgo80DKwu0+q9ac6PRtvFYs+4kTS1YUjguOB0O/CZxgmG
b2vcL3ogn7kAsNpGBsoY0fv8NMWsMz4Lg/dB+mzMKEvQytkVVl6JfvVuhCjmTonTomkTu3dE2NTP
mlrfRVC531SKzSHZjidpn2IEOS9J+ySGWjG+Z9ojWLaNZtgWP89CiVHJIK4RlGt93ZAdblFVNMve
l97J2P/LQ4x1gAMahhzD3GZfNDM+4ymwk+7CE86SLCjuKH/QGv2hJYV81w3SLMNRlipvgJenIdYg
oZExqfEkl8JcuceIHAO2LhErWg7keK2egxKwMVaa4ALrorOPqqhlLWtz8U+IbdZQCLTRm6p3M4a0
Q7apcXZxEOxoE3Vy7wOA85kjKtHNpInbUKkPBzqIj+zfMust6SGlwgWeJ2DEYayWmKjh+k++6neL
yfbLna62y6gX6f49dlsxOcyYuqfYWhda+6keNDj+LrYnBgyjA0e8TX9OsFSw+PVxvw5jcECdeO+p
eaQYv6fWfxx4H9mIboQEDzATWko9qeqv/CDQxJcj6BNCgpomhf07h60CtyoVTy4/BIv8HFmb7uxv
tzsh5vfTsUgd0RM63yyNDRj0dxET/yyFIwRhy93vwNkD5UndB2adYjjbM+NLwdvts2UwTpcZUYx5
LZCeSXPXjs9EozaZ6D0uWiqzHHIalSsarKSCwzsmfnnkM0QzwM+mBUF/J6RUsHoYrelsqI3nfYlE
7XA8NBzGynGxNbnKVHyx6QUMNvkmJmdY5Sf8RsPNJfT/qEQE9CMaoNat+Oz7tW8BJFcqp8s4hWa4
8MM4Ch5k3nFkFWPCo7LjrKD7NbuQRnebC3MREOe35U9rlc9U3ZHZ052iDLzGXNB+QjF+eLE0lxUI
BHi0u73ibabJxNGPtoNQLIgmJLkYhSV2IKvfsZUI2FNyAI97w1e/R7+9DDS4+mEJLvCw7b44JNBy
Lw6HInpoQGGQbXREwW81oJRWOSpBpTcMYXzCqt4qWQDQWIHqkI2j0ApkpDpHrf9E+/JtvFamQP0F
jLQVo8pZLZFygr6zbbq/4gQWteCOV/dCIrIRFgel0vXgaZ0VFC7Tl5GMJSfNamDjxr9W2uJhPycR
viiI6JW/2d1ExoFl891VqT+1O9eayshrujS/aYQ/EkOCi31ssOIlh1x22zzW+x+yB3EDtn3HasNv
CNG4kQJOC21i5LROXS1hTU55GFVsiIKVLu0quOww0mEFx9Ae7E+ywZNEz+qtbFb1q9Cin7Iq6ErB
wYVDbLLar+MwkuwBvpisUs/d3FazQ7TmEsOv2YIdvaTSox3QCbUEoBWa3VNhkXL3k/GcmxGJgQhC
aw/jklZZJGK2lSXHeLNJjNkgMEWaDTmPTpCAZZCyfJOuCe8X8NbsKWhuvrOZQo7sp2JqweoevD4Y
Wm/7yHv8x7pKgmKgRDAO8VjIw2I2O4h2gXxhHPRgQ3YT9xN8VASRPegZNCSp8szRG3GGgPvajDmz
RJzOQPbQRMn//TwpMs00IyJP+N5HKfcZE1aYt2OK49jSsKhV+nBrUF0XMXBwC5QLqNgpdNYJjiqB
r/Y3pB4HY6LZ+rDqSvDZMRinzFLHkO+l+HVSKa7gK1vsIyMHph45QPDGFnIOfQpUQCHobuqVvEgM
xjipGfsgxL9ZbJrgh3/a3aKogmXHwEvkguxzJy8HRiyv2/FDA9n31YyrsOMVfarwnffrNSkfez80
NANiamtq2zdNVTMMEll0iiWyUuFnD2gHKyPJKtBm3lVLttW/QJUTlSGCk+15/94oAedYlxppJ5mf
0149OChSsKf6sTdJX6KHkJuiyLCVfFil2NgzF90Q9JY9Yq3onaA2BDpPQy3IKTMEKXV4ge/KVOVf
mf7Ijb49F3+evyiT8QIpLeCUKXmVzHYCpUmCktmqGGYOHVtO4hSr0mphcVyhLM2NsCaiO5Py4dab
XMPVTqw77spQ+QafuZvS3/0IoNnafomzPRJjUa5dGbEPm0RTtU2UYyY3ga8Maes1iSFKGari2l19
s3TXSEweNZZ/WMvkv3L7x+XwItZVBhlxkhnq6XxqyDCxH1VWY/RCmZElvNsLR1jW9DTpBVBtrs9j
qpQSiEji6+7pt3NViSAYp1raAD5Awh6+LonyZMpZiiVNldXKLSsVATkPYJUJkgZO009OFYKJhfsz
rLMwAAP8DStRL7qSiwJhvIfSYPtZeBc2eBR4iQh2d6lVd0Qy9mmmOytce1HYKiB7Bdw+WiTnmm54
3+C/PjlVFSW2gObHkFyvqJwxdx8jlJ5ng0G8KBy3oJw//RCWOmOCf29t6/844ZObc6W3ir9AERyH
R14YNycOFMIvM0GR3PyqT3PXftLCU6aBrOM7jfVYgC5AJP+ex1DThl7lWhx+dQM9Hmusqv4febr6
op1Gc1dpJaJdqV7YOYZ4ZHZvYfP2xsXLWYwdhbliO8H2MZ/5aPf7qWkXzwdU5zVcyHPV7aMajnJF
ci4DrNyw086fdaenP8hY0HSLb9HJEjBuTBhMSnrJeNbzC3a5yzS3tS4/dH+e8v5AHuR/RFpiEI71
Mk4YiqXUMhzw+kb+U934JbV5dplPTIshdlJwgCQRPRXlfp++W6pIJgEiXIoG4Kn1WoT6FgpwxUDA
7QAXKSluB/cqvYUC8ZSiO3tdCMIgu6H7hlQ0cSHzBt9ShuA7w0ullWuQipqFSA2YAquCXDRHZBcw
7LxwCgbpt7/d4zvc26750OrzhaQGVCP5IzhJfw2iH8aA5Ub4aQXvOk9337wIPRck0piOKFbkXSyW
8P+rryGa63yHxsCn9irgaz5xcqrU3E2JkbD5OMwGr4RRkpsXBhKfwFK3uCQ1NB6nRM2I29tfQ0t0
dMJSSsFnvrFDNz1XPD0KfmApB6Z9HG1FHB8UpExEeZQhLCoQ5+37cKlu05T89LJoo6BHLhJNGPws
NqGCg9t8HVf1GCl67Qkltyipt85WoxNyqLooVL/9/ZQU+pRLXg8+cJRNGerCO7A3a8L/JrhykKbR
Z8SmYw8b+Ve6SeXXD5Bc2xU6znkV60pp1ors3AnRysIpinSO7lJq12oTP/mZCjxoepJX/tzln2W1
xXOuWSTOBiDpOpymNqKiwp56NY2X74s+RS9OI0xrl8Z1kyb6tZ+le3JxVSVP4oLygKiXzu1Y1HIJ
9BlriMHxWzUmg9taaxSClZeLu4jEBF7OT1jbeTsbKfkdpCPUZW2HMQu1qhXuEbkgPpaQWjeYZr7i
hpwalGTT6Cvmeuq8nUIfJvT5Wgg9+Tw9leT0w5h5q1FVgPN998OpQILmjG4sow6YGwzCWt6aFLQI
HWclrUXBeWgq2iIPbDc9bySaQJk88rz+8O6qKwZM58wTkCZa1bemoubxT2xJee4IiMu5pHtEOjul
f3Ivyq82EBn+yckm413p87iGg7IkGXP9pIdIs7OgFibmzHNNuh0fz4X7OhrTtIeKYMGlroZrITz0
CKfCkyw6I10AfhzjEZnC0PorBKUs6NFAqfLwsIqtIZS/9AdbXgMVi0y5pTjb+NIFY/JkPPNcnSNK
7B2MaYUe6T/TMLpFseDJiM17SXuG4g9epHq9hnvvdrnCj9ElxtPWI2x30TTdEYBD1IdeDmihqsAH
cnQ0uZ0qUcRtE53pkHGEoBb+zs1pGpedTONBgLvUlMR4ECZO2XCtsDgxuE5uFllVGSgXHP2D/H97
XQjbtmPYUgRihmzgZakKl+OrDRM5UgjWzbjErd5xtjQawPp7F1weswStui7m5tO1qyiu8T1Hlxm/
zTkfPmdBpIMAZvfs6+3vg4y2WXuw7c/lahmaF+Cu5jMbxXnHvy6ZEkj3Ch6bERtaMCZoh/z2aHK1
7PGqfd0mixoHGZhYyl3OOfTbcbmK9GNuLHMGWCdVnQwPtywIyRhalmq5wwP442QnLM7TZkQJKETM
4yFj/NHrTFxd82zU2r3AsHtpFZxwQx2nqp+s9cVt3W8UmDql8aEq1Pi+cqMP3fn82HV+uSMlq5No
59hmzUJTqVn3hYpE6RZGZY9Z4anof2pMA+rKZIhsrco/p1bpMhH1enVVvI2CeNYMhlyEKlc82UKe
4+qW/z6eHo53mUGmCeSs7ynzygJPM7QJ+cjbssivW59sq+P8UzouEs/0VG/+0VGXqhu5gaY47I7P
9mF0gzwjES1sw4vXyjSSRJc9AL1yUFX2KEKzFrGs10FL1uTXPhFd6mQjPpOy07gwhdCK2Ttswjzg
3f+uBlTKSbYmlsyXubyvUQGYSLpankuoGVFDrEcCFwfBnNDOL4tPBkvYnXCOL5doZun5hzDc1gOO
phU1a1B++K52FFUSgww/XXJeTq7SsExucT3rg0ni64hHzeNL4yrfoQsWWllb1rPbwGtAB6FqD/Y7
1JgXeALpRlNHS8S5CG+WdHN1abq0wJppMrYmgAobn6vLEhF1fJ92GgQjrQzt63oy3JeBVEuOSfzG
VH34w8HSdtlVwe4n6lAt0doCUxKoS81A4ePVgILXZzF1aO9v+ilpgN9x3bi4oVUhByTKBqyd4XVs
jkiFPHi7EnEpKLj9Ynk9i37h1NE0JsPIzmiZl/q56yCUWYx8CWVuGoWeAscDe6OAvyXTXIF2x071
jl/cRURrw6VJF0gj2wGpUevvYN/RrRd2N48ia3OL1dD3nOpRXcw5kyiAmHyOLnP9jQmOwKl3xFTS
wadVRACm4YJ2XP/8Ki5tFFT4OiwH4TvugyZLOBKgtT+R66091UJr9Xv5blqX5xnFw5xOX7Upp5UD
FMqirTSykje4omLB60B3njhrUGnJqY/7yE26E/WjWrQIBL8Doy3r2Jcc/DvaFcm8guWzU3lsEtSG
D9YasryKndQMzTqVsbXErEoNzEDHK9/1HoGnVUvrAm37S/F+Zk0GbJoGQETPIF5vXu24+TfWTbrX
TZgR2bodUnZcWltF2eHCHY+yWan40np3L8RsMJkF7IuhDQk/dyTZkkPssgU+HoQP99hwVYzIvS7J
u9toyx3++KH/YPq7Gjdm7opg+vtJyVLtgvN3qnFak2LKu3KoQCrpKZ06XMx8i7jQzF5jcVd72xgS
SVLPIXEPZLyxbDm7y5AGB3rSYWwi9/o7GCDRfF9sNMkvfF3Zw2Eoyf+sdXI+EuLxFvsJu+EQeFwU
eYeY2xLPG/QpEMhCOjZwP5s+Y6sO891luT2bGFw0IWXBWO78PCkVjZcG3lW9UzMWVQSyeDjjKlmb
LMu+/Hbfo5PIo5o0ByB9QxK4JayApQIxPI76ec536eXFgugmFvMbm2IBcElwpf+loSuRvZEpECfM
MvQr2JQzId3PX0PFo8exhBqZO3/x8CJR9Qk4Ry8pbtoPSUTPC5OrHimnFBJ1w27yMl4WhI/+1ujR
2YsXQhmhl/Y0v/bOUPQ6DIRMzSgM004ZN3g/jQnBrwljDaSkKVsPsZRoOVbL2UPreUm5JwhAKtm4
h8qN2zfUbr3lO+voGA5JCu9XT02CfEo/PZyIBSrSnmX1jzmarxHh4/iPFJwW5qnb/SgdJ+GrTNHA
KYvIk1xbUYhypiSpDtfzsQtLGHtChh7eeDl5DS7XTh3iLcJpOAQNO360wEexH7X+OImfb20zQ8l1
PqlrDjCh4TO61jaeZpG6FlqrzssR1Dyi0wbRm4pgmgtQdliZ35U8GfaJJYJSotfRrmab2FBkCaTX
bOwg+ELaH1BOvIwEMmqVAJj+NcOTAzW9QXsR0hUVUiDeb5xdTa5VokHI1G42X0f51WY8+ve1zBRJ
2i+G0t4zmLvlJabBp4y4gssCrx0OT92qwq9SVUKex5eTAUvFBbqKAq/zXSuBvKl3mo7WMz1H978R
4u8pGqvfD/Mv/woB6g9XwfvpreI2RROlyMRWyIDzaIpvErikAFPnxgOL/FMx34sh9gOMTAm0OAy3
c7W1K9HX/5XMnyJbnG84RHNaWMlPsuIytpqU6pEDxEkschC6hawox+cvmWaeJ4oSK6qQ/i/y8NS/
nXoSUMbYB8/HKaFKQyAjD7VcahOK4K7bbmO7NvOLl3lqimcJ1AZXuw7LNQ2TILPtH5Oba+xMa80v
QgueV4fz9EdCDDGoFBPx+is1rph9e+M4MkMGUjhNxyyNrh9lOtTEgy0XEiZ00zG9hrFCGvWZpYO6
IJofO4i81UXWbSmwdCjQjctXuUIB4UrXI1CHZ7rLDw7XEEcS6NffVNU7UY86gIfd00Jhn3SEE38M
6xhvcjBHh3eukeRrqcDp45p15DgmbLWhKUQouIJgQkbFKClktP12PYPI7WBnNE9pz7EDNHpZ1UTK
wSweJ0ys1n32g8PMla/QGDaD63g03G2kPg1SZLzKxHhM+p9OUbcMuF67NmiWtl+qm1jf9LQQiIc5
79ZUXEDoTJpXBFFBQH2WJ8yLXfv0jaMyPwf37qkrhzXJ/px1hIdNpHYlTlBpo/IbYPJ7CldOIfsr
CidraNg6CrWDWIN9yPZ1ISm6F2X1F3BriziJ2KVe6QolRqmpOuZdrtSbkcQ/UJw3K47u8+YSve2e
XqyEacbcQP9wwweSicVip4y7dxpUoA/TU2z9SC/ezdRUkbAJXZKC44x4mht5/N1hvda8ZZXs0A64
WF2WMZuZGS0Ef4ooC96ctUdWVT/bTmqayssPWs8elN0XsXUt07rH5sFPmyhgDb1cyF2XcrKw0lEn
A5lwdJtqRa3OhOy8S9SQmqxPJnKnW1Z3KbvCmihN7zFYZ9nCPD3Iwjjot1M7YxJEcxjqbWzbLGOS
tjgUja6vHl/3zCZ/A4ViWgk6gn66vf7Ic9fvqzXKWaIb4pZyjcGHq6J/Vhm2r7ePyDzJAKP+fnm3
f0KzNMqjVwQs45XISxLzOUF8/BOaMkpQM6lG2LPGF+HTEgZGhYt2Fu0gaG//niSE0cYlR6uoz+uH
Pj/2NWj67MYdiwKbPKQMTISyKyvntokKNU+nclqMtcN2BWlJ+S/+lauuhQ6UF9HVkb9kMCBd3O2J
hHFUdgrkgbxiBA9Pdub5n4Q45qhmsZ308DCDlx24eHpe2fRQKr0qWZjf2dr0fkiFA0Svsw2GQpaS
3jDZ0uHoKMq0Lb5xvAbqhLf1QFe9DqOVBPCyzyPQjk/o3ErF6KNCWuFDNitiuW2o8RyJF59UuVSg
Bg/sxcG8C901Uy6Om/S0gcs65DHqKNKTCjJz5+fKGUnuIrwiAQJqGCTphVlQtWzIPJiouxsDo5Pa
dhhfgwcPEpyVCmdYYDs2gIRuBlyyJrxhrPLfmNGE8dVbQlL7ON23Soj7/wW2QLokGg4IEnNrLY1y
xhpN76Gv6RrZihzw+/zt6c3DHYV3CoePeU/fibmIyOR+3HuhfbFWZL4ngJKB0T/uyhkGN5FwCIsV
OwytnNC/+yU2F2h8eFq3QDWlGTJG1xkBq6bshw9YS3stS3e+JJ/7ntPdpExsx8zGB8qNi2QlD/N3
tZyrmbW/HfrVKW6PCK5wwhcVyrX4iop/tPp1cb6iz5+4nL2/j36IlCrSPmjzz51wgJtVt2y4TKut
MbdVpoNK5L5J/X6Op21bVV85QKJsTkHs/VNEQc7c8hf+YmgkCG6yxSlSPIui98T5ma1yi9D3In3y
rnflUlZBFVE6ooyaySPlvbdFxPvzHNxpIXjNcHf7PJ8Uc82iw1Td4cJmpYGsaOs4SntmMv+2Pt/x
uWygzocAiypTe+M74Xlbz9cOHtwbDa6V7FCrpIP830Y8/Js46HEDmkisFxTmOzSxHCtQq9gvG/Fh
tL35G2TAx0jQ36VVT98gAisXjlwiGNqOSowDjGiXHFuctKJejTO2AFza5CdW7e5PHSttFisyD6Ka
uoMin6CD1brrmWzDTz7uzai3VeXY+G0+Oj98e+chUoiSd+70fBxU+FpHG/G8HZ+N+CEug7JDT4CW
MLheCfKEAFQuoNLJsfql0ltmITUOhmB/VVsEzhuh0c5zzc4Pk+s2T22e+EpeUCqCdAbSINQsRQVk
DLk5ThTzVjFuSrqU1cFlbfD5Gwx3rEJLjlvGK7Tp1+k0Mj2C4s88We7gMvavFoRX3yjK4MTE4kq0
W7W+SAaFLRyqxNOKpEof6QztLwWX7aeJiuLvhaZuSBH7hjbsCBStSQqwxmaV0flVyqxWbzE/2KIB
UMHhVVaMjknhiIc4mCDJ5oMTXT15JPaX7O+Y19saWt0X/q86edtsc/hDYL4BZNC++L9S6aqQLiu6
XUnBPhXXKfl5vS2zEnFbRBuh0eM+LZ0U6C+Ko7Ilwtw/JNuZgx5JpA5IIsMYmP2b1Q/FTiiKeUp4
PbTJ5Wzgo+O7o7cFYjyO5Zf/mnJXZO5rwW3De2E+LFx2EOYZAocim6JZILGekK7JzaEdU2S6lA3T
qkwiys/V/AndGkJWsp5kHMqOpTfnmnxNKcoZt+mi3yyBTpEgmd2qrwLn+paWxu/8GZduxjtCWJnC
hGSVr7B/SINwu0LhGol61SR9gSf+4LN2tnYGrxEd2Dqz5UfW6IXzDW5C/fRficcCWVgzQ6BHTJzU
+wCYiHN2FhgRfudEB2eSk1pszjWMJUMVh9CCtiN2kDDe1JejvaSJbc/PjMRsuKgHtkQWGC8aqXyE
jV3Zmnelxu8LNgYQUo7i7YEfpGA5hL2qPZUo+lMQR3qYAh8c/uf+RF7bfweRDhCIxLeT1m1j3Qi1
W1Su3tP6jLGzPE6iXtiabfY1hEBUsZRq6MpBee+5r9if7hugiW3VxORVIGwERPlTmXFsSsUAh6gJ
j4n2U6ounMgFDEkYNkxzFqO+TY12r+wVdh0rlSsHy7ZLp8zSeHlzxK9TTnCElHohWbUybAhE2EVb
GAtAdNu6nXq0tWxlRfC4NllfLmK3P2VsC31Md3XzBNgNV6km8UT9cuWA4RMSWJwLgcCnXj1osQZb
wfH2iPnh3bNxr+gfPFWu0XprfpjT92SEStRfJw0+zB7QNVsYpdmHWS4U+k7Bn/AYVUspjIioIJ68
vBnwnAN4ESxXdGkX0/Ux+BtSNu7vYglfR+NbaI8bP++n8zF644a6OBJoHv8NKZYNqMbSZ/6H3Pqo
E4kvv5Faw2Sb/4SM87aKoR2zEvacYrmJVN38Wj77I3CY7gkA98P2vSVRRrdWDPHtwij6tLVXc1zP
eVmlsmg0xzlMnltWAZCr30SNewa68FZEIebEsJwDPCCAsapr8dtEy1ZoXDk6oA0p1K1ig4Z3zIIC
Nqj2rUnHyB0rkiTEfFoaqqgaY9h24IwP5l6lat+hCzvzi/CAtPnySL9riylmzqBCObP3yLvERbKE
36UjZ3Lb0dnBCeY9v33sBt6Pp6s4EPYHmxffLhNuRvNrMW/Y+rAiwa9sw8vmY6zluQ1/Zv+UqHou
i8qNZjYDAHlpcybLPHLE6ft2l0Ma6jaoG7S7mbTRGAI0dW/82U/E1811Iq9e9xDau5jKvW8SmyNL
XuyHho9YOytwhsqAHP1aFlYmmYBGA0L7mmMvCw0vbTJiJgmfmJDZvkPzp7SZ3DW1gbwAoohe8iJp
Saps1SS2WqDzTdKf3fOJHi95KVSQLPXFFHNjoafn2vrC9pud4PVVJze2a+6ZDT+cjpy210fo9ntG
92OgPqxHaM6NpkHYhFFwpmqRVFyN45pdG7rD26+YARK/NugzmqqJCZlG3q217G69tdjQA9vJR8mg
pX871+c1gZnPl1Cb30LlrPbATSj96lCL7bwdVfjCHKC0a5+yMRu7zqmsMUipE+8JkEor8eB45CP3
9Btg1mhs8klwJ7GLx/KRvjfPqp3R/Mj/+wwoweXUsPc3NsK2qM+fpEYS6g3gfWImmt7PIZsm9Knp
VpTNj6O7O0CejBD0cm8k7xLFcJbc9MYGm3XE6com0NCfotp88HX7cXmjodEl9Kuwcty299o0YoD8
5UXWbqXvws/7y8vh0mKQPXYpzyimF/3grL9zRtjqErjyNBqAAQ17z7NEnDwJBZu8fs10hVJQe8m6
aDNc72t/ZM31Doq+YuwNSkXtjoMJj9Ov/pGDwUejiIMbCnpv1KyO1vY11vgvnId4gjuGub2nRg+q
cC9t19e5GfYFT4yRy/bHkN0ngiSTu9fGG0KigdRk7QsNaWDiPNTXHZJqSBRPGID/bYcv73+Qy7Qg
jRSFa+QAuhIJ0ChQfBNs2JFzoZchynLWxZMIqetCLO8DbmCJeESZFBr4AdBh/bCiadUVO+J7e26R
8kHnHIcZGfVPrtZyGf+H8v0vTn/1iwecoCimFBkdmr7HUZUmvmHjUVqGDTUaLQU48IFtLtT299tR
exhHYgry3XapvwLUQdW7/L/N7UaPTsGbSR0p9CTxTqLqZrHLiD7En0A3G11Li1IzNBTDVru8rGKa
9b6P1EqoAkXTq9mOgYBVJNi19cbE7yxEzjhZJHj5igtHLzvfjePdQr/8B+327R8g4zBDs5sSaSwc
cpCzQlvactHPAO3KK53+wiy5WJM9N7tBsuHw/f1iBRd14LyGH7VAJ2dqvvh4NcasxGyZi/ehReFU
oQmFjWaiyxv2noE8ofccio4XdnuA2zfHbvAbtEV6cYjZ9QmSVMjWSnrXnwwkgm9r7CVqcDsm2LeG
yImx/HOdCg41xnuaJ7Rd+T4Dlo2XGgNcY+4Mf+NtVO3G9lDEzUBP5xTBqi5cjgGGB/oTsnrj59D1
s78d7c7OJLDsX9mNQki41yuWLICCsxe749f2QSXr4VrefSJS1XT45qc0d8F1y2ANvDmbt+BrhmEB
J5E77arkZ5UximValJe1/F2ScDFaSd/92L3MX5gfQyZGJTj38dXeZyezYG+jDA+Da7a2P3U3eZqP
S6NPm2s10CaZlPmH9W4vmLXtlaJh9cZjb99cneBuqsWx/qx9/WljJVCWmzXWOIM9ZdbNgzeOk3Pw
1eSi4bO5X4Ov4NscO3BMmjRmNmI1GtI/dzDIOcXnS7HMjMCeCjyo0bOzt494Tx6m16t/UKXOdgPB
/rR1SPoTNUMomU9d8kHpZNMctGP2WRGEM7fjtDJBunHyUnQi937S1Yr3NXoO6kt+A8TJXRbFEAQR
kOwV35IUNx8XuwJDA6YxOrHt+YUaPVDT5fDh254u7fD6etpUPZ7If8JfXfPHwBcEEKJjjOYPnANI
d5+gyCcOFKWbL+h1Jip/sA9Wu6tGpRj80q60xi8F38P9fA0Xo1dFPwKE59S1pkPKzbiHbaglMTRZ
d1as4Hv9A7yMTPrkjWZRsMgewPO+Pxm8ppK1nEPM4zCKN1HuH1Wh7p8eNUwtHGcsQzLQivjH/CMD
iP/idylWGSCgjj3md7TNq3eV7ZiV/lnEdIzAOPpbdn5Z80JWeXRuRtZp+81sNZzOHyaokkRrJwpv
4/oMbS9vI2Xzlg/ZDGrI2pbSVPjWbgADmRjSqRo25fxqi/WaAcLFGU1+0gK6566jnWUQlRdR7oFY
v1aidKEvSzkZvlsr1pNURkd+0O5f2RT9zezuWmRrVb1pEG74cPc3HKxiaF3ZZ4IRWTK8Z5bK20YV
m05BcZe9/IMv1zcK7BLqY6AQCymrBqkeE52m/eynoIfzu+aLcFiQl37AOHsPcvL07fLUjmFPZfht
26QN9Y2/dwsDpsJSQna12ZojKZEOo6SQWptqlFC7FnnGEKeWLt1UTPzA8Umn0DBWYYyspwnhri1l
h3CVzjTM2geeqlXbdVj35avj6GybSCCQtTYz+5k6UPmbuvzD7Oypu63a1YQrYrN4eKFTV7bdAKci
d4AgKWQDA85HUD2/e3aqLlZw/BPuLT6Cl0CDZK3gpcRO11zkDiZ1uq3CjOHhEOGhoGR6lrj8uW2Q
Nx7BxMFNMiSKSpp42n/wV7FjHyW7Dd+iT+l2658TBz2Hg+UpMZrPo6dqrkLKFB5+IZxxQkXxp+Ae
V6Nb4dw4hYlyfIfz9gYpQq0a5Pt1D+2p2AM8H8zJfCofHVZByRKH+eLXwFX175BqyFcThuMJdgnH
mwHXb+1a969eiwMVrU9Wudm3tJ7zGdr8cTs9t/ZEtGTzQav8Vsc1EDuZpwmwVYiOcRwQ/1XThPr7
BD8grC4SIH8nfKTB4qZrkDXwoh4+c+uTe1JNXX1ZPca5wk5+34CKbAsdFDzOyyIQ5dgQ5wwRQ3k/
nJNx9lKHzUJzk6sKy595HYmIrBeSmxQfHOaFKlgHGscLke87FbBALn4GurhJVYyRXY5DllcqI//R
KdRB5FHv+qvu0sm2Ram3/FZMMC9afPCzfiAInpopm192k9JGxOyn+VkYN1PT8156HIHPOjRbjzBT
0QNzWnTDutwhDG4LVpnld9/d//NS115Ok7zvBQ15Cs1b3tPGF617u7dLupNVsgjMUBU3LRum9Spx
dMVcU0CG5heXptGYC93yO7zFnp16mOtIGur1wmfcidbru7ddE0fQ2J0czpQFKLmCmOIXIh/OHVg1
XJ1LsOKu2x9gDTOX59hMEwHrHPUGxk9j+1FlyvkAnfDRsYaL9x5QUhbO/YQIttSocDRWD6ryauZu
lB6MaXjbESYdzhF6v46oG++/Fh80VLLnSfEMY9FutxH/F33dYHExQpxVRTUGdKPF60UJ8NESJnUC
0IdDyguQbIPiaXokAj1jg+azJ58+o2OEJ4yXvCG/J1KWSJt2m83HDv489RoYGZ6rB7pC9diT1nOT
lYdeDjdvrUyn7Aw8HGM+B81By8m1tPBb0vuw+l/CdWWAZDbuTFy/lakttSxflX64tMv1BLZEleWe
olcD/rbTyOJaeIK/0rzIGmml/o0DQIcedMhlIwDpeZgC2qo02XxwffJ+bJbyyS+yIooG2ZpnW+/A
5R0IP4tbAmoPMuc9TnbiJxhpgwFXC9xPNRhTUYUs/GX7zV+fIPSsqpjB3SlsR/nndvaWOmpiz0De
sjihTAQbAZ2HXDtfyp8EqXtL0hr2Er3G4Wahyrw0kngHasYkE2tyu1yT9kl7HrstJQ71Y4tn5wE6
tAZzvB8vGO6ZOcXLHX+fbJZ7WS6NKpgjf33JC9QyXJ0UMRovp9c/hyaQnodQ0T6Ccw7gzpavC+R8
Z9+hh+f8bPpnsizSduMXHKpK340f/FVyuXEav9cIrI/7CKNikSSeofKXaTKa6hnzVrBtdoWzXtGN
CsRWaWsNtRHGEcg4ZiL3QMqshs8ZSmlvR99Y9x2mg7hkduDPaWIwbPcJorDIlBjaaamHDPkKXyko
oY+EbdStQLL8N8yyn0MJUb3xm2QoGRDb/l8tAiRTY5Uu79PuIUf9Ek3pDG7pgvegFJtjv9UWQwK/
GpPjxtZ1BGsT6D//wU1illfU8NaQa/2vHBs9WdB1G1bNOYHD8PzwBGRy1lV1s2JioqE2RrQMlMg7
USxeBX+5h3Ij9YDhQDJusodtG5Zr34Echb7sveTD9S8jx23w7RAhekRXYEF1zk0f+/vkNtw0qQG3
yI+klGxOcyxw4c6ayRvqIJmdVj8XulZ8WjVAhV5oczXzQuU09uQDL6bJncmONjIGzAB59mLz4Xbj
MsN/cJ/qoYatVkWSaCJLXT/8wwYrJ1i65il3nyBhj6VNrD4h/MRbgQG3t3BtRwRq7dC3ROFkvA8Y
r2YX7VS67bwx/sPnm2BMf0F0sQc/OVbwpeQwuleR7G3XuTFhrW+JeyWNiPX0jtUXbanyh+HEMtkq
aAnkwBX0+65oeBHLzZQyyXoDwYyXkwsw9sdYSQGjMChl/Kej+RyQWEEHFTtbeuc6vOCc1hzYzwAO
F9m2W8cNLk5bVgGbs8jiHcFKc7PJZxg5FZHfk0vY6YR3PiZC5+gqtT3dUwwGY1Vk8WTLMm8nJ35n
Hhbpx2NiYKo1IxzM59NRRv0yx0yRL0mwIgYTfPULGabRPgqi8tmDVSEaoxq4oO/wGTUmb+cMRBTW
ke6cJlr4O4QkQl/KpVHnxa5C7qRmZnA4cQCZIC0t4ZdcixiiCrN8jV0Uf2oga92VIXVLgN/78+6G
5XmNC7DEMVer7avJPzmIH96YFNnhZYyhq74EPcMSRG6148PwVkYzEG5nGNWHja44fc5uSD7S3A9/
5dzt/Dc6dva7lCzRvzigSBauVcjqBF3+NrWP6waOlUlLziu7Cn7oPZBwuYfSRoYhsOKBv51WQVaf
+Sg5+cOfEQwTbFRNUzm1sx1xKorfltZrxyxPHVwL8NmT18ccnRzrq96dnNlexcuaS3rkCuQ8AcWa
GFKU2UL3WQ+pBxUVB8md7eqqfkZWwEtQe7EkZcGEvPuFG5YeDMyH6CAi9s2QoFAXXbSC0bJ1qCyc
TRwdzkXxTBInqWVt/ZbKozJOq2llSzBwbB5exAVlaYIjOk9WlaOhV2yY/JFxexhupXlCG+p8FsjQ
2vP2SHAlD5M7gXT0Q+mUU2M0JSdmQ97EZYLoEGXbLZm+9WHU8r1gQU5sW3ntiWwNuxRDJgL7x6jc
aAJz59OQAOuaNxV/4+c6ocN0YWPlfsUHebkbX6aen202Q6EIn2U/6J3JicvC1IDP8AffhpvWsfCh
6DHDiNsLQXVSoNY3jsWqMMgkbNuz4QNbU5Csr1hH7GvYgYgttqU2UE+eqbW/J0UnQgVF3PVboF3D
n1BqSCDdnh3/vg2LbF8HLkubkzdm7E1JCLGDYYRM2ydcImR6kllVI7Pq0P4aYxKlvkPAtjnRiEqv
Y/3NF5Gv5adUQ4DVbSycC3VF+VMAwVbMR+fpbyj3TH10ie3wheAQ7quJ+vkbi9/oVNlIlcQZemB/
DdndfTKV82tDB2d5M3sQEWc1+rRwV92t1PRLaZi1iMQM1mIuPqMVG1orXHcXzY2yeS32UiUAG60U
OQT7snjxN9yxxnT03ZO80d4+nZoIwZbXU85VEkDfm6URkCDY8kqgXVdbVcM2S3FAkpIAMGp4tC0X
xVhTqY33pkJJXu7l8cWpwnYJMEVT1XujlKUa1iuc+3z78H0jeypMp8SynH1TMrLpoiVemiaWGKEd
YB3HICUJIKqVqqlc26rYgHWJ7mo+Zz3ou6ruUyaU4Ikp9OWOiXnjwK8SFt+zisrPW/dvEYd7RK50
jlo3qZoaUHlGxFPl9LuI24ZwpkSdjv5uoW4vq2Xtk60wZDMUBGskzTunPDZVdvkO1nPXptiTSDef
NTZW/nHHWVaqxT6gkEZvnU5m3wL1biSgQY7J8d0uOle1RIVD7XrX09rzTw1xI9tRgAKPyNARtP4V
Dqz6Uj4Q7cmKh7sTHJy9l4HY8Z0179Cl2+5hTyG1Rds2tnPhst7yLJm+XKZvAdksrOn0E5hEw3hr
wm/d7TCM7vND+3dn/85I89cnw551XT0XWguGM+0/uakgMz8GgLSmJFUTuRDVlmFs3oZGgQIaiW60
EiW6nbIs8oLZmUTOLzF2kKrPS47WVfORqv/ECmxfVKPq7anMl1GXH88MIruRYotnDTU3QMqclEO+
KLica35rhceOsAopw9Xes08C0lxONn5PcXG0vS2U2zbHK1RnTIaQ3Wa6HwDCQc3Py1YoagZHMepC
SoEXwtzQK6NMo2bTzpRKHXuLGvIFUAO6YcC8/LnsUnsbh+V7f+7LWgFiLGNIZs1oVX4Bt0g7RdQV
dJFvxTzklViO8KhojPws2eSqS29Y6q6EDamSzl2mfcdF2/LjUD6oXUABIwHHyR2Mb10s+jtUXMlM
Jabb0GR+I5q8yJmxuS4z4IenXtnRlBm1H3HFdvlidNjwuvWMYUsY4iw3tzavaG8Wjrntd8+d0/T0
hjHptt4eAOCrHMBrqJt17cMSGs8moxxk0SGRHtmO24xGWB6sP8irqgGT27SbNyz6H8iC+ZX1VLnB
benX6Gmbz/EOCQGty/oeYa6O4MHtJ5vv0xyG9wj4PT2s9Nved0/rG7QAzhUzr39RUFI5Tdzh5/Qa
SwMeg4+wcvHQaprKhsGaj9bz5WBIRdc6WY98RuXcyUNng/VNHL/ICrKlZywgpQsSCZzB5NAaQ5Bk
i/1m/nkIRpmd/BeHs6PK4kQH9vgZA0KzC0OiJAXCvbnqnf7VGtdOlvdDeaUIp9zooqzQGTMPXiLQ
uN5bjHJZp2VwrK7t4D791y+lDu7OSnW2xRuvpMUoE9nqN0xoidsCpUrqhMfP3qKBMLDLQzUZx9hj
HV54MrM++sEfTkVCyrs3A7cd04kL0S+1FDp5VED5wuaFgtKvJoOIpuQs2w+yC2s7t42qEC+Bczv2
9h5AgZn6f74YtKsKpzdwG2A+PbCAryQXlqCYRP/naH0gRzjUDqFePkUfHZLW8FnZwAjEiAkaKOr/
VVMb0EnI1+RdAacMJBVlu0ggNh59RviV+ieG/4fw9gmwBLn+na6iwlDeK5UDuIrhY8UBgb8iCaRy
GpeFxUMjm4BDS5l+WX0cRKLR7LTOdy9LqAA7UQzVml2sUtZssPk7wrUMWTIbQZIFGzNIBv2HjHnT
fRCkSmx/AsS/+dsexpZlZrcVBhuhyl/3SoKD7nQk/LKeH7LkMNmVVyWVnAOwRA/TnCvG8QtMYzK/
xYFE7tQnGB9rW6LFSJey8qmY+2EFu4PwNnBMSt3T1nxnOwTutAdh1NKRRZ9vsltBnG61++7m95gg
J2ROh/CnWkADCTbwCZK6P8iUobbpF2Omd7WL+FIesj+MKQU3tKpubUvQKcsAnd/zrRxDUNA8NmZB
Y3pyxUgnyjHdDMHAkjhJlAb2+FcLrXyLC0w4t6qlQRoYkAzo+PWhKNbhgA8/MNstdTSzlnBxPX88
Qq40jH6NT/7x727Hx2VKHVRYdEMEqMJZqp/hbcnh9kER4yHphn/d8YQ4a2cr3D6K8cEvbJHe1XvU
C35wQk54ITkJthRfL86OtG6KhtFj5F0ov9v04OILyebwaYeW7D9JjpMw5gcIfkRI5OcQgnqdn+7T
0cntdt08bWZqTSRUyrSYf3I3pNauMOuz1rjEYENNKOBXcgeW+z9J+apOK882lOjEFYfc6Gm4VhoW
uSp9rv8LnTUXq0UwQGoXo/GtrZV3fNORrL21yfhAN6RL3QXHfUAxcCYOiiWRmeUHXrEtdId591Yc
FGZyifIyP3XCH+FZ1WTBfqM0LNIM5ov0dwcz7ey31q40UoIQ0iCBhUwVdEN53WdGegXBwvVaoBaG
VvcX1CUM3ntiNbGmaAwAp35nxCKTZjGpwEWzwvIpkEvmB7Ra/krc2fe5RPgHC2cEp+umHbOlOtdX
igpjnt2Aj1e7vZVFYzYSDmKJyi/7Qu7Ltetiwe2P0IBlWK9/YKS/Nw1b/rIye7zh110wOXI0UK7i
wH4mEWsmEj0A13f2OeDE9kOZxU7mI23BUTmt4Cvfu9gABW3pzuUKVKiJCw0s+4Bj5bHmXm43VwY5
2KK+QVr+hRUYAZol6FNK3fThclKsFH48gcMacPoZjlhMpCTAKo5KId2bIZPAmGKr2qrwShJuzD95
aBh1DxGfI2JPurQL3dRHQt3nQnB/E539Rap7TC02xrMgLq3yiPJowtWLnAfjF0EppPhuCAreUv6z
RgsCYWzUnTdOX49QInYOeBwZo3cGEfzcNnS3zTC2EVj9bkJ7NDJzlUuH8mPZwOETfnhmEK1tGDwE
OVqaZLwHZpRji8fMj6PzoILPnwLthctu11kKZdwUZu+QV8QorLZuAdYTadaer7rDyqwMforU2+HC
QRn0I2HcRRuRdYqE7jl05IkTYAO9jhTIT2OQsEkUojy/JDPcJPX3+fNe4fRjkIy7Cx/HzKy+VbjB
La9yzNdK4eh9Na9kdvnxjhUf42oOXMty7dYZe9vuNHNAVQmBHlTo4xCQh7O1BZuX2zJJGd+laTPT
L4yoxsoqT+cSfqGVcnDHEy6CpXLLghEGDmyh3YXAydMAOJ5KDGwc5lzFRS5L2U3vtZtPQ3x5hpwb
lr/wonBif2pgDDEc5QdDilNCssAGf06ZKDd1UCSoZ7Sc0aJOYn+/WHr0URsE5iODoF/qhG0YF6hH
cxACNF1z/5Ff/m2AZWwnk134zTZ44tFQzyHYBpX6qJ1/rtubW/HqJrzHPb9iubZJmf0vDLAiu6G4
B80MRBTZ7cn1efGnevoJ8zOBaYFYhthVJ4Z0ylvv1A9vDe7xFyEsMaBDuDG/LJxJ2z3SsDQt1CAB
qpJbGeFiQg9I6IGXwRD3Fc+H8IZ0HYSEP/+nfSUDb1mzERmZpJ8AOTMziPFBQh85+p4HWG6qIjPG
WTiRdQYA0t5ZcB4rkgk0xCtGu0Fl0to4OXJjBmEVdSzDkuLwloadqroMjX+Qvz6TkV7DMu9xFrwm
3nYtnoOFIzoVsNJxlGjehByZv3H0EVgLmyjTC1dI7M2s8XPRcT+dlYP004TxYK9AgABse4wY9Rei
pzv3tnxi2w76GSbsc+EPR8nDlO+RbD9dZ3WU250woKTmUfTF/XQpy+/rnjowV2Jt/45GGmQtAI81
O5hDTBaGnA3eq6DiEbDh/Myphmoduu4aqVMLqh7/iE9a7c5qhbRv9aopBtPQdK1CbGlkDWzwurnp
ES8arDt/oKF67pSB025gtsY/oN0S1aw1Q3We+9+cOsotaE6/pZLjJcO5vb1Q+mlvOltkKTcpCgRd
VnTvNOXdgj6DJq+/evFFpK2o1UxJYhkc3pu/FHhP0OeGqbR7zSWKsQPOyz1hjeJolcXXQD//L4Ld
UfosdqO06aLZDlKREdARU1vEQZ2tfmG1VzfBhDzNXNxWNB3XKqKUTMSFfcm+WKzmS9iNRWBpWpyv
e7HkCrYmOOo5xV39leln889fXTGJ0wIPlqcVGuILGseedbnBC8Ff2yjTHOkR1EOT/z89kgGuYVXM
hyRK60ml8+HlB6r+OJVT6nwAKSkvavJvz5f+nrql1VB40SoXZfqnvyTe4sysdFiVas3YqmGbJMwV
e6QcvwL5GQQZGjwZDgHKPE0/wqyO2Z3eO86svyAKBz4ZNTjbppAzpN5lioMv25WCgy+WpLgghvM1
8bSeThwJ7GL1vPbtTbu5lWNIaPNRRDlonY49wGy2goqR4ibeLbkUqALoUokRly81mEQVcZLqM2Q4
NmbBF7h7Kaj8uLGGZeUwEp4eR+cIvNSvsEnqGQ/e6HpbAs8uhRzGzHaOei0aA8UL+kR4n32rn/NQ
1R3Sqot+yf8sUrlyLjr7OP/HU5qO3kVzPYGKNMjYbOKg5oDkDZ6aJb534SFXA0tUYfMfrT+8nKmt
XhmOiDxIl2RNdOGUGgRD/37ueXO1hS+hKvn4V9Qp+HS9RpkDtuyI5dXGY88QJz8/56yUJd4QtdIx
RJfLjjzq4ymlKEhoj+rkG+N4xqMlAv9wzHlrF19uPkcxalFENDLHO0EeY7bz7hYzhkn4MztYYpwU
N+pX+4novW9qhef16JoFKWBoqaLV3oFf1wT5pOzNm7OJONfu+heH/0FemhN9vqss3Y65Hk0R5gww
2vxnlLxYV6uGn/uApY7nHLk/tVhhDAREwa/1jdT66TJ1chz4hXUJX6hCv5NzT9Hxgigc8HwcYzUb
dsrAqhx0voXtn38SxkTNXbxV452BOV9XQyZsnKsXfSyQJ5zzFSlk4vkGS+FeqNZDOpEImLLJKgox
FVpoG2GhBF+PM5PprJ6uqOWNilbNGqNBfnEB4P13c9OHwag6Y2mfExBFFYrNWIaWxb3DiYmDq+SI
wfxthw0nndEGBb7w2FTIpKhoY7NjxnvsjuVl8mwVz683RFW/swaoNDmWbzDRfS+D85JBYkXLRgyd
7hoaVjV/yktAm97JrcFU7PYa6eS8s4H0MXIk372yeQ92u8lyHE+m1Qts4QY0NG/v65l+7k73CqmN
6dOG5ElFCPTN0xJfzqwN9o60waa+Vkpt5d+RwcgF6VFVRpbNutGKdYev4RrAXTFmKPyycqBCSo+u
DH5iT8gZeaDIiLd//aXHxdsAss2dqBRD6mke6zjJAyiPJam+XF/KcCu9c5VSVzkIJTPb+EHnaSAu
t7Stdw94oeSM30A1mHzN48iZf/WZtv9JpdzY8nlf8fqBbNgvZfM2r02GG07aZC4VgMRfRaujtttz
czuv6dSFDrmSMOHB7plZsjL7ruE7paQrCbmZMLWScHxYwhbYg0hbjtfS49fuYs+M5lYx68Imw5W6
6rfGEM1iCEEna1P43puNQoCGMyHyhnkq5O9+39p26cNLklownSG5crbn6LlQLCn7ev97sMtD7nex
TYWVPGiuPdeVGTWb+MtDnKkIiMnYiFEIgkCSCkpASJGEe1XcsASUBK1SQEnkz3HI+mAvAE1qiP1d
an3OJehJph4r/idiGP5z3dDpzENfVkBb5ZufU4fiyPXDJZqXS3dUy179jHix5f8QTA9OwD8NkjU6
HAiACCVHTMtx7ccvLVSIk0zoBwyPqxMsqDllZJuxhvgB4cStj3ZhKk8tFhXMC1Qv9PdluowcLmfG
LH+94JdEwDUpItdtluW9TvDJIc5YsH2WMQsjI/gMjKHSvPtME8LPIJ36C0hplrO4HV7nHDqFPLKO
c2TInC0XFRPmZ0mtd+gEID99Hd3XOgnIRtNkGQGSqHqSi3JlNZddwDZZaxhaSe+cwea+2Pvh0CDq
reQr9QzuH1Ji2BpTinakBV4hIXH90DYgtm1dqM5cvut+vYgYASPxykpTDvHsBXBQ+A6Dvp2WtmvC
Nn5ZPc9EGdqtfNvaPAKPqLyJqYDtF1xwuX1Ur9z6Tc2P7EgdJ4Ifmy5Lb+qdZnlPpI8CCLkHMqh0
L0TFbkn1sRZ6OV1ZGqZUwS759IMgiLwwEbIV6ic57gml4RgBDGXdgZKwlkb9zJeDVYjjFTs1Imqn
2+lZ+JrFupqXQ1oPxhf8ncogm3RtVNushnz72tb+cE5R6pdQb6rw8EGo7SkBfrNV1o2K0SLfqcny
zsaVg5MRbtGR2anmvBhYffAKHzGm7m+2GqT65O15MEBFrJSwNNHHDk7mV8aHplxD0vejvDwvSRkL
j2FLwU/CKTNsTeE4qMEQYL6HhPAfv2C0PKKDnmNTJmfjPCCkirut0E/QwvVavMgrOXS58ljJ3fDs
dSy5/A22l13yM6HPCGGIsn3Qs61pzM117xV/nF10aZfx93Xb1jIzNrDUMCf87dcDFnkkbIvZwqy4
HajZAQR2JWfESmKhLb6uagGP03sdd9bS340NYzImqI9thLeSPxGOrvhHX5xy9B+7nlD1WuKYx+AH
Brv608CkD4FR72JoUQWGScVFFfnWZiYliaXtePxZ2Pbm+psKvFw9HIRpo/E+cSGu64ZnbnxSeu1z
7+OIi8CxQLhSRM5oTf7eADSnOQqz6sDwgTMWYJLc6eYibSMjF9hU7W51BrvABk7GR20zem4DoOkY
/51hOcESR2W4JinD2mq3TKXed9/ug1Ouiy7kIpmb9B4E01aV/sWizXiu2AEMsS7jpfIM/QNqvJCW
TBT2uaGS91bohnqXvbkCbLoHGi73B9cqE/FAUcNWJ68CrCizztYrJYFEcoYbZxpvEVLEaisMlwsE
jv89AOrdIXI5W5ozek9pV+ZX1pdX8Y8Uv2T1Q8GRxrthx/muSoIDnsGwcyrhjV4Jyw9cHA6xly9C
AYy51BvNxBPE1Fr+lNv0REJc55Fe9f/mDBT1IA6ny+Jd+hpEPfOmfMiMp1NjRWk1Yh9a+ATtFiC7
sy13hZeqsVUZ/cDdoYUthwi1KvwDTRTYVMNFJoYFSP+R3mV+L+WVqQ3SppIJE8a7VNgmum96RqSw
a8VdcwrhV13mQ6ZLPs2WAYCVokhDiwX9KZ6iBduhoHvSrO0K0RFErLEaYgGYYjzmO40Wp1ZS2DbL
9/IxlW4/CTIkGyyQAhdPc1h4bpeuTMPB3uDfJUJhR79abSQZl6AnZ9yfSte36Zz9S8oGk54PcFyW
ctKhFhLUhqG0x/O2ZzO7w5wxzE/9FZEA9HJtwUvBd9OwXpMk2GuT97KBchYjk48T0Ep+FXJCB75q
bm33c0vwuL5hoooMS/vlSLa97voR2baebj/ikFbrnOBgFrCH+UGs2j2dVQ8ODvZTrUhztdViydy/
jNLt4f09ooYdixhR3APhfSXJrxRejw4ZAQtl+vyVBDrULTPcZgCgArJB0aKu0LsqqyYmQzj5zQBa
E3pTzzf6NGvj92fFnAMbFpgwW2ijaQgXlrJiPLUemUPBcYJY6BsTtTrgtXpFfi9hwZm1bu9uzlTp
oFqAx63i5HrKA6g2I77Jpr2LnV+jVHGYy4IS2Ak1BDybYe3ewz3j4RcvcYoYe4B3LPOvNWeB2dCL
hwham1tI4mUXAbqKjYrtRVqpncA0HuXT3Kq5MQS11seKhP1xIeoAAAZb8Fb+s0eykO7GkOVAcf3g
KbBXtZPnfeBUoiCYdJ+zz4U9arnI0nqQ1yjSDNr68pManqo1vg3s4MLZFaAkqa0eeAtFNf8sFUAm
BHGEYksdwL6koOWZHsCcpJ05vaEmHq+KJp56qHJAxqL4gb+dAU7ehKxwQ47AnNkGhQHG9/8i0Bfu
HtEP6+dbSUSwQ/CaQGW0JTB+0TAlolsXooMqexTvZtv5fEiu0JUoH0bzSlDXyD7dspadunHQIVlL
FK47eLegNiG9m/g5/7jYQDPkS4DFq9m8L5Ir7dqMaKkAh+xb1m4R4EbnRfaKxr9Kwr9srDtfbQ0y
rHmbCtzx5QqC1ntdP1NKimE3WIiE258jNqfnglo2wi5IFUalMV85Fx1CQax+nn/aw9qLpKoEnxS9
Hx7C/VyZqBtPHm0yCbUoAyBLPg0XQm+09E/XxT0G7+HsKfK9vaTBxnc0B3QoMfZ0Ulo8ShR0ycj0
O3oafPAlPs7AR2BIpItx09clua2MngfKak2vmVMN0isCLMpNUQFXY425guaQop+dOxzWlx/iXMSX
mZcSk1mN46MTeYkc8detU3tyDWioM6E373y1VPyzFHu91n9luerdh1HbgyczLbeMshkLGpebW3vw
7cmojZTb8cKOHfLG2GZSdAbnYFC6YyKPafDuHgi+mHWcFWlCU9NVTT+0GWHFNyLUnoyTS9P5vHIt
m9rCwmEF2t4LOIzcZKMccyIKJ++p/FrkNekVZ7jejrNZnq/K/C22uW51xnzC7o193DcWfR1oVQeZ
KQjIkeUofClG1n5msoYwQttYd/T7P9ErgKUbA6BPLnANZgAftEfjVM6xt1Au+Q2XxThFlV62zCOJ
twCe18yLgXSDgpm+nEGVHn01W5bq44onSPBLXkS3p8uAHOFytQjCclViLoY88Fzofx/SKPmsy0S6
nINM9X+oyrvSKZlim0jr+yaqEvWSQbCrJHKfQl5BJUrORiDUS+IEuf7fgPubdIRX4TG5JOdPnkK1
Jm29bcVtYW+e1RG0hgXDgBudfzhFN4lZmAeIhAg5wYD66Yk7q5ZzH67to7mlkMu7NL45MRdCO7Ii
xhl19vhsvqtU6q2NtRYc/wHrXk1P+i/bru5zTaYhZw0rwvcbvopdFhz1EesOu3x7ZgZKEp4pPG56
AnX7zA1TSuaURXEEQgyA2TUo5vdvIwwkYaHCKFwHJrEy9Qwz+4B17sHHFbMrzWnAUbd7V5hyxqpX
s25kr2MLH5MwEXdh/2Qogs8VyEsFKDwRRiwc2v31fnMUxlBIw+hMZ1EoTvcutc3mop4XjINs5TvL
z4z2QxPQWnI2dohtoLu6sejGglb8EnydMyfrZekCcuRcbQ2yImLLuKdsaGNMyYAuIkhuY4xYKQWf
KiVlxvGHSsuTrOGzAASpQrrK6Y2B/UDHPmKLS0nvCFLKz2K6oj1JPB0F8c2KQQwFRyyNpeajFj/O
yfd7GPNrUurj1Kl30MuFVz9j1QGL606ua6V6yFcrv+rpdC1/x00gacOoir+CBog8RHoxKGQE/vDo
LfMysbbV6suOt4sBEEsK45Hd/KVzBr10udSFsct0ScWjTn+1fcvX/fwClNkYFMIfXOYGELhPZOGS
N11Fo1FiJmWZgZzpUmECEApC0NMwqN7FJPE6ve0bOOYT5bjsT2o+fgeitofb/LM8WWIs7vmDPxKH
/0lo6yZ8L5gLGm4EHSSqdBRa2Plqc/oELADDDfsJQFVgfF4lFWk6JlrDtdirfOioI5cx0VehRN0+
YymVWy2IdXn73+L5DdEpppTPrK4ySNk8l5JnF6gscXwaA7try8/c2MwjRk1ztz1QiarGaqxCMnM/
J33bLrnoMAdT6PcnhTRsR0N3usA0ST28OEupLxZPkW3tg4I74wluzKOoKC7rACOO02vYPsA42UvS
ClkfjXRoGTvse2pxGVSUbDZt571Ez8oXs6HqxJ36rCh5x3v3LuDAtcmzVEf9fssIB23ViD1A2cbB
3PWR5Vpr1EmePB4uSTT4lFHnMy7In3fKkIOWeJl02mL5nNt9F7aMmkF/FVQDbKvbfZcepiHvZ6Ja
s9nB/xxbEuf6U77siOyivLVvNPuRVyAjzjOE+7wHoDMozlTLsYFvcwRc5KkfvOzipW/3HGC6nDpJ
pr018ejrSNL1kkFvZN5zMe9y+JaekkePggKXEGa6c41wFDk5eNE1zs6YWk2RcKO7r+R6FcR051ku
PHXxg5l1oRUH++7txbd3XfVjehG4jjFGUp9fD2BDYAv29W+j6Eaji4TKwGqHhMy6DnUWGjp0xPv6
f1XIs/CHG54S6P50GXq+Vjv9ii9KooyOPDIhr0mJVYWNwAMeDw76U+6mcuQvIBDrN+GDsGFE4kNm
OfUEE/65mMuQDKLZgxVzsxk5HfTE7hGEqCbn7oN5l9pd14DvT3NgLS5CvH7Ni4N3scxTBIS0J+v2
AbQXmTY9sou9nPDf2pIcReTMpghfPCfLzeMWLnUw35scm3yfRFJpcK8rgBqPvjjKvEd9F3WrVeBg
DD0WEHd4blsJYvMfV3nLV4curPWbrtBjsP3ODXYJm20/rmwWUX+oTOWh3KU1cL0Zto9YVsMJNRBP
RrunhEo8hN0VeDk8btBbXHZOlWFDP73xVpMtXMpyImy3Qj32bkqlGP1aMxNN9ELjfqQ2Bslx7o4A
FT+3pA8l0LdHWxZ2UC8RCt1wzZU4blrB8imVRRJdJWA+Y+gbToBfLwF9rSfPo9hS/qfUub0U0GWW
j8sEh2JX9lJtKUpKiBEsoeDlXYhqcmzrKsmsSv3DSG1qjLNK12sVJ0ObTENPB89OLlbGPn0SfmwF
sEx+9J9iFR9oAGjykLKYCry+M+KfhveI32y+7RSX8AFfl2PJUMM2Dn0+zByNz09rgknC/muBSLyf
YKXodfrdWYAVyFfQEFTqbQuVNSy9jbOolpRijCgablVWxA89vsYikaZFnHf7swYIQ7qriyt7qOIZ
YgM01YraAYyjo5SUhoEEFat0zFLYVgFqXb5mY9+RFLfexW9rVzTPrcq6DfdnXi1y0ASsIYznJj9U
ngf5UjR2kNp3rZYTmwNeIlovxq4g97BrdJ4lEhnaoxAmxzAGISYKHaZNor9gQymlNjqOLTyV34UB
nLhr9EPm+N+hyPoVxq7t3FGakWXwTPizKY+T6XtKZjjyGYpVuPJNQRNKUzBnXO9ALnopFlAMzotG
cRuVKbg6s+yRPOOEauhQrQtdAGGU9VKhiunfZ8ibLkuHvDANCXXyNW+lFJoSRCAWJdTM7d/VeC2p
jixv4XhI9pphWZj8KdaV+Ws3yjDfRuJE2Z6uqIEZQscaPaqLnmV0DYsbps4+Te52SW7GYCaNpeV9
6wn4UMsAKfZ00Bcfntvr16AiPK/Czouc9T2djPqwCE6qMpstQKaYzk9ninqkkq7FHy6xqhe4pDPY
ZXil7L9m1blAVm52sz08jo/cn1MTvgKxTCkG2KhNkGczRJu7/3pZ1gL4QfvnC7JPYi4jvVN0zIbx
fd0XzK5LU/0yI1Z3nkmuHtjh/LvkMO9WDxC8F2riQRKueFg4RbCWXzT9nGBkueLYHHjM4mp+7aBd
LRf+LhoejDaT3lEfyVTOOlPfrpXizvO1hTEINFAYjTlrImAtjERqFjSgESXkZ1j9dY/UVyenxwEP
YiThwcU0+WvdEwGpCCdWOqlKPRIWi6GceZef3C5TxtnZb6AMhQF83bymywfI+R0D3ZOpA01radd6
WooVNFs4lV85G6nXX3Syl07DRl3l2/Uw05Uf8kQvYr8CPpRxCzbnsmww+rUfRFy9g3xkbJ69R4Nu
ICFXm+pvLh9gz3tIZusFKnoU8aiFyKVNG7c+uPvP56avZrRjDvwWLdOCcqnIW7+pVDpuTbjwq81J
Il3CiTznQTvDCNhiP1ShEs7wWf2APqCUgJAOFLWkZ3QPmbkkyxwmgt5EqS4zE+jRWu3J1aE/AZs/
q2h93DSKQdI/T0D3Owe/8JAKBFKFWrK8zf9noP/N78trOsxipHLG3thzIlsmhmioOkFAVSKlxxAo
HJvaKe4FuLMB6ujShzJPYvikEf/nUEwg9xs88q11cxXWTZB6WLtIWIKGydRvHuLCm3u7h3sfWIvr
f+4DZBzdYcU3Hk6uDYunGGANC44UKOLTjo/SwpWP/DqsePuU/Rh6fV7UhTvix35Jvo4M/NnoTGgD
W8D8EoEyg+rbhz9Lir9PG1+T2HwXzgtPm2nAFC4QW+aJSgE6iiFthBl/t9/kgprnm0a27SnMr3M5
/axEgFbnYg8TMR+CleQRvhYxOekU7tFj5+dbxbCi6J/TD5BA0AQ1xQ1EvQuQARw0FlpMRnKOgRl+
Jtl9W0cC42ZdNB/qLFwtwCSc3eFX0uYDKA4Fq884YcpsD5h5R7i8CSZLb5bcWknUvZfmiv6ZZYPS
rPWuUaTSiRSMWZ5DH+c9Kiy78WIPGiKzOxxq+rqNqXP99+juZHMzf0n/96vWUTDKf4EJHKZi1r4w
BMtjlG4SLVaDSO5jdfRJq17BU3bN27KfSIh7o/E+CpGitjGAQ3acGpZDXgsFG8KtWN1m1yecLrW6
ddmceCHG0qROiG72fU9LqxZq48VE6SKiVWpAfMSa/AZDuIT0DMUI7WjX6q6kY1Q2GOn45foBNCnc
9Vkd8EzgMA5/NHzfXQr8YBqxx8fI+5LMlWLhllKVKD2Uj/0TErXXFBlJurBJr8nIEBRetgeS9had
/ttDPd66U4bQpLsiyPNSHcaANuspUwRbDiq6dxBgeqpc+oRIthXZv8RO9QiV8YiMgiVn0BFyi5E6
aMc4QCf4TCVAMcnNougNiSQm1QnKRfeJBJdJxUcME65WJEbwExeUlPG0QH10SoOq/sdXfu8LccUB
k0lQsNvSE5ZUBE0v2w7jAlqLg9Lcd6bq6PXS++W0IVwHHUFBpQOXNd1hGD+R1gyT+nutr0M+MctM
lIBe5jdvhsvzbVSoNuIt03CIhqg5JeIX6YrjGANPZm34X5Nzs+qvxGEkZEOJ9l0aYYzNgSOHzAMS
ielMfHNVxRxkIBvZ8yQeigQsMc6/dMicrdwnpH9SFK/pRf+X1gkcuPtemXmMI1LOkcBvvE5nI+RL
HhuXLAbbRU4NXYiIociynDh82derOJJ+F4yQmQYGyOgsSYXeIFPKVvHeEqQ9igKZyq0Mlgnw5WW+
RlA91g4E7OzGzmVJTLWICUQ6vMhvLOs35C7HMSr1fi8y1fm6n/ZwYZrjPdRG0NFtzNIxiWOYGaA/
Zozc4lij8XgkaDxsrAXFk9qUwUrjCvYX6qkhAO9WhaTWX/fh/XKjbz5zjlKSoSis4YvEUACr6Sgj
TUveCwoeGXUDyEBYpGaJ2wkwnJXapdj3qmZHLmAS0XuvcR1vooiITx083clOiOyNZwzhSP+TZ60C
Qix5+zg54WgJW/DEiQrjSn71s1IqjsV+3AGWcDKppgHDw3AMlK837TfxHR/oLR/iQWXR5j9L7lLj
UjhGgPj/YrXTeOc+/NUxgjx9K7yKECJkFglOoedsD+ogqHwWQCeS+02V/Y+dbbNhzP6Lkbcq4fSG
K9+TZPGnHc80FFE5C3a29wFLEJllnhlB6LKRzUreABIaXDV5sLwQbRBJlN3+FPt0bUbuTjM484sO
p2EzjlXkSTNN6UX4AB9Q9v9x6kbCWKKxLLzax6m+uFEmI4ocPBZoAipNUOhFgGh57j/qPUQ5C7a0
f/Y+VIOfmaQmBi3M1glg8id52CDdIDPiy47+JN6XfzeLalSLIYqS/lQah7YajI6vnKa39a0Jry7J
Bp5yaCyKD2j0lvNuxVxmdaVUCEUuJv2EnH5VeSi6kanp7d66mF203/LlHv7rV2hxIOoGvXByTYf7
9Y6mX/e1gz0Ciy36FJTO5o1Uk+Ds0BQJ0q3Zq4TpSXMvr0my4NQRA5W9FYYV0G6nu0o3f15zEmQY
VF4z3tBj03LT297vqyOSYNVEv3+KcbJrJBqEVmtGsor6T3aPE2M+Kb6/cxlIyYfUh/BXnWuBiEhf
IJBngicPbZQuR+qB3DaawNh19RUMveVNr5dZ0f2eeSk6krtE077kFMp3ZoFTmv25qeYZ55cDLG8R
cf8H+0sWPmWdWNkoVbgC4EcPXfdLHVKNx4WoEZZFCHQk6h+J2al4VVbMlZWyUC63o7F8l0SCEaJF
Kj3LRvpGM/nmiC9uKX8JXVyaJmWlmuT6nHdkzLLgg0dGuKqz86WFUvMoiFby+qJI8J4s9bsKyTCu
015pcZxXOFsJnlrYTPEPrVKREPYXiRcp3r8e2Gn1jULXx5wj8wZ3Pf+NixiI+vzLRaKazGIWXA4v
+sVJZi/O9hVnCSklREt/6IA/IFL9j65O/1epzFzUXO9UNBM5QItyUJZ9Cb0CmX3lHhWr7QXQeWyY
SoCIIKq3L1SvMIyNjyQjus2yoD7Lq5y43E9pEpnZ9bcA/4iSec5J89uZPg0fzxnCYNuJbqsk9HQI
3/AoHi0PK83aY019UlAOxwYr8er4iE7dKuWQG8thzc4TgPU6DSk6LymkWaER9lHLvMs0Y4Rt69Lj
3AZzDJ+nrUnciXMNCSB9AD+DvAn4tcXRxaUI3h2PyEFd8sHnv4AP4NAXQmPn9f4JwtKNk2z210R7
uXB8DxVfD1lRMeIEGEwx/WTD4rjF4a2BbyR07B4uDsjjT9Y38FvfXZ4xehH/+rj8ULUsP42zIBiM
uyzNuHwR+fYq1veS8rrOGRQln9Z0d+WQexWmGOtqYQZku9xwmdPx3TqYdBoHZJnaZkDR62E8d8D8
dAoEE5BnoAnPTx7U/17YMfRXeElRbsknKSZfCpOfJjFbaIi06JDUhU2J3RyKjfItgSNSkQYJqGiG
ZP4WkUETGrqJ5cZq2xWju6UzWY9UX649pjpCaSA45dIUcVpPUUnbuQGzgJ3QVnS6yuoOv/kaJYKS
oaIIdJ7NoxdJ1NgFc4k6VV+4A/S+3SwFwHTcQuGnGjFqoSZ6+zEWzNDvCqCnhd9bnDp0AEg8CwIn
EzwDmUFXaNeEBq4wMOJni2zVZhjrSUto+aQCIpBh1ddvcNLZtgcl+ndhvIkxl7PkHWmXeH/mIAsd
indk7Tz8HnOrqUPDSxxliXCngq6wXC9THqbqnyc9VF6YUyiNVhB9eMc/tZaPvK2KsGDL2LKVeMuU
dlMhiXPWzCVGUGkiyF3mbKA3nGzYcVhr5BW1Lqo18KaBKWAdcfPBW6DaT8XPJOLYkUJeTvzOuXR6
3N1GKLY/4kOeN0ubDKsm3Xzu3+Ascj3lmySU3Z2fcsyxHCFazcpV2NcOQdwAbd9ljCNyCAYwQpM+
9nf8ASGZjUTTZtimo5TI0ggJTf/eoyA5SWvvhIqIHFuGuSRdNd/DRhLrEJukFjX0y9v5XiF0ePq8
gM6h3xjRcoLFlcR/jyQIlUo8UVqtDziQj7FkC3GbdX2iv9GiiUCZaAxFxSJlrxBMVdf7YDS1zbfX
EcBXwrHp9HusLb9gKVUJbIkxthY4t4D590tRz3h/uiYsWLNIL6HYN+Mo4brmnWT0xksdq1NTHhBf
yvuwj/Ep8QCZKKs8/p8NLdOekn2x6rbrMj0yHvY+MJOKUmaNq0R9VHMQaCBQWeSTNgZ8SXkez+WB
RMcB9AqJdqN4stxlv6MYdZGVT+d2IHcoAt1NYfa4INMO7tWYVt4ss34AV6V/kAhXBbV2KxNKIIVD
XKldbk/dKlf0qrH7D1KKMcBFi1l8z/BKecyjeJ//Ln39xLRBxM0bEZEsRSf0Wc8BLC703Pw7CIoW
mGmG4PZEL7Co345bR4SydSEzt8jx3OIcTLXBLGcTwjhTCLvXSF3dDp7dHef5ZX7BMonLBGghiinH
5uI1Ahd72BIHx4rPt/Ikf1YICrpBx4zJLtAud2IFvtiHma3waRezTpe5pjCUHQd7rifhKP94kwkN
KWR0cxBhSSeu/9dmFOQnCpI8naPB3cJ0nk4w0wDpXSiLDzKVwvH3EFOEYgKcLzaoQVzuGRvh8Ytq
i9pclrs1ilIuI2NO5XnoEo0SmXYnxykEDEXRwE5ja370eNIAtX3zjo6EqLhNnRibV2vI9BUnxmPO
SZynSA9qNImMQ4nPHjOczTselboQ5Ka/lq0bLtXexm1IMgZswSKvyysR/RLVyJs/LGHNHJ1axRWK
kULKQetPMeI//4FV3erhP2zKxwPlk4vGKpQjhbPUq07Ruu582MbRaUEfeVyfLFzZt+AS75EmG6uj
kDhkiA69GnwejGTwIVKIlgLh3NrUOAW2NhBjRHEGyuKiVHbBl+IXsm4yNh/yoa3al1F1kXl6Bn6a
gJV6CDUSBXzcWdXBSYvQEJUqBdDIPTZzJhOL6CSlulOkgGZ/ZkqywSFGg0MnpweNVKxhjDniORls
5N8BPs3e8okAphXK/9PMiPtBrEuzL5FCTqamAB1RbRKmUlYEYlH31v74abA0UJw9k6BgaTQtoBkp
4kiNhXIQBlfgreBHZyleOZXkNb67xs8rxXq81xoBQNm+VEUCNyvPxGgRmuEUEYdkjqNstyqzS5lk
lMLQzveN47VdRzbHkeRTwdSXNDPm+66rCtMqr6KGs9qnLG2RKKpQKfAvKNXAP5iC156yAlUG1qLc
HGFyPU8Ncb9vUqXf+44dUnH2CbchYeMtiVzwfaXyJQ/V7ck74ekX5HJfEBJbfnItu8TuesQdTOuA
JODgRJ2PJ9eNI6+I7XJDvORknZtTSbE4n6/JN8+OnPbtm9bO0SW2PNBD1hH79YezZSPGF211ytAK
8/Eln+3ZnYBPNVv7pNihirt7Tefxu3jS4G0G1tjy39Ke3qnUGtTIPdXOpAa3O2jyJ9+Y6rc1kpfK
ccdWwRmmKDHZytI1vLQ6ldTj6qTjizQvSwBgj5nxAmL/eJyuVrNOmoJP33yiPJ1uNtjVD6MMtJ0r
uFOCHpVumldLDj1Kdj1wOOA963O0vOuMYUDTpDPjyQJl+ZWuUUpXvq3BkU6u/pe4E/QJLHCUK4lq
CSilTlHYwefArrWh8vUOK26TPdJz/DJbZRojQKsITQtxOVT9DMP+0SkwYj51lkq8ghp8r8ZYv6yM
Q4bwEe+VB7K7oR6zvzZitLL+PH7CEz/c651CPho55FKHgAC/amn9GhjHnkB1VMnzSZwz/l0DttLa
vtl9uvfDk1sazvwRQeMvb2TsRGFt5NeHJUmoevtov5qnZqitnvC+VOdNEIdabDT4nizeLAr7AR7M
6Nmv2FFbxdXc6+QgVZp475aIL/lHfJ7XX7TZ/w2PjHVO0R4iRIJ0R+yx+w9wYr6eLnQ6daZSJAmW
6HNGj5KEdxmRsp15NSQWfOyzQ2QZ/VpeNY8g1zgcptlrLvI5xSUzjhpibkvyngGQzaWRcObCMznq
avI10+eVC7kAIsOF+2AKxOUlbN2W5lrKXOua67mFecz48ijExj5Qxn1adlTK3qVI5tPCgZFMZ1CO
BCFK7MptxxLvYpqmm3c4XcbKePICddRZ8lqEn/13i1BkrO0bsDdKsYZrTcMN65MBVazPDyWWVqfb
mHTonsZYyQoPtZuR12sOfkFJq5VFC3tOGSiOQ5VBcLShC8dDLbBOS+rQkU1tREwknhvockKzX0xs
IHqR/L9BhPeqPRNFrDZUa7NZmR2ea2VsILnBY5l6lmXlKi8ths0/EAJGSS7leWRAKZ8NDsO94W3s
xXK5giUKvtxYwVl7iq42XzAJcbw4NklDsFxcCdzXVPcHjNmvAZE1q1aIBG/MNcwRIx4SyDpTgTDd
CN/jgACfFPDYvwk0UoWQn7jVWFVuodfz7PPcaxCisAKKvWr3QRRC+Yzd0tFKwdjEXuwv76QOSmcA
GCX9kJARnrERNcZgvQz0xUtD5DhuIIBW7aoeTC8BLszj7dBUk5nnOlYRN0Z+8M+bsNgeNPrk6qTX
aAfN6Qs7rVCRq8UCUjgLt2P9CqV64LtVK81FvEOeWaa/brKZk1qkAQqzXtu55SeN/iN/Ymf+Ix90
jXMDMBM/CBDKokX552w8BSVNVp/agc6DtVSzLiU4K/Nw4N140THYeb6yNtdAwHcz7sAfifhrUIgs
dYliKXead2NSo270quW/mPpT3b7ydfXZoaIzIQ1T1cRGrrRmmz4uUkEDK2T0gtqVFRcxmVoihs6A
85tZzLDe92M/lgndlQsFcKnUA/Ntfcov1N8rsoGinw91V+RTTsDZq6Mv//tlGqzRojs5wti5rJL0
hI+tFplDz4WyYZx46XHW2MecSbvlPmdPThM/h9jPJnAOn84VruyR5NdoBUe7Eom3VMUsjBZWDu/u
24iuOi4m99OdGAAfiMdb2B7hmZ73M07dYXUrk8BQn0lfswmN4nbMAAMjtYtAFXho7dyOr2ARAnkW
OelfNtEIkoFtUf6Bk9j3iaRnATIyHsnE+EG1XvQY2+TYBLDBFpSHMQo/RTNX17gJkEZyDUhhBY2h
d9h4BuUchBKpNeR1IG3N/OngUWn9/1pHSyNxa6Z5xM+ERejlP3TqvsZ8XEo8IfGqhV+sqIXg3azP
6PSs9fI3Zw0xczy7Vs5WG4Yz5dK6C+Rj3ktKf+cHYudMBseBDxqaxIkv/qIfcSp7nc6JLykZ6I9n
7AjMM0tV9JthWcBpUBcFxTT8uSf5QIYxIrDE7GYoobyVSr2rR679d3TuolVuLh+FHr8wNDXpHcSX
5M3y6z3VqiuPuUeVOTRTLlvgtYcFNHtMgP8jMjXMb3m3iKE4H6znG3SDdRhBK4BazhdQVFKCYAsa
gTjUvSAhvy2jn7u/AFp842DlSAPujKO/qheE2zgITL8HRF8d/XIR4RooCJGWOCS2uR5NXrjkQd9Y
eJNlCcAMloVh8pSQMfYU/ngzAoruVKCHf94ld7DU6EANoAxlu7pYf3rgXRZeyYhlwpYgtHJ7VesO
9G8pKriOZFJ7Xrr9+HVO0nsllzw/SF7bYf7AXVURnTHZl1WCdYQdENGTqziljccsECaXAl/ZxJnR
TIsYxQ2d+MAbm5DOEDHmQkdLxoIjYJzLvWhD+zfTAmVhjZlqJC16VD4nX3URcUAShkc1ns9+36z8
uBEQBopYZTAb/tDYoWUeqV9FKYYzGuYHG2Pnljiq5FngC9ngq75MGuGtmSiPnJN4ntxPt9xkMOt9
ocgn2kAPAxhmqP6ofE3556DMKYzFezz+zMfEaHvNj2b7gyXJnwT2HZ+1pK2sz3CV48PhGkhIOXWF
7bF4bGkaUEb8o53TjlKV9Z9klX5p99CN+sEI2Ot2N98j7+QXdE8El9LG8fBtNEDUDv8+CfT9F/W1
Gksl90l08h26gS7j6G1OKQS5Z80P8Cu4r1GGCXyWnXxgOjUT/3nH9ejkK/2aj1ygCPWINatqHZAS
n2QBzggOxjcp2WVbbUuJkRbRt22HNaGfW0ltc/hpC9S/cFE/w97TK7kcViTzZt1u9FJkx/TqORj0
k1KeMbzrttY9NjjEnXd0fgopwOsn/1EzFIAHQEfL/DBLsrjAJigyzTn/pSnoK/3wviGxqSNf6Eao
wIUsQVhHvzgIre6z85vhTHF3n4tIN5aE7T3Sg2TAM2JFXFCoAr/ALpzXKbQHPpzszNYsiM3k+tsc
AIZqipaxkmfu4KWMCAJN8yfuhkjhNGKW73qQ4M7/VWxdLBl9ojDeul9THnaqEA7tevJQ0ezuZncy
u6fhRq35TChZxX6oIUkVGG1AQkk28F6cB1fb5TluEOrRMJMx8/eIQbaezGkcB6fkJg5Y860JWjEq
CMXZHh70qg+3H4b+fGuSbO5JCrpP0R6fM6QbCIHPBXWNRbDa9s7/qkTShd9JyzfmfeARZ8cJXh5V
bWFhZQEbT+ew3l1iw7ffKcEfzFHFKU+SF/9MlBkuw2fF4+nh+Vz5X3QvowVs5ZZywU+8lJumqcn6
o3BybTv+JWoqR2sjV8nAuKYHHKzmOfoEJt3au1kSSyRkg1QGVf+ErBksBhnMopoETiwgNvKGBLxc
hz59jKHcThET6orCGclHwjvJsVqnb6XInw4MLsO671oh+MXWMtnLbYlPHbDnyyjeMATY2LnXEr/n
c/gTQCKB8VAS/6AdGdSj5KUt/87R8O9tPyt8mvSbggFsy7GXyEzXzSPuBi4UdbZEFoYiDcx/UOt2
4RM5+ZYa/z6SlnbCVpRuhbY4MDnV5TwF+Fz5veQwmOfeVxEjqRnP5mZ+1ORjdlEwOVVR+SQkf3dX
56SgUwv1f6v+s/00SMcBBRNb6indqnkzmwctZwaPkL6dlZZubEEKaa27H9rfgqSX/KW5CP6r35Bo
lahMXgfsLA/lDonWi1Wt5DQE+4eYBnX26ImIJ4lS1TyDz/pWxmtbDZbfHnFRVSMhPMI0Y8yByQF6
i0gf0icZqky2bV4EoGQ0I/tZ2U8sjF6pa7nT6tTPOYENkllFL3nS4EutxGHSdbABsZXPALixd+Y+
ovkMuTOXCsiDqNmxzSGtoTKjIGTcK2oZ2Z858GZ9wN9RrA27ALWlWyOtRJL49mbnUlmsf/dupB/a
+gzVEum4t3Ka4dXBR/Dis2uvGmHHKKR6tWGXStA5J4KLrFoQdVteuW/7YF/i2Ush/WY7FoyXbod0
quK2OTw9jGs91lXdqZdPceqAxAIqE0FyAzKzD4lgIgCWExabim/j/rccKp4Icsk6nYk3wZHhs0Ka
247+JugXsRblCty3aXs1/B72iBKqRxiWKu49rqtW+cDVJhVp+h5lk6aDqxrtcX2H6LLCJreEV3lc
G8S7EOVJOsFOjMA9ZVycInC66nGMAWCqYo57259qL3wBHhSSdnFtY1gsr1n7VtA4PuYOtXNipeqh
Tl4NqOfrYjbbI8XUSQX1aycbtgWIqAeSwrNB4SghSHmgNtIEmvxIy9U+rToTk7cX1yzGr18kShPd
71f1xWpUNdFfqoYG50RfdpLojV0tpV9PVoLxpXwVS/34SY8DaPtPtPteqHqLtZo/UMMGV14hrsuL
J/XdwmQML5SQvKAHDMZNSd/8Og43kbhbj3nd7SalurMvW2USSSGZ7KUlg9igPlq0O19mJYa6IW+S
4NjlTOezQ31tHAx7POMhcYFg2k92ZbSao6BIGDWazeXbzFG7fK+wLREY9XIQDqlh72jD4bQFzan4
NHS5+w4guzT/enKMoAKxmTmubg3rOjQAKeiNP0Zrub76tDqNy8yVu4/tSgKB3gfRA6ML12Gdt9Uv
epmq/blKQkSYfS6mdOWaFaeaV9VaGxOb8KiQU45Dvcrf0Png4sUhr1N/4u7kPkDM4RNqlNnOqdSA
2yZ4sjdUc+He2lLJnW227o7rN4529cHFnWADCRrRpqNzGHu4vN/MiLiM/3vhRauyop2MqcX0MHu5
4N7YsKr32h/COD4MfvCfuLuoyhYBkrrnFOyxIlYldx6F9l1ECqFstFsqlJLs33d/OOQw8B0t+V1/
ghUmf4M9q1/BF/yPQq/Q0OLAr+WhbZ69NSLmRCRinbGHt782TRbGUNt5KgIf9yczAX7XuO+tz1t7
xwSkX7skp80piclR94LhsoASteVEqGGbll2tG1Xt+am+22pU/9775Bq3gOfMHmB7nWfWfdT1P754
rag3DELQp1xkzEvZBw0aR5M4786EX1WJujF87SCLJR/FKKRu3V6AqP3qN6zWM4wIfRpyxtj17ZE3
lSUg7pQba131wNqF9qypxUY5rRa9X6MEs/0sMAhJTD9MerJO7jwUPMpw6Sd//KVTATN4SxMqoA+h
T1391jK4dxoxrPNF6X45QHUNOpdX0h61anMCzx63mfAFF/X4Is9fqlFPq5+0Q78hp2zUHTLqIynM
blUVo46aMxN9RupL2IQtT9mpFjy+NvsjFpnb4eImsyCl8BJBnMOXbdh2Wf2pAmtikquF2JxVQbHm
MS2C+d2NSMr28U4ZjKlA6ACxV0OFYiwRqrgHiVdbosAq3RO5h06h0gN9D55EFzK9yHo8P5vqXR/t
EvIB5lkJ1olJEXwiwBNl+1MZhPOogINt5oRmxbdLi6afsOh97c8MnSpcCy2DhfWslbEBILphwlTD
d4fiKNAMzlUWEz4IamOV7pT0h0YjXU009Cz/LGADOWkK/v4W8eA9NsoeBL24gYDG81WeDbEEyX/q
5wKnSH1HHy/G/67DFKfNVFL56DiWDTegJiC9Xmap5pu+5WJ6NxXxNvy64bCiJFeB8+DFq6Q/XWIN
2pkN/D1/NUwVA6sDEVOLt3RIZBK9O5NWqwdnLMFBPLpk4uwSz4M7JP6+4OfgeaHadD8B2ONTEREl
ZFqv9D6CFnmWlNZxbCwqj96XsJDpsqysEMGa5cPCF0EK1ou94wBN++QxFj8l9d2G3Mw8uv59Fmzf
FxOMVJcHjX5YWZyCb8KGqOtLfSr2HsSwh7zqbeSYofQTyKeOPhT3rUG+/vWbeOBpCvzlc7WZMaHW
y7qZyYa/HV0S34iZGtAaqJqJBBakhJ1iuDwNX7WvzqMpRZvGtAFQ5+7rw+T+MlsZMPPfoAcaFRFx
9ORP/T7C9hCmZ/kcDYeSmNTH3rgtecoNjzGqWgTvUd2GoMOmtR0PwnB0knZOJ7JIXTEG+mlUFfpu
y2KnEFM/BCECshF+xye3q7+avJ58IhqcMQTE96jvSYdmwktX0MMal+WTvubARcE2dAIFIuzxFd6M
gUYavDkHmQcqXzgtJgYbUM+dtj1tzmE408hY5TNHqykGV41D6Sa6xcoQNnZPTpNgYhuCT5GeBSK2
e2RcLIH0/sak0B/XQ+q2RYojhrPhOiuDeq8H3SA5vFQT8xFkO4xiwu4gZogfH7ENPT8fH49C0DiD
OWxEo0pmZwJhG/Q5fJYjCOgOB9OjwuS34WWUkMkt/3Z0EPzgeWUMpLzP1Hj7BI2J+tx8G59wp2DD
GOLs/JeIcUFwbrGsf0sJERXYiEF5RcHnbmVFvYEsMVdqbKztQUVNOqOT1dLSfZEYj5xAn29NLotT
mNHJ+YANuhuCSP3OPZHZ/I1qEsPKHtmOIdZb2+wMGVwSVMhpuIQw6Q/ii8swphzdoBZyDRt+VJUY
86kjS8ZVXKygaGWlOY/4GmWXgkkLTgNFibZgDL9xBHkKhRLU1XcTFdaDqKZhabq75z7ahJKtLnQO
W8vNoDbuC+a6e7oldZibaD62jfahu11gI3RJSl23EL2spjjhI3/ZIDlnLNGwivlmyh+r1O9vzqJ1
gTEXyDejO2GYedSbnnUOQK2OzWdy09jSQ48Fq44K0Jh5zIlE0D16F27LT4IoZLZExJfQE9J3I+iV
2Wpvi15fQgdFWt3SlQIVDFymxmukFZPJSA5m4HL9FDrxJbtlWPcieuXT64VltyMrkNNjN/gUHzG4
XJKYPuKkCfcgGMBml5+WjKUbqxuvTkeD6u2vtWT/3i5Aq0THzEmfHbdou/zkCeONmiXjD0TWVNET
7UwZZFGV3jVqgu1e66Wf6XgABE78FbPLSM3TCQ3Cny5gtpbqRkIVOpVj9cdcRBA20Z+uAMe0JQLU
f0cGgMHgMeZCd1UDBw3GJ0ePfLsXMpKBMUGJKwkdocpGNSkbSVAi5Bb4T7ltJINkavaVKdMdPXaK
4gdEleSMH7r3mNZUOmol8o8F/UzcV0zM+aWHykwR0MJotqN9Xj+eXx0/u0GhgNDxyN5RrAS/4QP8
QNqkCrAkIrbA6s+OxWBgJDd36cNMbzqnTg93ne9/QYFZxumtXr2NMOTagKvRY/t15+AgoMdoMoCk
7SNS7aS8Vyf7yfjHqchteG2ITDzbUCZe5R0bVxxvhxbudJQUdaceZM6HiTVlUTy180ALzEJXcOQf
XVC6/uqmwsC7DXvh6XnAEKJ7P1cqseZ2Qfalt4J+rZ9lmxcWKevS8o1yaDaM2waoNTGvDDXJP+lj
b6KHCAV1LX4z9GLHqL85dmhUOIm3h7eJNNA7ww3qWhnuiCLmby0cn+J4LmYPmF3lCWBE+sZRTVas
f52cRbcqU7DtvDmDmBdtYc6tfHjBMxf6XinOpNRoOatejG6+9G8dsD9UEzvvA5MlypERKchYWL+s
jyeWPvCH7Zh6OjMRHSud/8Wb/MCxgs9qjo/c1y0dlztJdjV3kifuzoY9M2+QpRJqSWFPEg0w9Bvy
bMG+A85acryHk+uMnv1/pTTOLmc/WTxYcox+SaJfi9RoDkuRaACszYYQk5x0Upt5tV1h/49sZH7H
QA16VSzpwxlmeyscETgnBDSHgRWwLiGPDK/VxelRZSQ0aW41yo9QDunpTBxF/Pklg7QcVa+yjVbH
lf0Go04rvMKFJkwCyhFKTu045NwB43UyA+GNFxiDpkHqzAkFAVZa9C/MNdlueAJKR++2sYPlO7cg
1F3Ro5YILqQyab07rFDJXqEk6M/hd+p0rRb+R1cIqSyR+YuS6ffQKA4PIDmSUqUEaRw60JUD8JLs
LbGkUyPMLBIvM38VVtKk5/ywVKLO/CwOU311iDB1vLtDrOr0Txsd9fPvEPg83mP6pgEapf3EaRYW
wsJqy+3njkRzCoxh6IfKlhz3CYLJd3QxyEQlPRDg4uo/2ui08mGfpEsqbIIjApmokewOzWpX8RwG
UYC+QUGTszckUblK+3nX1Q95Nl4QCxiF8wiNy6AYsvihAGI5qczx2siwHA8sr+MeG/Hx57xvaqm9
QnCC0YJTlf3BNmXugW4TDb3PfotRlmNixvJ76xBXuw25Oi09VsqiPai7rPyxA5xYrMuXh0c72IJS
XqKk27Ote765mv2YYOCmvfkVPWnv6TgnX75U9l/U3unAeXS+qnIrr8n7JOTqteSLVfTHaPNgxgTD
l/RK/OL520BhGGYzup3kMJPGoqVUMC9yJC6Iw+Znlm7NQVPkRCHZmdhUwBv7AalgbldmFfYgRLjF
KOYEo6pOeeDTv/3D1tldaAP36FMI+Lo32yJf9BEnq7TX0QQ5PR5DclDZjWxHKGBzOMSQ9F6NKb88
rChYFIrERN+XDtmJXat2gEvIQVYyTgczVV7IJINHwuuoK0hVBCjTEqfUTKtPQiOt38gjvJe6X3Z3
qD4Wc4/XM7DaWroTH+31cJBioNLUjCDT3leRgTlqJno5NeOpxmWEel/sR8kH0pRwRJtI32ZVdYK6
BfDF1xKM4A1db8c7/5OTDLPgnSa3Va0hCZ9KTLXKkUIvMvGaO8Xyy0M+msM7//O6vw2zE8kpEg6J
8N8jKp+YQNb9yS1a0HXvjvVqVmcRq+18lntoddnHaE6P5Kl7QLRvPUtAYeQxu34/XWLHx9RbgOFz
QwsfWLZupRKFkvMKFAGV4+p25svk0l/8TqieGYDN1JpvWNS/6lloQcAQGRHtfgXi57qBxlStR8wH
YgMDEysupiwNjlnJ4g+4SUY4dHW3zv9809Z1NyYru4UJbpV9a1NrrfJfO7+5Bq4BxZb8GxAnDQhM
YZdHG7Fn9DSRj8s/AEZALhv+3WC5s9/DNgFoeSeuB5CndoDTAR7ROMaEVRMpvwM8R2x/0BlrHzsD
hEzzDYunhKanOw98IafMGnpBpybDgSZfb+YJN37+4Ka31egJDibYqCxeD8rPRmXthUfPv2oGWJi5
pfmZLw7mJadK0VE3hif2N3WF5J3VamSWwPoMjFwbG2Dik7KgNh0jKNPaEogeayZgJC65L+gbxzz2
nwQRIOV2mVO0Zma9pGEWL/0gLVVUUJSzObx5lIZcilL2aeyD/ILTSh1wgOMPDl9YS7Zafu28BpHE
z/DL2Fjap56z5Wab7uWJCKVWi5RIgvY/9KC0RfKZf/tHdeyJ2QP6ZSvkLgMptiVw/F4dhWJBzhKk
wWiO0X8Me87qHJa9IenT36P85Ajn1PpYX9UVbZ1xQsUjFDKQqg7OQ+KE8wRJk2bFoodMWizcK337
ZWPSHZKaAwNAhS8M8kCrqvlsQLRvRgEu2AVJWoZep5ClBuAClhgACw7XlgjGMwrsm6xb+VgHc9kF
e3oKW53IrxF2QxvQcB98dg9ZLBhLvZmYCWQNvo7kSHzpdDa3sU6oD0Y4EgBVuROh4aVo4jSsnnTw
mdVlwQjcPGBhaToVyWjhWOFSzR5Xm+KpS4e7eYvMH4l1E3f/Vc18bUTmdqvOBpSGJNNxcM4vKMJN
6yOlqSY0QpuGG2mme6XuTDzSc0fMaJ16C0voxdxgYFpU27xb+UP4elITthKNFnCsgjylgRO8R0Hs
NI0Rfy+L1a4+12zzrH+Ur0/3lFPnfppnDBeGd6JVpnkHCOD4C/A+WFu+dwHM/g3uU+6wQGEEq1cB
pbMSTV/SdwklGTkgfGkGI6YNBVrwL9UxCpOKetCgBTSKTa5SAgM+IPk6m/jR3sROOphcCMSRFlBy
s+hEATWPLL5nYpJOKET2cYSdtvCAAWyYvZ1fp91jS6kBJRNxhgudLp6FGFuGjZXOMIfyoIatJZUX
cvxyZ3FPVci0cZ7wA4G5vQpfXhWmcWb0pYucoyWqoxNjq4qXhBit2/tzejl+enXPC9skrL9gQzkh
o+1Dsa+UM3NnDlIWkNuzRtMuvnDOINxzb3D3livS04MxoxNHy5sLFuaYdw3zGng46APrmzrtMG6G
N4Z/VD6YWCJHAw/fq912VF9/yDFt2GsyXiBYiKq/mL2Y8ySCl2moNwKsaxTzxxWcja9+JYgiYEB9
egU6G43aafrcd2wJGr//yvGbsLX1t4BNjPIsi6gQ26JmCiLTQ7rGhKaYtHafmdNg8OB9FC9zYwY7
SUXNJz11r8yQf7wGa+z8fP+oTy3HpkDCcyW9RqdjygmvLYeT0TJmEBQHFqdKVUHDXNXDw6PAwJKy
oGISQoQuhbTbWFA3J2WnkaV8yHDd1wxbJzJOba+8iXJbW2RnoJjelK86DIHg9jtV7G7Hj9zjKwLQ
BIwyZEPsbPTT7r9kW9w7BLLzglUp4b0Ddvm3eXi67MzgOKuaZnTnPbPGzdjLoUt6T0x4xs1cG4W9
dmfQfk+bNxcPvQI0oP7iEIf6v5iMyLzZC1kmomtrlH+N8dXrP29zo/CIy5WSUUcl3Fsv0YgdgO/8
GWMTqfkAUMLcC3W/+VyK7j6rTobbAhMunYOjgVp7zciuJ3xfL8CFmndGlJmRM2s8s6SGbbjsNqFM
lCDOr7PXmuZfIy2tcbLXqupGRpKigpiUk4CE3FOq7CA1+TLLGqjHa5OpAzSSPT5hdhTAqRfpZxZx
a3AvAS0/cZ4dqLCEHvQ9zxKORbh2+qgDOcfsitRlHt498/9GpcbUmCW7+VwK1VkpBjga9GPNix3U
qTJLGaDkqD62sKsT/cKu0xFeZ2lv43ojnWyJ8IEEa5pqsW7faSoEeHxcGiVPPzmWmGqdRn4H5IhN
oVt+jCux6ys3W533+XLW1F0mXtPy56IEyynlafjuWrHFk+0b7PeQv3RG+Gr1MGDDqMFPwM88eO0i
aDp4a3SYeHGQgVt7efYPO4qo/weRA0zUZ2LWaOoxWZ0tB7FvkF83vhDl8c/zTE89YrWRSEh6sXLC
Z8QPr7vVfOC6hsEBOCgq3mKgiqweVVBj6UopwycMnUSJ6rU472ua1bwY1GcPoGW0LwglakjaizBy
NCCIdWUYCkmYLGd1+xWhTkvS/ofAQ0cPp3TmcdW9losjRF5hNUe5bgZJpql3qOM9sZkQgnTv40xb
NkB05PSqYL2kuvHNdH9AR0qB9vwBe+53tDe5t/Gv3DiFikwDL3Fjl7Hmm++lkYOZJIPelYVaeB10
UXgyGbdQKwuFAeT6nhZ6lp8g8RSns6EtE/kkQH6j/Ba3wU+QzdboOVJzRNte04Y9mxA6fpkR5zMW
jOC4NSqC96Dq54XhnHnG0Gpi9lgpCK5W5FUwAexwgwtP5ZrdnButLjJWTYkNuev3t4j2Ik7hSHS7
lYt+1amfsm1i0hgLx4eS1ICKMI7nSU1hM7Nig3+vp8ZbjB6EpMFcOeVptod7PFlnBVFyDyHw+U/B
OwBGleWxjbOCpzJNCuRbOvJC80+JTrSV5Q17wBgPBY2FdeKX9ewjkSAwJUEV/sSGvANFkABzkVNA
W8GOA+bHCWNZfroQBHgxqNBn1ncr6L24kRu4gFbB0Mpu2GNwPumnyxpLhk91pE7ppWzWGZuTVW48
c+0vhwejs2rww+eBh9eB0o2RK+T209A1gp6qRLlvZIehsE/lbQ+XF21+dFWIfqF+DS9swgvtyu5n
AWdS5bywtBdQJ6OmsgAGyDtUI2ecfS3tprBdChn8w56GuD4czD7q7JCgmh48gvCUQX8nq2mpH10s
dagOha1kESCw3SxTT7LEAEdiRDKyyK65kkt1ciKl85EJrmWX2SX4+YLO/JbaUpdcM0/E1fm70DoY
VfgQVIMR1Z1vfHQfRMTfwQtFUaRR1Ds8pmgUl7d7sDuBcD5+J3XUCdQBHcZ0nmmvbjk7Ytxy2RZ6
xWI0PHrZwSTrb8D8PXbcs0bLiiCUo0lU1RY52QcqUtQGGUTowbx1h0t3qSigxglQi23/37TxBCbh
oiwttZN6/pO664OIloHUX3RY6Pc/pQUSu0I0xexFQmyX2CdiUNDhuR6fdN8WClxP11hIAEOGRzmI
HpVhIIVrZZbrqoSXXP2iMEXcQtLOdvkCwDFor0r23U0GoRxruWpOt379nDve4xZASrYk5GTmD05M
9xYM5c+g0ODWW90ncheIM2QJQoa/jOm0MbBw6Ifokb6jAjGW7gtsuQJ6ZDwqTeHX/fL8wL7l1JZw
saUAMs+o8LRs6gIfLGM1zLJrOy0Xx8mvAZAOIqO/kkgNSl3QuqA2+z6O0+9S6PdPevGrYk4FTbNz
Xc/4jtIP75Ogk4y96kiTpeeQYLVRKxGxyHffVtayPdvxbBYX1+l8VeTnGeZ8YKQuFcxjBt2GS6yD
4b7eUre/t63eZGvxCXPcUQreCvOaAN5OnDgPL5k/+Zl8XY3HgnnNdZDWiWrRTDHN8Cysrli9Hd4s
1jxi7bQ8j8dTzT5E3KIR4PixunlGDHwCIMFX7/c+5MhcAnRrghUo4w3rW+qQQJWF+HabI155C4Av
U2QvOoB7uW9MNl9Ty4rbjeLZWemLtFbW1k9QaOqX11lPOunUH+5Y6OyHzPoYnVL+V+DVC5NG/8EM
4YuANL0tF1ZFMRmU7PcRnbAYVddMbRCwr3mNx9Ce4alfAhesXhmmKyyhD71YkLRAAacuojp8hJd4
v7MmQkdEzZopp77GvhVsyN/h9QWtdj+tQTMG9bUuTex3Ve59fpLQFxrqPhBof1dgXnJVC1BTMr7c
f/bE9WbV/4vcQWoJNlldAuQE8sLdn3meVnrQguv1yf9yk10q/v8dZXnopWpcMIDs1gFrd9rw9nXW
uurrDl0zqp7IGF58PEjOJxaHcYUWT1MllQkE8i4AIo9pypirCFbewkIeVDHAxZOZTYvn2yzpyMSo
3Eky8vXVmx0IwRo9IyuyHNARKfqic/cvjZ3G4FArwToQfEYPgrOf2zztDdqsTBls7cSR5yZ216BR
STJ7Kzhs16S7v7CMdI6gSK0Ykkb8KRiabkSEEDZQaAjXVQlqSQaIFMJCmWCvG6uVkO0p8iiJhe8z
Yj+su6xhpJUNhjOXHNvMcEQF25BjIORbMKCqX3WR7KsWy9ZJAQlfLxa3N5EOXmXC9fzafO7zz7sK
snBmLUQEnUT0cQgC2WKI/hEr07zNygNQfn0MgB1/uMrgl5qCBPcwXNAv9MRNhHIo2eoyWQS6k5z7
tWTsS6OXpAVHZOS8Wt1sdRUiq6Cc0CWb5J8hRI1o9m1P0nW/L6OZjgAvg+dgfQqrrVXm8BHUFXBZ
kd3rPW9oRDvInGSjgxHIeSC1HPZG9B7AOitoIeELNQGQR64DH4NNFk9b3uZ3Wih/MliSB1Bb00Rg
AdIu/uxKi4FNmj3I53PIAMjNn8toRYzyqnNs07JDsSqKZK+rf0lrmbyo1Y6TtIz47sOrkiJhN0eX
e9+4ATKSGiSuGxHpMPhjo6VEtMhaSmr9H2nNgWSuK87fC2inu6OFnt7lHJKXzKcyzjV1UOREm38G
zKaO4u34NJNzFs/nnDs1gEEwMWm4hvETVyazUtvtbEnqbaVtJAq0QTU5gP3ctilG+oAciLO/Fhi+
OgoHRTnnZIBuonbZpMQh1ujLMj93bIFPwOED62Qt9Ek26dgccS7N38PN/7po0RwSH/go26HX8Fek
ikbhHPHzuCRDlVdq6vh8xA4XctaiA1K8w8fo17E8TJ0iQh2oqqP2ZYPllkD+/LpeGGUkuOUrw4pb
1N2mEHu62/wOblbJzRS8wTLuofRDTbAAS8iQt5/FIXKUH+bTRF9KmN+yvD0W5LMQYUQE9feAv7Wt
I2V77134AlTNHB+JJbcCGEOcmjE3nVPJBbs+VlvfloHlrWWQC7g5JlwZjMsPZ15AAqwaWZR/KqvV
6kHdR0UnqDQEL4spJ83559eq/B8Qf+37YyF/aiHxYkGr9GRrJ+3aCUmPg/NSJqkLBEoxCKFh+7aW
vPtkKJ5Lv14KNW0G4COABJeGXDcgazHja8u4i5mUfpUkYOULwi000plqC/FDBVy5x5JvdWIMFBdp
eIE7Js755dsL10oou3hBBrbyjs1CjYB/hpCQt1Q2GEcMxBIAIlihClOQqfS9gBFfFlI/TfK8P+Z1
tnzM+mBN38S1kMU+h91wjqzYq32dZyE21M5O7bQ2BhV5nYMz/cuw1JX6VfMkJ4Q8KuOoF6Gi01tE
cGw9UuNc3ZI7BZSqcY/eMxjdDFq162Mvf4rzRl3CHuCPGFDbbtxWZeyXYrtgcw6/y7wYq5FI15NY
9hNPistVyJuGYb8oVyqcP9Yh/5y50N6pOeJTXoWrz3eP8JZc7bLCubEMoO7w+jN3g+k0d+RIZWhv
kgVXnHEQ+KIW1baeS1UvSkPt1Izqiaso6EFsf4PQBVwcBNeegKmFxN0r0FS5jZN5aNz7dMs3Vi0U
MvivenqRFe6xavDYQYAzLCFqcFF6CFVBXkUlpq20VtbkxgJDlrLKxW5F2ergP7qAnJg8J6yf4ztl
SIROHGjs2kz3zfCab8gEQYtXSZUW94sZ6xM7hJAUsaXsUvFxbNVjq+/pZP4+/BIScXuC1Mcw2vFH
F8AtQ7DpzYOSSVCeTY/o73qgRjBeUjAb/pMNQX3xmBC0+4YF+ZHKYlWyvG9tr8sTRzfmWjuSnuHV
jGDvI9fABP10weFOqFDonQdg2lyo5KG5ETFTN3L2QrKhHsv6ZfCw+iEDBsRA84yWXNJNscscY0eu
2t3ljcpXhBZ4hY75v8x0z0yanjzVbhQms0LhO1efungoqLAmsVIrMYaw7xl202UuKQMq1QzOvOqf
INrCKdR6fG3dwjV21cV8wspHttS/2u+IYRa/Sy0DISImJZ3N4m2zxXTS+VU08iurjJ6zC5s30FSe
SQWEYu7jaNDNw1wpGbb8PksoPfH/qLBbKHJDFrBtLgdYkUhBBf3H2lPAhO0MpOAUp2kf7amfTR+I
RViHLnMHJQVqe6wmCXuZTTcb6QyVLGovrBLtCQrmtvsna/57auvn4S1lTzbv2rU8lUhRJONM5Cpo
xrxRtA+gW49qkarGY0DI02m9EB3OcQMRW6s1OyWd3L/A2KnU4+zbkvJQATj9B66nj2cIRWBtEpaR
JUNJZToy0zWUPpGqcGZrZ8RO7jwCY2M4XG+m8r77NE9O1CuwdZkwYzgI9RBwR75VonUSefhvyABQ
7zuONtNZ/9KdzD/JUOza7658thdB9tYXl3/NGxH7UsQDoQa2FT96NjQv6T8B2/N+Yr60puKtyS2m
WTOOx4zz0uylWLwmqs9UgiVvEr455ECIanMO/VH4YwH57kj1pfNXc6PRkwcM+7Ffb94hF7a4JBUK
Rao7v4cYLJHqlBU0YQkuk1GhiuYUdcSy5PXXavObdzKuNJkvjC/U8HnfRCD+ILTG4+c78KFrwCml
yRAFyp3D0p0iQmNiJJ0QIYVHt9OqgnFexbUkUzJH8zl0EAcFB0UyfLfvXll9rovXyJdsJmfa8DNC
oPDfDaE/MNs6VRZDFsCPRUMkNBm1lL8MrITYiuW5N+aiA/hszReaGkVTkKDxIkJfpkBZL0RnDM9K
da9D4LI5DL+iIKWMgW17tjdLPASVFWvpE6dje/8Sg8Ql2vRP+VJCGqV5CVw2xpkWlIJjcTO2CwSO
MJ+GKK7mcy9wS+yjWZi9f25cxTQNcAEg2OvkE902RtIVFxQm5RX/q6cpX1uTWNd2MSHNlaQncyGD
Kax4Xfx6wMqFI9XbGwxJvFuYwm3O9EyJHS4KLsTCOdZB/m8CutHvgwWOA2+xbb01+MPZa3PYkQVW
oXYAGWgj4h7IwYeP+arumF6lbWo9MighR+BrIP5pNHrA5sX3fpFyR3pLm5Fy76d9hMjCxIrLejkJ
4Wve5WdsLWmaBHAplMHpFnCsw591/979dcP4aB2f9f5DoSPcDrJSsCrdrabXhpBn4BajLYCgxicH
J84Y92/VX9M22EjIU0IpSinhiXDt1A4HSq6qbHbYJ1gnTNgQt3jLTXOULgRaulrfPnMT5qaDZcer
K3vF7/Y1C4ha4q/am1d4N7YRgth5naWPd7GZ2ANRggpoPGdGiZdbNJBX+lqI5stVMs7iUjwcSnkg
V4yy4I/mPO+UfonwGGRdf/5AjlSyOMcs8i3Rsa6iDKXJgpxYBafn8RWCJgYlf+vve3vtLc3MTVqs
1Hxq2h3XqQUiTovQIoucsarb2qaKVzNG28BOexmPF8KhwPrOh9hsvhPRrluiFxA8S5ytVGF2Ls74
IX2e8E5o6PcHPJdVQ5gtSmP4OqYKYZID1oM9kBv8T+hqrUgi5+3gVfvcwwdJyQRhzyBgxBESu7dI
WBvAcV/7Bqd6mVR57WiKZgmsXq1BJU3QuvTxIxV3KvvWOFbafRcKkuxZSuOq/aGDAH19DGyk0Bob
tRCzjyBtVMm3CM44ecDX6oFudMswZlXxuwRaGIToagShUncjn+E92Wajs8TV+dqFKeKZ1wdvAr8f
06j7GRu/qBHSxY7UI74otF2Aeq5mRng+YkQUiXUD0Yq7J9kkHOg76pGWVEfUnXVwalO8KpsfrqUF
x5nJ3r1evm5nWRemVDl4zCnRWgQH9rLIokOZl+dem7nH2EacUCd1/a/oXhlInADmvhz30Xr6KxQE
6XR7dsYyI5RJo1uOlKugG+oVEqmBLc+aHHiBxYOG9yt5l06hFtifiOONyCPv+AIaJ4UfuJxlYHJE
2l5Atrp4eGGzud24F3ukOrhyxPHOAnYzjrymbt35kSB0+YyxoXDqoU1L9qA65HOfiyAPmNVNUmor
kwh9Ucxw5kKQUAqkUpZBQL5cNgx8DC0ANS8CBTaulod8MSlTPjocj/mQTPnXkgeS1e4LOXa4UZwt
PrH5DCIJZeQD7uIPLp28UGTuvzRHbHd4DIVCde5Loi3OmyXZGHsZg/t7bmTdVrlJ+OtcUFt5h+K7
drH7Fng9osGZolldP5PJHmBOsIxh+PIuRMgm5r3mr3Ld8N7QTYx02ZE/KRCT/sb7cnTzkiUT8svs
wqjgektypWgHlw10gzXKZW7fEMEZ1EvkDD2wSF8HYsaHv8+Yo/6E5pSF/B/ezawv2j9Fnp4us8aV
miKrHgaj941jIPFsu2PpTugVkI88OWiD9iy+a8SujesbA/Nr0gBFDzoK9R411pxx2A2O0jx7HY1y
WPWgWrc1spRHl9VvqxCLm7crNjGPOcL5dbTw5ZwVtijXu3LE6R0Tpnhpunam2yGzDrmUcY7s0SEs
OHDuGm2ZdTvfDS6U4tKm3zpPplnERQVU32rvotkit5FcB57Lfo80zhkEI83NDbmq+RE+qliGh/JM
we6dvi6bVomnu7TamfrbzHIttv0YvatlCse5UfppjK2AeZ4874ZqJEKopkkAb06wdUrIsjpme5Vd
VaO7rHMnGjmPKfT4X1X5K/cIpI5Y7ICsrjbgnHD7AeOtGrB3a2NJs6yej+2+TD1fz8n3oO/gfXHt
xNkokWUXQPTpO2+zS03BrVjEDUChlQLQmhzyhI95JB870NMs+MNs4Mb8LodPoGuL3ev8XJnSg45w
X/A4pZvaHRw6x8B/JkHMBZl+GN/VpJpCLQ6f/mbrxbTU75ujYZQdcYK08HpD/+segxNpGYTFI0yQ
YFdMvdmoUI7xcYGpol7a8M3YocGSMcatfPU0cQ8vCmS1tfsworHAMpMnh7ZGQL35yRdDhvlMrBsC
Z2uia7iH0H9GH5h3lrJso4isJGA+/UH9Ddw/SLh0V3IDXzBgWbVS01t2j/CQwa3ux2UHseU1xBx3
RLCfLx5PAODV7MUZNlHhUapqX5yFlnLcqrN/zM1uOaIK/igKw8hAAHSxZqUe8y67F6GZkJffATZv
PkeFGzHTKYMF1qvlw6Pv7w8yfi7c/zpMuo38nhz95tk4UgAOHFB606vpnXiIwbuQ2iNXInqLCM9k
XcqBeRAVGIF85wb/EsTJssQSnsEw1aTLUcXZUgTs0956ETlNFE4I20jINmip/nTpyivM+U8M5a54
aT2ZE2C3HKvHNGN6C2DuFfz4TZ3kHhNCW6r3gaGS2Z+r8JioEHEBn0i2kpbxGXYHCxaqnOmDOJu9
aw5ppWsDlP7i+IbVzRVHXrYq0paaAntDbXGg5UYP5ed0ePEY1IZPVBNgcXHHeWDiAs56/3pNJK4Q
37v9sEtllxJYVASfNhJcKHf+FRxU+PiHPnXxGA1MQxVp4SmBlJ/n1h5u8Bw54WZtEny8O4ywemyQ
yRWR2pkLqglqAoI7n2rWMWTHA5xWmyc9PveQYj3k5sZOYzadFr45/IewP/ZeQrhFbcmLvsxSisSj
Dd9ATIN0ARTbBDhaY5+c6Z6XWt+lMkxNGxRamjaad9XU7cwRG5u5feQUfyifChQqixuKGDpIQ3pm
65vedrlMGO24S4VMIiWhApc0EDOMLX3bHsDqLCV0Od4LXo0yC3K6/ps0aNVflVRdEa1ZV4WkT30D
SMNF4zEFbq0RDy48caPmpRUTC+4OPJ9nqwS3HbIfAqdeNFArS9hBgYycQ84rcuRuIqB7qZW7vs3Z
Ra2FQmMo42LU7Zjj03atvtJoU3TtkkUtGDRt1FfH9c0IfFpwMpvafdPftdCZNrVUMgNWV/Q7ZchJ
pHvuxzhCWn7Zmm/s/MMXAMLVJnnynsZVvrv82FcYfgEO2SqeCanVyCV0uVHZ0xE8igrqqX29UP12
rkBsicZYPeTjBycyK+7/mwoGIUesU10HF/YHfoHb/2Yt+kS926D00x/ymRYhh00ba3JBV5uGxdD+
BZmgnRQ+OEOHeV7JStK1ojH2Y5DnXtJWwgYXbdqv2YT9tPCSEU3Oj3PSu4pOPx32edjwyUbzeWOy
AkNOSYpWyIvThjhpG4WfK6Ict96cOyBfFYo5EobTedW2DG2K/zaT/4o3UQeY20kGLL2NjX9Ewwma
Ek5Iji6mK7pbhciayPM6+9p4bHXZn2fKOjDdP1fcv/c9rPwGIFpXh2Zi1C4jDwjdca1l8e4USBwh
Z8xxw3FU1vqkNvs9hR3JO+pwLHUYbdpqjkvY+lHcRKaCUIU+vq9jhVPIFSZ/31/nDlJ6lGcbbOnv
dzN/6WsdK6G8p5CPa06fI1A6D1rftdpPpZitAS/gCndguMsiHNmy95hTDRr73RUoABFn0uz9IRtl
rdF7NH1vAxzmOJGNsUX/f7VeybJtgc+YjSf+QXaQ0wECRJQ+nF6nD2qwk++2Ymtm1NHSxiEDgHES
v/PDjz88UMOAapGqfGgtazKBmouyzmRSXdWsOxnCpTIg2uoQSgXH3qGxamRFCbF00t29H/2VpSs0
D6RsOdkvOgzUxWoOc2iimfXb05Rke08IkqDJb3d1DlbVEYvoWhpbcJ8OVzyiXRnCm1BLD+ClQFM9
iX8dUnJLNganeNzncKrCaCmjr44oH4V2vmhkvG6aSQCARI7d4uTo63FjpfmKMBUUtlE3oSP5n7Yg
EgVHMjIOaLRydO5504YVr8BMjg3Fiom6ddQwj7/Yn8IunwVD+ghfhlWcfCdvhFL46UkHmX47NpRr
3FzNZxqTfOMU/lNGdPhM6D5XY8QiolU7R45aYyRVPBNHu5gfEtD5BjxYpg71vGfwbAJEQJCZcStG
Evb3LfxtrOBADDeENxG92hTaKt6r5mP7rF7Sf5SHCtlxv37livXP3kwbVui24x7Jql0YttMdps/K
THnQ7S7WKr4kjyK4LgfyjjXFZpUkvZAlca9GO8VkuU/FpiUgdxxZaFvbNPF/s6M9oABpfxM7Rlsa
6nE288YVLT4YHrNHAeDn+keUY6ODuHv6XVBfOh2Mz1U0OwLOJEZp6FyuNkJsiKiiZ6cNkIn07KSM
mVX6F3Vts38sjsX8EJnSpCYZAjJ0Z2K86jAZUqzuF/3mZ/I1YhJC2i49Pinwm2AtxMr/G9GlmaJh
AIyuGO+is+r0+5mFAdJcID8qP3m4f1CXTPr3cAtRIN7IlD8jz6ZOelMmsONrJAvGm1kCzBPWNURU
b5kfxyGvTXbYOCGkz0i7tAWiIkQkSyfoxdMslPabFJK9Fk0nRr6MqE9sV1j2uN4f3HoNEU2OaK4S
gHiBGMOM+J6zhzrrrfi9ufMNYQc4cDN+b5dXKiGMyK6acOYuscPIbo+MMn1LIKQCVUKxylbeMdiC
P3M0hNb02iKJRZn8GX6Bw3qz6VkfWxL8awGWcSmoaSjh+ALlhiCJsOsi3+dlVLHDVSnzu/hS6KOM
LYObGb4qaRG+8waYTeBwO/EFV6kR/vOZIY3PY7V7dJPPi1l3wQeCbepdf6pulEsVzrWsScTcWLlP
1YGTvOo3JwrXdEw+Ob32xPdzIBJsPs9i3adSFI+dhJSQFCy6Gpov7N76RJVktA5g6rjdo9lOmBuh
n25UNxViGQLfcbGT6P3CY/Jh9ZpGxLbrljgfkkhUNH973VL3/bXffeoyRVHRdLB5+yJF9KzWu/I8
RZxxNlhF5kKnHFXVCUnG2qYKtCn4kPbFuOIRKnEiyRVRJEOCx/Y21khG6SbWXf2q1yZHVrF3CzWk
w4nIUStr/i4utzIs3zOIOUarb6C7/0qzn3qBL4xBWsdTbDFp+EXpzwiMmiuKbdhO36a41wbXUh7Z
i3cQG9ySZQVeff1gWUxdtnkcp4ccL1P9ia1XifGwHob/WZ3d4iPDm+ttPB/iFkOFW+zw4dw679JD
3LjLjO1QW/1OOfRo5KyF+Hzd5IVX6zSL9f/KuaCGNlsb3UHNAEjLUZEFMF+jYjwp9bkqmMiuqqd1
vultOtIuN4qaLgPtlzMf3JVfR/LcNQvyxLNDZALfXDNFHKFZiiUULb4RHLMiG5OsEEvEH8ts+1CE
xNUJZErwABQcOsh8u6Y5mc7a1as/3hmzVUpQbTLMPQe62wbBUCTPcTVbGqRIEvHQQOQtC7ZsN626
5JR7V9Yz3VTQjS8ckTwGNtQcbglMNta7t9kpoeqsKMmKZcT+faTCmjpVowu2vi2yaMIFlkFNkvam
4U8OF+eny1aWhEQ7XgUOor5zdt0rYox4hK2z27LDhb8ia/jRpucX+zDPqmfZY/t8S3Js7U1Ym8iq
HfXmaEu0D4T27v8EpvanttDKWtckUInGT2buAERj7PuYA1vsS+WhCft18wCUi9l5jRN4L85Jl7Ed
pfKZT+w21+6j6j6Te73DcPucQh3WuGNL4zaJmYg+tCeXl0MUxaDAepCxHqx4idR3ieRRBW3H0qAl
z21iBYeorN7TWMzJlFCayCf1kR5UtMkV25kW0lgJp7Smq83syZJjM1aoCp2GFmcosEcalw1grGB7
Ya7l+xtExVDrVuX0k4OMwTySBOSMFXBnVM+2sN2sCo715qCd3pXH16HWYAHOvoT2/YXvGBHah8RD
XshSBg4s/iMGHHs2lz1cm6ihvFDg5mZ95iSv7h+NS+pMXr216egZO9MMCQ7OYGdTGvWkCg/9S4ch
DeMG5O+EGHHy17WhQUnj+dukXtUevirH2DMU4a4fqh193kAG/yApd7pxB4upQeZfvDJvjHMeRwu5
gxHGdF1pDhsu22IcYxDydndvnYIRbdGYe0GhJeiUYVooURXy/7+x5WLUODzDAhkCssBJ7n2nVf6o
gDjg8nTjcXCix8BUAmfXOQGikX9s7oWCLbLqnhR6R1KibP/v+FHyCq/ekEEqzBz5Z/Wao3nPE92q
IIKiRjvc4kRhrEPumPxY6C6r0CTS89+MMI3CrvY8Mt4t6honJkovx80FR9aiRATt+Ke1EzYgwT+c
Kf69FHDRO6Wt+ujt5MMw18uOR0PkTm4XLt+FTBWmR3B49NyFyHYW1aorfayCHXPJ3YCxW3QCWG7M
7nueBceNzkb8FZ34880Hb5vSwn4A1bBVfomg7v7pG0Qqqd4eFpBQ993u9YQNG3QM+ZGpToB96siz
YPEvpb0nDi/KLLgiLk/UdWUm4GolEL9hedvfFuS/nOCZ/q0cYpGuNySTLX5Cp2t6QXxhZbzxcy05
yrxBhbLEusPuJLeBBbijErCdFw7mTnaTxovT3UoOgCEBNMDPGkPMG7y9mEKBGNE0bEOlTKEnppdN
vsqAQAGuqgHvbaTKa0p/Y82Pj4ztcXDwkBwYRUNIeTfgG9lCD7dWXqVqq9NmRiLDEiSiJ6fj/Tgs
xWS58+hhE50Dz92TOuL9wyY1QVkBTKWXQ+H98/eDPNwzhjgDDbOf7r//QuH2OrK/97b0f0eAY8Ie
kfF2XowE7/q4oPC69fBERIX1xz4f+r52GShS73F4x+/SuFuZPe888aUNBzkAsGjEVBPHPiAYV5Ci
L3LKxTs5pdkhxLF/LOlhSDTnjA+OubCu+X+Tkh7kNJAoWWsqizHv8BfpQIlthOFKuAWJu0rThamF
Nf/P4WYg3HKsiFKzk2eDpXPOI7MRgZMK0ncr1G7OiDbtf1XguCXGu1CyXf3RbcEeznB0PxpUxPuE
RxOmUnyxLKo42OE+VdQMWEF5J3ErAP/ylyXNCGgdtFZ77c54DQrcQIrHp7gUjBSVL7e1DKe6VsXS
nah7Yi8W3ntxkOLxVFoj4eE2rEh0hsRf0RrumogIo2GZ/qjSAlmnhfLDomOx3BpiXNd3Nmi4sPqc
L+DV3W3tKPhPI+w7GLqdeXrYPW98g2ptto5ZnJrhMLsdiIsFVqGos6Ua38nanCCa2FN77wjSMQrZ
J4zYfiekmK9rphbT0W52rfaMytXYWI289e24PAtZNY82dBm9i5cZ2f/lYlvMJlGEOMrp7s32kUr/
o8x5xvPocQWnFEw6zKGyQydVEj8emQ8PY8HffD6xrvJPvWuq8kQUQ48lEK8dFn2ye6qCxD1eDxB2
FczBD1oePLq55V4i0EnOfO7hC1HDB5ENDQaqz6nOAQah/wI1pIHY1GXrwsmeOX9LjqI9O2ycV9YH
UyE0AjgwD+se9TC81JDLuXDubeLBXiKdx5zj9N8u81L88flUxrkADgzrDnflFTN1k7new882l+5E
QIkKr0ctkKNF9R9O+gVmpzTqvr59O475uvLecs0gQ3ejewWgsZLoriboDl8tQStTh2Fmq5HnQQNI
/yR+9D4UvfXJsXMsQz5xW51In1Lq1uFsT0bBSa7rYji/jhV0/jtmwf+JGeQrqKWWydN+Kx56CbOn
Ez6+yV65TEqwnKLan1N/LKXiv4Zdm4nyg3MhZhvdM6cxtDsa5JOXYpqbfVa7qcK5uc+kt5VhVfgu
CL0U1IFsBNCS1QTbADgt7AppZMZaC5g3t5y2AHwf1Gn1vHM9zAMdQ2wK1OYkEjRAKKwnblC9li3S
TnsaGE/+MLyRBpd06zfZcuAo4SUyTLRYLkJbpVXp7aigapq9oHJsdYkx8iVretTFx6+HSYmWi1oD
REqCI0x2oHYXJMJURwJ5TFJjv7UAaXICYcc1WOu/RDcaupDaDvzrs8FVjLLzNweBwfunK63Lwkfz
HwOJZciJOuemwv7z5GnDAfa/Iy+S+2SGN4La2UkI+0XKT5OqIaW2sm/k35ghCgHyApmGWoZmZHst
uZCfiEACMeNaApc1vnwAOSe6fO+grtA9TeU6kczl6nQNvs1vsVHn0GqCdJYkD+HI1h6ahn7bC9X5
2SQztgoADI7MIEJhh+kSLQZ0suEJIBZFYjD/V/l4rNnfKRqVmumRiqtc4X80Xr8EGt0M7yTKfpef
SHJoT64NkBTNq269694SsOhGpKW6OFs2Jkem218jb91VlXzO29aTZ9Jjhh/pyte8wANYGEZmv3Tg
xv5fUbJSvmEF3oUY/qa8SV3ce6mqwOUIZQqI6707WdW5Zwft6HmNW/eqWtJ/dvDwSabmjZqye0+J
fJJHrgH05u1FsXSGxZwasVLTHpOoUTZmP0sNJCyoiagZ1XafrivkcspWCwSCtdcquxYXpoC8lNEb
VwsOR5KT5usky3yv5S5u7+6stjqhCWC5cQB3VlTnRNE3WUTwu+fkdxhcJQr7dibmIFDAY0OUfV9l
b/3R7aWEdO+t5nZU2y9NotWWbrPSXaHrGUxFCBPtdk5OicKhT2bnwGr8b5N01TgDZ+0zbv2UY2jv
86DhKHvht/T4K14VMqvaWW1uPT8WomgTBFrNaw+bYEp/RGVnL55kKuwckd9KImvjJs6cFtUrL+Ua
q6LYe7CzhZ/Tq7nP9w0ACHsrA667NCkzwo0u/DcXe8nRhySyydD3L6jYdClbHMbN3559NssO8b9E
lFnyI9854jbKD5O4JkssUfzgPfGNX3ZsAAjYUeLMZ7sltmyFJp9+zWku8A3QOiwsJ/jcF/raEe+r
FsmmLCiWcqiuk7YxjpP98cgyvgCOOX1TEtlVAtbzdCjO+gC8TDWaWsV6flE7QU7Bv7H3aafCntrw
egrzCMxPWLJtxJ6etHR44axlkT1BtCKsrN7wHZHJBT/fchfydy5qsF/RKTedyFu0xktgQIrb6ZmV
pKhiNXnz7z6AhruQtiJCojnr5sPyA9rRNaHe1LVJ5/RQ0r69s6COTOnRQ4zDiSi+LPalVAvpqSez
n9FhbeTU0pvFp36dZxMHp0dhkqwcpFs1B6jToi9kb7e3SbvI8Sl0h9cqvrmHSjDopDenh8GaiqvH
tt0OwGy45kk5fr5s91KXovtVjspkN2wkM2qAlMV9iVye3GR1linZDg0SIA1ZoXO4CWIlbW8uPajH
q7Q8+lsGXmUwhtuVpwPiJbeqrWoZUNUJRHA3VrYLBhEzoyG77gHZ+YJ7cCZ6SXeq3wPSDBIwim3S
3vDkREMRcQQq7fho5fndatAt2b32wF7MRFaO/l50HhCyNfV1YStEY3WBCaxCrNnrcgcZ8SNyUKt7
2pweBQ2FgLor/1q/JN6uXr6mODmxLN6yMITWXHj38eatVzINnnKBWebFHIvXAj+omOlLJx8mIJx0
KJh0IUBp3R/5TXq24j06dphmxqIDkdlTHXshuV+6WoCe/ZyPb5oSPky3FdLnDhmTwWJ+NqNQoMyl
EVbfNjX1hJfAianItgSxZZ/l2znJQJPE9ofIVzmP8aEhrJV7h963wNnt/sykJlYmu6s85MpXJt4w
cxg067hbW28QpdNp3shQGumAAv234jn46oBDZ4ldGhuPVrSzFKbGF5LhzfeP6UmTWWHpw4mZxpdF
QbRD1Z1VLZcxAWoOft+2ix0zD20MdceJUcjqE/C5glxBHnpPvNXEsmtwJY3IWJibA4OmQ54rZ9Go
Q6bLKFleOF7NLmT0MfvSJUj04diW0gLSnJ1muDqMAotWDqot5mM9SN0sZySqDzvHhM0CyRFsIjVF
hsgDpKx8+Ek6fGNzPR+Nzrj/hzirJ41VVFkToJHxABrd/nPxmv5rjuIVFIWH+7h16mjRzK7kBZCT
VjC0CJ/NZ+6fGUYuAQ44zFLl+JiEBe9HnmEZbvi2AGkC7z4RE+NR1HaDj2rxMl8nv1vjkZ2FZlB8
A29iRgWIwV6/Vq9Cya2FZc/MdfVrXSv8En7LJYbDWIO/rKfpbZqohJmOEoIcIrKEMqmwx31LC4SY
1/lpFK4AkZBMk/TDfPuYezLxB4lEd2oj6jH05sTefZs8r3utfJ+NppbchaGIn+tErkk+PRqXa+to
yac6/SgziZ3V0edg4chOapecM+5EhNyuvo7Fm+BvpIebl/1e2jywGqJ7V1st3MjZ8AhfYXn+mYDs
8JvmrE+a3jMk9xYRwmrEgtPcH6/EJRy1/NJ0eBTY/aycvdGaDTLzMJoT+5tNCx3nn5x5CnOuR698
tUXvilmfFVJDVPy9m2Q0rFcnnP+xuQfk6tSbK5DYKuAvkyVPPqLsgWVZC9fQDUXl1QvUuX8R4STu
vGlfH0cd7pPJfatqEBO3kdlfCxXlURYUbV/lhsRsfIvY8jDwknSbMJykJsrzPDIwoUAwASm1h/Ky
O1Nyh6u0lqq6HXhWGXFnByht49/mSPZ23+htUMgx1cD1dmkJxoXAMQtZCUsklZ90WdupUS7ISlge
/Bg3lIIuScWnhKhFCFFZGC5BQKY2yV9haZe/iIfse950QJS1IEplS04a5zXt5TX8q+djWMQg0vdk
jLUem16kpAnFwWcaHQZyNgbzbHJSjyyFk+NrgH+E19E5jrdpKUKDk9zwujuDLmecjQKRVUIs+t1B
3nZuLtD8i+arFwAM4YzoCPxcPM7PoJClUjcaNkU3GcMB+1K3oHqttXzYxvidFM84bskYxrgI2kRn
D+EHS/g6YzVUTWt/tCQSOJe80GPchcH7daLGI920H8MvvIMqTMzN64QPJVIpGzxIKkxef8izz5Cc
zC9DFgjvEq852Qdtwy3KbwgR7Hzx+YpDU/VQQjuoPXyuXIV4HQmMQTMvOgxyXx4FJpfkVMfSlm4l
4x9Xe6y047aMnkCrBqet1EsfddrTfFfXoJGeXRu8ksWf250t5wWY9taKMt/0icfYX3a3+3rkdUHM
Nu2iDFUiOKGaBwYJXdi9ZQ9kcaJl8sz3wp+Cx0yqM03H2lZmiCdIRyfUYvIckIGUK2KfYY8PSpY/
yDMbhKluUhCb3rl6yuQtVHGqyObKmYQqcjXWXv5O/yEkAUxmRbEDRwUDXu9GPsk4C6igapkrnR7I
Lz1AwMDj1xUC6VtPBhkZ7DZbWa8PGM+LeNEsHBpangBRcm+VzRvY8p0hTtosw4UHXZHdcXpEBZrY
W5be31GvgFbtWW6ENeNpZgudnpJfSO3br1mnFhd0VnMJTOIekmNN8qoghcpt4z9kG7x5eHOfCiSV
ze714VW/ZgixkLUd72oJbwDfitblAaYe95Epl7wXfwib4oUDQEHR4SxMVxI+mYvCZIljiT4ouwvU
GPNR0ZcKbPRVsQhB2PMmwN3TjtBqIC/J5VlqfYv7UD6DpT4c50hWYWkTDMF07WHS0CLG+DqjQnoo
hByqqWCtF0Z9m7DHyP5dU6Om7rRE9dMnXmLH1GjzLiJu0BB66vWNooo+Ie3TCNtRar/NLFnnlJ7C
kFZo+RO2VLPj4SSmZDsKyx4WmnB472RwqPYAH/Lmv4levmAHAwhT+uT0WthD9c3/oDMOHnzqI7ZA
aSKhH5rWaLZbWAw4UP6dt6fs7dZtIuOzwl6ZGZlntVPmM482avJ9jhP3SDqFL84vRvnaNIlTuvu3
u4ngGzn4PJBEEzM5xDw+6HjjByqu//sNuojJ0OyYY/k/Lu35R4t1/MEssdsA/kzoZp/eqv1WLLRv
lZ57hVyWtVWVGYdBgZnqZ06Fw9Z/oQutJN5Sc/uEgDUiBMPrSI2ni1LyccSYOQ5cTvdlwxNwwRv6
iLodivsf/1X/aBhvO8LrS4Edx/1L1yA4d5pfHDMHVlBMBX74gIecC1uPdYv1Ab5kX/DZKIvSsXPA
iTcHjNwO62Q3htxhpzYeF2Ah422Vojmt10Ug5Hduqu6Ls+9mk87ruNXaFgAlmqrMwxnn1fgTfN70
kEPybt6sDZqCDfFmYhi1eE9H0q59T+IG5+Pc0zAQ67+/OOu2WOC7b/HZhfgbCpofQBUxO/v0szwr
nGqV7dKBh9WDaEXT23fup1DugGA2QiOxW6cP+GfmWvK5a7rgrZi7Q/CtML9aGJbRyBT3Is6+ig7k
+BK8pzPBahFIdROf9+EqrOhRAL7MGpBPjQhywWIYXjuXcxLtwaysUDG46AtEbHHNMJZhizRY7Fay
tz8RgQRYG7PafzQuKoEACbl63397Cs1j2jI9U25qI299ClwN5KKw3Pn7xK2wxKljWH7UejQwvgNw
r0r0Pds09gOke6jYp1GFadr4IQLQFRaJ8ZGVxND2ARHvtNkoqZCZLYSuO8A3xV5J5uta28bKFuBK
cogHCBqEVDEPcFcLvvP7/qajNnZPcv8xBXai0rzhLap2YXG9+W8fyNtw4p+hFG4I+7HrB5ZEhU2A
jbuVNoKm9nNf4kG2YOjmuQAMoqnYUnLkw5mWEkkt0n8Z77l1S1uO/FGVIYfzyHc4RlqwOGxXFc+J
EN/W/yY2ILLGPNy4A/o7hdMj/dtpbkmave1C8BNg7+1NxJ00xhpk7A8gwe29HJ9nPNrFLf1rGakq
BHhvqV5W5us/1hoVfAJNs1WE4q3HE4aBXrQtbv2dB2ZOaV9gY6sEP11xyHe4wvcnzYlgD4rgPaJE
2nruqCvYS+Zif15+KHCIQA82HqYfnKnHS0x4lGb2+B+vOFm+6aJNqh33lx5xGiVMhKRtCPRkvHHK
tonOJazhKzYmnvWPdnnVfKpbcExe70GQIJFi5MJ7JS3aR1s9kcsQ0SomKyZTKVtuqRYzFMjgamGu
0SKjNI3usW06l8wUu66TgV0eexzoeVKKNwm4hyoiq1gjaqmjG/2BUnfJBCzaHTwg0cPR4RQhYXlR
wfhb02ht+cUV3o04moTZH3JDrrmxLa/Cp1e66rBneawv+CKft8C6MFrI6MESbcAwfRkTanwA3BA1
0fOZgZAZNTVyvIBBCJU2kuoTjM9v/+yXxpgwB9zhDm3HNCTICOX2GXhRsDZLVMnmWGasZ6kYqT2k
PHJJK/Bg6cB1Np1K1UpyWOF+XrtIoPg9zzZZOslKRDV1V8zhuck5xUEKkp4kJcf1Duu/cb2tA+ng
kpyuOPz10wC6Cn2/91HcZwVmhpO1xBNCSxf8d+5QB5IV8X3f/gXx+l/r3/Y+6RTjxt1Ik/1JObvX
89WRzskRyqok1b/SVxrbqGMg6mvL8dNxOmBKLn0syv+zU5awkQdSEJVWZYNx1musPpxwTT7ZlS/K
aO89tzNhwYnQCxJj5eEkFYw4URfLe1G6qXvmnygQfI9C+9mo5/zQvylBCevDnlAu4xKlM41EgyCT
eZDxDM52JvbnpoQ8JODsnsiVVgbZl8uuuzuPR14OwoLNQXev61FcWUlbfaGv998KAqeibhIVt4O6
D7QpdwlVWNrk/dqNGTVEGGfY1zVjb3ArP9pTTtooo15J6XXh3aG5uGsBG08h3Jvcq7RIR2+iVKfB
sQEKXCoA6Gqc4YD4K6zuyalK5WyCc0vgtV9P1ITnfzk0Aoi4TD4FDdMSUYI41facdLdP8QhLsSsd
auWxkhEcHabGMaWhYhvXfz9e7bYb54k8P8iBX0OldVhbizGhwkxyCEVHcxFx/AWT/tiVsRr+a0Tm
MOliQ3rav+Mx8ibe00GZ5ajoz6IkdTwyu8fds50SpyRHq0l3UOgOxIJ2tKbDi7+QSBOHUZUfh0oH
+8x+Oa6YUSAux2hNgokfuSawpCy521mJ6y9XVweFyVTQ5ReFX5psGZDp0XYZwNrdcTq0jWIbKE7K
rlSWkNra6YXRN4tWjA/be5kkVUPRjZbWWQR83AG4ANIp+HCguOlOa4eOyL/dC7AJj2fzLfZ9+Bif
MW/mpk4Ooy1c/qJm6s44iqftyPy6qEm0JFwNRZpPhqt0qnpFcdFbX9MDo8L/TR+vl4PlEXGHptov
7cyTMrL/ZiZFaarivFIjnCJPFEATkRMwwi/+71yoD8K9WvwfCodPSZAdAnO7teysF8KRBciNW53o
b21NgXP69i/yt+6oFeWjzq73lv1+xFIDcBnYs9HDgNhF4UlZlpI707vD+E5Gt6lvsM55j5zBLKOW
p6eP6Wr3YS9hz8sklrRBMcmOrFUxUhbLTVCCH2MJZh2lCOPPusmS52wyb2epdvzHjalZJCdngkzu
6NotesTquDNlnZ2ftud6M3lmR0i29NbI5KV7gMaSDjtKxQVXPXGywQNWeyOl9MHfE7faQnTPjbMN
bw29U0wfc0J8nX5sutOcdnjcAVzJObttHigQV2zWw7bZ7iRetLyJq7oz8bDcX/u1LfhzsDPR31dt
k8i1uoaK6DKY03ttBAuBQ1948C4j9EOF2srZP11NIzSUqm4Nob7HKX04CAjdgiNeoW/tBU2TsPzI
vShBCV9LU+w1sEwsdl+0I7P4NEkhl63e15anX4Eg6RITkNMIeloL/X5SgNpP3neTtYM8LFc2e4xr
MMdBgfXQ9oB6JZyPBLh3YFgm2cSZxlwtWVSQhNqgb+sOSyW0ij9VD0SnMiO5rd1A24vzfSpLks0Q
aK4XKcopuKczdSHe/fCI1HleuFjR1CFDuK7vpZx3yrNxetDvxGeWKXQCUOhDV+o6rvOe+GpFoZ8m
zbPVFwHVKQiQnjYBbAXgB/HTIVK7nyNLPBHOaYAjE8RpwDPnyJvHcoY7SZ5WpEOwuFMtDWTuK6bS
6OM56RZ4yM03tafkrCrcNs9Sm6pLXjOUCSTf2qy9FBt0KiMT3bBL6sNAJtiDYk0pff2KrBIXzbCo
JOBTjhALCfhidhcKXpGRPwJfSzwFKCY8PEgRNYVU1AdmNwM57YmX1aKIVSCSU8Kxqy1NaTtakaMy
l/ok0PMIZuDyBEAYrhNwDlohUiDOE3SqK1YZGWyYrHMXin2akF0wsUruKCPTkUzaPO4eDvuFf4gC
AWiS8+1Zk30aA+Dg9u4SRDKoM9HnICkj57UuiFq7hug8idxlEct7krjTG9akIMikRTd+EepA1EqB
GMy2G4jt1lfhvkps3RwFS26JHfaMOmE6EGMZ1WcwFjkD9nEPwvRqI87UJlQLKD+Rb3KDErZKk0Ii
RHartrNtZJJrsTKGyA06jeEkhSW4FSMhQ0vlZbclr8qRqxIIqF8bsSTO2PS0eb1vG9W2fv6MdyWt
ptk5UCXuaqryC94RfFY2Y4W1kU/iADG2gEH9CcpwLQ4hnD8W8CksBf5m1W+z5WwagAHcSIm8WbHZ
0qNzB0NgOUGgd8I9Vg48NcjJX7nwE/mvNWQ/U4VQrserw0MkOF/T2JfBEdwC4vXZ80hNHWLFKiat
bShr25B3sLHblcFFj7KE0+PJASKQGiQuAOSsrsX6/sVGypyRY+7RWQfUgbdACoTfkhxq0S1TfmcQ
PXrsIMNCkmFgXIhsUo/GgXkgvOL8HN8wmkAJtIZji3ABPYOGjIXrCl+EPnbufFyDC3bFU4kmdt+8
OMh6JCwE4TmkpDGR69Bx3V8BYawAgwn++u4ick6SxeGNtG0ezcIP+g/kGNxjdkKyl0WwCa+mqXAT
Cl003DC5adEeA6O8BE5f3gJIir3aRHRtuSTcI6Cb1ZIhikFDmPTddXLSjjYBafQHGjEEyXpbK6ul
KFAxaSy79iy5Z2Y63Y9l0uzE5AcPnpDpFYr3Q+y4hoYne0yeUS9849sSGVfqT7xOt+qghdk3FPu4
vBHgkuT/IgtE4p13UBNtIBZ9g+cGGgjLeg63PqbNF0Cl50jb6xyeOk/pA3ygM3HLuZS4WZ8yWdZs
xbuoe0GH8lkFMpha2ABuutckUZP/gC+AGelEq9DcW47+H8cjyKKGeNs65Z+CmphD9sJmuxdRiJlm
5Yk56R0Qp5XYmwhd/+38VkREC8EggCBer57j5y3EEmSW8jn3UOXhxsrPz1QK9WomtUttD5ptQLN8
lIY3ymyqAD/XS/R8DpNGtztUdEy8nT/uFjK9MLz/OY09P4OGcrUrlKcAUAQYvsOX6eH/Ffm5Ito2
TFZtu9w3Dv+tzCglDYN2Ue3TNDoCM4j5AJmO3amoWc/81iy6Benn4+nEB0QuuLVauHMnj70BTAtq
86KD36oBFIZiuTs+HkGG+laWIwGfnC5OO/ONlILEv+oUcxef8UcOwnXhpauFaILlUgT8DhSq2Onz
qr1hV2zQOtSBqDgpB6RHtSt0pkewNAc+PzsW+2uEltkHRzFR6RD018eqzwuNWRbLn8/toL+w5jlK
D5/70AjkTnWW7V/PTCFcETf692ViBXjx5oZt0unh2PIq7eyV3IQKzKI8cdQbrWOAqJlIovCRpQE7
hlnxj5vwFEVAEleJjma5VibgXcRdGgCJTwMNsExzSEtK/jacaU/WCu+yMdhdcpHSNtpZe60Nxjjs
UhSTqtA9LTKaPa6LXVqlxo6DTnNQnS01XRJwOCUHfNtDbVcUEBe24N+EHBx44D/FWXFje+r9rxJS
E0gWom02bCVufPb+glVsaafYqmra2+CCx2Nvwy7XAA41i5v3fiN14JLOlzPFx7Mlh0IUE0rqpKFH
QSQlI4vVR/qc2kJ1IBRDhC10lMd8mQ6mmGVYqvXhcpyrYWCQT3oh7EzWtSXLbUxcRZf0JbjLVhAg
iDJY4E3GVdrXefMiMHW5GMjOXmnaPpxWeAJnIrSZbOOcwUIRh92uR7uIe9obgZAl8qbF57aTG/o1
HtW3wOIcE5ApW1fpNFAvzuxJgxpWg2TRloPyqupD/6OZ/XUxFKrgAnrosyk1947qpZ2MUdBOOCk5
KpgVGoBXLZRvFGvq/sem9bDm/e3/W+O3r7jmyFIupXV7Mcp5nY8X5UFtPH9zIrjn3WS9lis6bRaQ
4Lt6/a11TFXhOIBeBfjvERjUVhzoSxCqPrq2OhT08OFGiBIaBGb4RQqmqMbzZ3Mf4fTieWt112Dr
iPvpJbR3i+44mb+/B4LjkHFluw2fi9IjiaZdiAo/UE0/vTYrJbqb6i62vML2xL7csiLub95n/Y7c
JBOCEnh/1v7kp9YnjhFujEJFsZjBMAWOMfRN/JAB2h3kpwQwGRGGKrufGYmMtVqKKXDynULZGJN3
RSZi82geaeRlqQql8OYG3XXfyjyLBFy5FsNyEfLAVWwXW8MgFTYtJrpR699BC9NYTxy5gGiubUl4
ubpKx//Lvq2/8vqwJjANWkduU+2LJLtG2KTbBuhmy4fYiIfOs8xkHeAO6xrz/HJs/pFdZF/fw93r
UZWD7ev1bKMqutesQxcv7pNtX38MPul+t7wledtATsgt3XPSTMohq5qoVWmHz+9JNenSz6VYnAeR
30urmoxrrMIw6+G9m+ougIJ0AF29CxdHqFKRWqenkBGQQPBC6g+kI5jh3WyjfDOIWtPJXWLORVaf
UvE05IFjvQ3ZNulMTSbp0Z0oTE+hPQ5eAQTkzavY6pzLm5YNSG5Nw2cGya3RURxgAXDfkLiAwjsq
OGZvyepms9A8axAC7HTmmefTHDv/JoOOW+WJlsJ6UvfCrqzAmsIvmrg5EPSmCzEwMelm4WvHHkNs
AjsQ9CUMBJtjJRhbZ3WJOa6Pp4RqxTrDjZV0ggEMEpeyJl7G9tULGzEjJ57sxK21hNQVGyp0vQAM
BFp5YmpqzxhcsuLZRxLcqLzBQ6HStD84W5fdaPo5VUn2QYeK9qvG9R7oiGZk3sr4Gu7nVhc9F1fo
OFSbzyO1eAqamuuA++9DE1e7UOX4aPp8UNShoc1+sLYxFk4cbYPPLHXR5v/hHTaZj9eFV9mvaQCv
FzsDloJM3z2K3ZAiPzWh+GQQeiNo/HE5HrhP7QR8H7/utSd09QhLPTadQSS/lYBL3z6B3VUmyDQQ
YKVXz5nrN5Yn/XbLm3Bd3u97TgUEyELKlA/F/uNO7yytLuSZXsE2K+FCw/5HTIMLLx0HthNvtpLL
wBEDuK48RPhFD8fIyJeonF4rjZMVH2eJlqusKcBuH3jdvnWeno2SvnCAwfsfGcqlBWhIL7qssxp4
7lQUAgbklY0aeVqJgBqPC/TRQDIRbhxk/RML4fOtCWTw6zraMM7KXhrQq82IK7s1jLcTbqIc+3/L
cq3j+vl+gtrpJxsxT/Yz4ry681t2Ev3COMY3eZfY9Tghc9MUmTARAkNoMsWEvxYyz1S5lXkyXwMs
U/9U1ztgc9zSWbb5w+dN56B0+yI9TPAiT77dHLeh/k/MOXuPTKWUULXzgtiS4iOC9qTdGTUIbVV6
JFHYCLDrBGzSrLICMEuqfV9lG4WqzpnGtS9HW1lfqW+C/IjQOSEl9s5pi8LrWz2anJGO9XqHKKaI
2S5OjJ11e1eOY8hBV6Us0lIAW/p5lRuJDG2V5oYBgrd9YRLWuhraqqwEbGrTjlLQbAx8Ocka7tnw
tswp7x/wzK0qFL0m4rB3xclbH9ZnSToCYXgHtWZAHdufkrq/I9gE3PSrp9R0hLGIU4/IG6iVWiXN
dpQ8+hKB8AGcURZLrQEWr8IY6aehF2W2aZ0Ub9n/sCbw0l/JuPJepvCOlHljjT5zpaWGIYH1ZnIm
5ebz9URnPkxxW5XZKAWmId9MhxXpAds40MBqSO0sOiykp04L3UO/v6hyoGGaDmgBU83reHVslaDz
hkAt905CA7YSmQcwl2DXFcyzjXbamizHWAv3JI2I41XJfj9bJ2dtXti0/dT70WW5cbI9Zm44HSFN
FAvZq8Zg+4g3s9bP3JRtI1LSmJTtSjitbr3U0cLr7FyURgpjCA56Jhgl71tP3S8AmpXzABnYxBKz
gsEqPoVSbdrxM+hg+qon0GitQH8lhjqzJlANmYOcOao+jzYKYV9ZM+NMD5CqJJ5ho5txXDIwgsLP
c5jEKfd9FSn9jxTmPCceRS+5JOqOsrIjbYhJtXmxfQyV3eX1o5uyhlTRI3LfCyKJI3wV4zweFncC
xDsZ1w7xyTtUMD56IwrRKiOU0hZOjan0tiyE+UviZoppiazEKFDKSZC6pYesClgMK98MOnzimb6v
POGx/4zDBHk0xW4E5BAf54ccXZ32tTCWENLfge8DuU7AE+KYq97WGahA9wKKsNNhR15qKRS4RU4m
MAxnImXSHDCvCenaAa1O7gfYS1RxVAJEWS8mUwgK8ZpNEVRzAIZI51TxNJ/xcIPpVO1wfUWvA0qb
glUGbDFRs5QcxQjB1lJ2MJ0OhXPrldkgSSe/3ktSit7DudbKG68mh2kZQ2Lhho2+CAXsN/BLJkBy
DxPzlSmySGkRT6ag3s0+zbBH6XXIzhA+xlv7j9D+OhIDxO6b6NMK0L3inbOTVamQeapLizwv31zc
qTyCE4p171cLHpYusGjCVWhv2sBVHMEoK66LzCVcgQHSXHwWZrvLCdWs75BXo/jRd/6BIgwciCpX
V51yvi4cfIO4fUFI7a4pkBDgfsxFIUWs2QWAdgX06wSs4OhbRMBsCTQYCP7T37C+eDMqPpaRpTtf
WbKFP2dpWoGOHyGU4XpPrg8AIlPI9XfUmnjf3jQewV1BfLQ0mXo0/tleA8bTIeb+QkvHw7akMQym
iOnJde0m9wfvHbQLDCcq5sHnU5VTNwi2T9Vf4mM7oQxVAs1BnKK7NMHFyIrOXwcJrW1MLJU8NDWc
ZHzaF4lR2lyET5ffPyWjgKqRLIj8i5FG9ZhkPvMsApAUgBnJxRGevtEMATqN0vCr5YVo1QdsTU4z
0l7j6PdAxFKkeisSYbBPu9OXx5LIrtef4Xgc3gwmu50SURX2dvvR3VFNytyWYk6WdyPrJP79+RyH
g45dAwa6iGwBoxX/3bXQId7OYXqjUITvUBtmq0BDTkAx0CmHYZefdDaMSdhpONWzBZjDoHv34Lsk
yDVTYLIA7fsS1Ovr8lT64m8AXU55XSx/0WWEScZOEWukfoOpUboKTpbZKmy0wpt+w/PDVMOcCfw8
k1ERDwxmVTzuY/y7p06T1I95Gruraf0vzmpimt85gkRnqGI0Z7HUjAy6HTgdXE+TIBaCWdURFWed
94sVCarDyc2mB/vOVqMBxjIAn/MFUbPErAJVp40kOUBLPxXsVWLW4Ql6YAk9HjzJt0RndtfnKeWD
Dl4EOSb+BDz1yxr7ywaWrsqzwPuHm52/1Q1J7QBT0vmSOBZKVRFbu2W7W+946t+DgPuwfPLmmacm
j+9SImFRJ34KpjEGFXFZqnirqynPY9xpoVFCuOvEjOv8fXc+fssbjnoDRSJT3/69QBnlKbMGQHxc
XMiyZAQ9qIBqCmcUMk0nTXyHOENIBxDW5ekhW/u+Kb7BY8B7Ph1gXmLuDJ/GlYwMVi8tAX/Ykcct
0ysPvDpwnRQRcdzgaYPHC2srEAPdsCs4Cdx3ByQp/DDsY8z43BM539e+6Lmh7JISRb42MmlmzboX
WP3lZotsDbiW/bKXeC9S1MRrMx33iTzDlkUnInEEN8TECXCfEDHCmAK5pcPrJaHBgxWGY9XBC4Nu
0nESdQ3jnrJTd7EUF9wd4jetfmQBQsonJ4/4+ofJu5PNWBwiePejTmHzR2fhmfWR6SRdlKrXTHVj
J0zjlgFDIL9PWHU5AdKM2/nzjE7XXuOS/bjI+3kRq7Xxb6Avb+TMutjE6qpD0t3iaxvsGZ6eeXpN
7KiNEemZRnKoPq/NN8B57v3S6GGjVt4tCxxzVEu/3gwss9lVzEPuyu//wFBed39l+ErMnoc2C7Om
FflmJLTs+e4hyPwQ0sfY5HRfAJmxo77hO2JeNE4Yih/UvQpQ2OAH9QvJf0YNjrR7+d+/+vorqbXb
tiOkW6g+AXbACRVQYMlWW60TyyjwaogVxBInWCXyD044pgfkRJuL7XN+dvxEFwPcngEgkVkl6DV2
wqUse90RQAi3iCrJCPfs7k7xmwEgM5UfjdcX3tVQiRs5kYkVUVARQidhAOtKIjmWcwZFV1jznmbn
u6QwfBsaMciAkmoaLJ1A571L+R9nDFSQ8pjhdighBGTqXPZtcbklGN5ll6QL+LdDI6XjI8rWcUAP
EVjKi526wotPj9Cq9+UjDnSpzAri0syHs+Al0X0yrNJq930+saTv1h0LZCtRW3R+Ljmjuzl0NMYs
SBPg6nR2Qlp7crROpPLZXHX4OqI2ymilnJccXAJxqfkknlaz+VkvOISM1jCVdNK3k6WPEP6uOqVX
KfgIyK3OWqxhzbDSuKg595cR8bY0AXfqruSwpclN5wsHDbl+tWsyvDmMFts88ECyzx/ySLRKcf7N
avU4VLddXCKbvw4SvjTT6Y47HSwSDVl/Nx5YHD9Sm8DqQxT1ivDhsLME8LNgbdUbbDSUnA+UJu29
5VS+He0/vnLCy6ZH/cS6Nwv4ui2PfXMDcGG5DPHotF9LBnyExAxyENppdlRKNj2SlRFtRpWSCyX9
BuI5886G1UMkOGMaePj/PtCeL890233yI7rRGIoXRcOZSmWGaXlorjVxon5Y72i3bM1bNPqOw/gT
bfl3D837iqQBrcx6iRvW7pwY2a5lc6ipadPcXvPmsX3cE4aa71JB87Q9qyrHkFSr++WWRAVFJqqD
mTCZYEl7uBU1mUTtEc59Xhhpb90WQtKS9eapJPtaif6Brd3zDoWGYFFNErh8TTw2DZHPXx+C9wdI
aocIRj8p0B5PK4K1SMBjBkRnpJ0HK+SBM6ChQ47zvyVpEED0cp8YOyz3p/9C+5zT7ebazuriYl3n
DSvsMa7qgzCB5ESMV2dHP7cIUD51QX2YzZvg1TF0iO6+pvqaiXFKdQj1kYgPcHA4TIHID0uWwzMb
okPlerYjGGRp6zbXXJEH5yX8bJqXF2ndwXDJO+QWNYNeN2zk+5OhW1sRDoABIy8yytR72p4PTClO
gg0e2BWA+iJO/HViBjld4z6cE6dEYcdDaM7E/CxPoc52JChBDZ7DiZfHTBeizfwrqtF7iAGlJFEi
2293J4y6ExqNTfhgiVHwSNsb0qsVRC1Eb5GLj0wEyucX7AS+y6IlFKsU19Er4Fv9dpM+38yuozVl
blfjmJhxucZs+gRiR+czPqGCX5axPy+jS3fkYFcXO+MwrGdzctToOhhvuRPPNSZ4szxWs2Ou8JaR
v4Gxj829tIT1UsFb1xxVuSvZG99pS7kLNFaRZ5BvExjtWICWMS7ovzRHwpYCXvLajkhuD9ZHi6E9
FnWr8XZObNjzX6zRugeQa9czTi8vVDFRuWOvoXkk/0ULF03S9vmdNc5AvLNlAF+bP7rJlGR3o7wS
wLqr1xJaUyXUEv2bkXa7S4xhgIcb+vf4TixjXGzlHIVZtuOK9Zmv5O8l9r5AAguViCHHgMTUjvSJ
TXeBJdeg8uEplis8oJqsnQW9PSc4iTivvYmjryGj0WJ0GbTScQAJAQIM58U9nb5wSAJvka8xCOBV
XfGy+/sahj1eNVEuC/rcUtHezHvjfk1YNI5n5WsiGxWZIDlGSeTuBt962w2i82C1Gik/Qg0gkTZT
3AHAmicZgtr1QFNwcS6ZmFyhtPOsOgN5MlMUxgy+wKUSBy+P9WRwnlEanWxB94G3W/rT/Gim8dlf
J9ggA346OdrLvgKzFtDQTcWoraJfHlKgBcXCOVEccSVxm7Zh+2gMbQXmLFu2yt3liKhTeIInWDad
X2nxteXC662oRHk4OqQRtDmx2dL5ehx8jSaY383fr8NBntvI7UKu9Os5Kx015La4Hh+rRX1vlGdk
EmazrJL87cpZwy1OWCdt8exfsDaS3uahjTJZUucHiYpQHijrNVVCFAX9+mvweXPtidqMRkrJOfxI
fzN1/fONNtN8nwXkItuqgeOY0jHAcF8xYm7b6gXKICWBnp+iSPE3ub24FyVXbgoUYCFTpT7tY7Bd
AftYLa8kSFDEzI7bNVbqHFz4fliCG004KUzkV4SWuF8KlLnHC+2QVVpkvUit9JhljrArzTdZvK4O
SQX97IFESi39bJXa+CNiC88QK9o79+7WGjnuAyLo3cQRQlqsG1IUICIayRP6RrvsZPwoSh5p3Sc+
vLOFaK664QPVuvI6OhCy6rYDDwA6mn/JZAnXNATZPOFQ+4rZ9cQVTbBfKpOTKoImoHAX8l4v/i6f
Jo5yKK/iXURMTeUKysnNT9JJ0xfz1Mi/xKVMcG/5ls15FZ00pbFw2vMrxPuxH1uwM1+U1XryxwnQ
FxNKDncOZmEQgaSjodeDyPs+3t1dgbOav/QzgFWZhO5lxT6cnjV0Nrq/JmX5U5r0gexd46vbtJ2M
I0EPZwrOSLd9+4dVf5hU8Xihv1SDmB2sp1MsMLzAB4QB3vZD+dqbDefHgZCM5ScVwUsr3Io3QMGQ
Geg9qHMwFrJ7c2jbOZQS0i4Gmx49f8iLQMFO4CqNXT4phuet99LGTTfQd6xk4/U1aIt1LzuZA+hW
yL7/HrYl7bm8bw+BVygP8PgTsKuPdAYFMKUJvsiySY/Uv6iSe5lakV/7M2gJ7DKfV6hW4kVrL6mC
O6KQlRJZwHfQHWdo3vRC5m8boO3QpF6MJyTmKOEg4JuN9yVvi7oJxIb2ClL6AqlhyogxV5FtPPUc
rnEos8VQwW1DOu0i92Yn7zmzZftd2iNgTtQ8DCwsC0nhRWilc+l6aPnWeB9u4VM6+omPFVY1RTxD
+mwj2az7pgpvrdnR/dDXVL3niHmpFTumMPJnxHEJsQtUecV6gvPNeLeup8KArXPMfoQ1A5ou0REL
LhuT4uYeJ9uc4WYqMs6DeHKU2Inr0I1orLXS0dYVlqdAwWgkffUKfnATV1Je6irrUUziGO8x4Dwu
o7/TUR8luF7iSxRN4tO72UqaPpmEJrCcCbNSHAzgHRDZnBLnBC9zuglUf3oFLeDYGaxJl4rcaVH8
kISOJM1eKWY9on/wTpFfTRoqJl+X534yV7j3l+BfPwPQn7JACP6GY1N7TrsLSWjbFR/SLimpjhG8
rqy1+Nu5UIAh/H0roR7/c6ruuBCnciqNK0qQCbi42TrILaX3vYZsYx1A1ioanFCPZHu2pgQoYwwQ
0oZwYOX7pf7ZehJ2EA88TXrmwhBB1Ez5zG6rLn062XyfF9FjcIFDhOiSRuiluzhmJBIstAd2luxl
QRii8BrydVBAQ82AplshBtlQQUxpEcxpbw/+1CSIVihZpVoTCHyefr5s1uo6bzoV2a3BrEvEsmK1
8ByL+JKWYxSiLfkpE261yfx1RYDY11RliHNAt9+afwh6qL49lER5Y8LzFKkiwGIOemySIhKge5Fo
mQX25+4pIuO39tEtGmOYuyBFnKnbWJ1x3jCQffuYWvItvQ+1jVE+UfZYmo1igzlUPuDIOtVrcWLm
FHebYmmDOKJe5Ui00XMwDUc/rVWuMIA+DizHRg+5WLrUf4XIgwMpNtK8ECKQ5OfutnPh4Bjv4Euc
wgWvcXshfNGBOdWuzzrdpUc1k6Y2q6NRnKXUUHWsK88rDSG2jZkt2B/TVwSNkv4cV4UjVJuEIBRd
OciXRifVcRBgvONlHi4LcFMquNIVu9o0UHqWG4srjMVr0jjcHRatRrFv/nt4R0YbS2uwu0OebVYm
Iz8M+cJrYIV8zz1dOBpjzV/CyV0Mvah91WBAWskQzDi7bCS1hyLR5llnPTKTOsQDul0jaiRpH8gV
l5djYfzKDwmnFaH0zwPTfje/SCKvmPJ5bM5+Ehoq+17IpKgEfhPVedE9HeMukTY5LkHbcAsM7jKL
RM032+xO6bs0kUx8qtNZ6uRcKCEd+tdwlSB8CuK+HZ1MyFdofTg4SiA3vWH684ei1GenGmC6WjfB
Dh0olGdoK29k76t3fVisrqu6x9+E6fbbH6+fZ+sD391KLeMfLLajmHb8ddJ4dy37/NF4C9AjsACZ
B7YJHhNp12dpweiqI05OD+ubkc8bd8iybxZITaCednaXuuN6ejQz5p2LBj8xB8hbIPrroXzI6buT
tzRFncnUz1if6JQuiRw0dZpt2e+aEgiUGbe1w8vlP25U0/hZMti84pQCWnQ/MONhr8o766lKjzLv
QH/dC6C37+dzuIlxP4dNgXD2hGiwCU4x8NFRt3wnwwX7wRB8Qeqp+Kj5qL8TH7OExVfVb/u5kPhA
Daf5DraRP1OBA8oECiv2hh1e1zqJFAbdTydb506Dn+ThF8mSWLuBsIGgyKTVmDAA2wQ+F5rNkg/r
l3Y0neGYogKSUtwC9Os80y+nnr1s1rV41Lm88RfHPnVs7Xeaj/gWEz68a9MWPo3dQ/sddfGNmCiD
zPyWhdujauc6kQtBF/Oqlw2Ui9j5PALrQVgQMrkL+56zrcN1i2lHSV3pvYg7/QPUxqVss3mjiUrQ
DX6889xLFy+9mfR1XhF+4AphQDSkKbdt5eog4TA4UOrJB+ECMefsBJRdiUIT8Oqg0cVdSfo1ON3o
oXQ5m4gQznUky34qte2EHk/mJFCRkSFQFPs19+inVXs0Qbr6P00UjNxKq3cnaY7T3BDpxzJ7MkA8
PJE/Bmq4gX1SsDO1+VdhuRV6jh9MfCdOuV94cx6zbhOYVjPVaA+WveRj5NPUsBvwMv8bim2Okp+/
mBXBZu3D41bDtU7fAQ0CX7gQPVcwh/iYTfZ/ig+gYwObKr2FFggcCwghfNb5A1Pq2QzDIvml6C8g
xiNFcfR9Q19PJ5FN/fkvV6vXuIP2MxReXtRFLmF+/EGjAtA5KV5Jcm/Ydcb3+l1CTXEkdGCV+8OJ
HivEaGI1vdS4/rtaMCviDor7RMdjN0MmFp6c5euPTGRRcabtOT9uyOnhp7A9KsfNPj68Ef4Sqo7m
ZlzBnrZVkUO36FPROIPJAbrvxXtcKPw6JltbN2/KBe1ejkDMKZxeKJfyvQnEJY+EbYKpJ306LUu0
ODqBmgiWnqJ78Ffl6NuzsyUwMqsjiAId+D7DWPc4sV33+faGFuq47XTOOXfzS+y8uLMqbbRl9Jl9
q0RwLdbi+V+XLbJj39FmiP1X1FnmsZwUfydsZ1zJNEmqCWEpNHG8PACsRsCP2KrdQ9s1ecjKgL+f
YCvRoYvOFcaBvY/emf8CnjXR/VDDQ8rj2b077udJBuIH+A0mMz2I+9KtBFMVM80VA9MALG/3atdy
kSpFROi4L7X9PwgrqgJSZAhE9v5h+jeSH5GFXN+uGLtITcA++AKKx+AxzVA/lmtrgoZBkVqCDWHN
xNQack/OhccKJ8GuorcTO3OHAm8I0dhEmZeTIs0C9wuVPXzwnK6xVTrItfNPMCWckbPr44FyTl6u
yBrRh7PQmv3aUmf/9fhgjkXx5leEaRReLABCQP0e0ZiFISK8EIpmSQ6d+7U495mjDXkAZDal8U9N
DWfB9ZA9rYSLgbj5wYiDGlgib+LjQljt3bt0RZn8BloCHUkaBY/lh4XCSKXiBBtnpgkZkFbX6zw2
rhe3E9ERBnHLrJgBcR/WALxjJPfHr7Lrt0x/0UjM1IOTm+s/M58PjhCbGsrcMlzdVGgBnG9R7Wn3
GA+v6QAb52FEoybpTdjzxofzBr2kwYha4lvtw+oq4k4kO2wzkP2gfBKZcatWty0uZSJQ/xnGiqtU
ygEGR2lGXjJn+ZqtlceT2SMQVQBXzxDfmcjWr5d/JOAv+mizJaVc2Rg9aRidSXtyveqEaXPg37Cm
0W1z5pwxhkmUC4Y79E2WkpPpBk1tROGT7YvVNV/wwT33pkDIl3vEsV09s8NQzJTX+xyHMq3NH3Rh
1YsUJB26qx2T852ThQg60qCGOFNT13g7iQWM8wKy7ejAY+W/94vUbLUIEEDuT9BaTi9J4TtODrQd
A7SJM8zBlu8EXdbS2+FWMWQv2GGenncQFCMTI4ebygaaU1/7V0JBvems0hr7L9Ic09boq9/pyLN2
NjNiTVXRW8O/+uc6lWq0UwvZHjcrR6r2MX+tKp6azKGM+6rut7RhUDtAoyhMcDIYsksRqDqHiFPv
R6zyBorhePT+iEhj4OHGHVMpT3vGj+z/6pP7B1xB2wifEf4KbZbVEXHVl5JgqTmAnTAwc70/LtC7
iCUyFh2ulV0GrrU6rF+S1GRgtlYA9YuW4Zz/gcCnX+SyUMEhRZt4s5rPgJy6qS61+JGZppHPliFN
5dNL7Dz66GPRMtpU8nuxb+34hHpQA4bHRk98+plT+8dPpxAJMHr1qlUR1/63OMsmsNDBMIZZAi22
cylWfiybV5Yld7UzZQpYNX/JQkFs7wkttdEkPDD5n/lfYFM5Bwo/J01hDSKKNnM7JeiDXSbqVu6Y
P4tImXuFyliMgsL9XhBfagA2UyH8bMVp+iXg+gIMtifreA4h7+N09Npg0jBWAeGk6vNoOXbd2OLu
W5MIc2QiZBsWcUvaSWXvuyE1va8y3WApAsTckts8mqXZ0nC3QK8adgdAbSNph26p98d8M4BeKdSY
+AKRnOe80MbYjLydosKK1RunFkkp0c7tzsSA3lxr9payRmleCNsYbIplrc8An/nlCSzHcCRvVzz+
ky7LehWH4Q1LN9If3e7pABZAS5z4nd9ukaWTmk/CuKyAt2Wx74ytaHpyB9u5z3insEk2ZwkHYKlp
/b+TXZd7Wpzozc4zLwXlDYdBHjDJUO7xMtQF2X3wIeRbja3TYwMPQWoL8BqCyxZ8j0UmnJozfTTw
zNHEcFTjor+Bnyw4FDqYZXvk03gem7j+6XU/nhz8i4QrruYGQN3pQcFHUJwvV+NNgw/HvzZi0ATq
6TShWEqbIMh4jzT3f8/osvR/74CqE4PVNZVXaj8OtD8V1eNhjfYSDtTaJttxMrPgAAKluEPRejgs
NN2tq65PrK7HWwRxg7vXjc+PInpT5I+ACGL075jeM2UNs5h6wtX4h8e6rwoTT9fyu4huHYHBk5Id
52wHG11qa9NkikdMax8XGl3aJZsJtrGEwS2PjVUmLXuWOPA3bF+ShoR/yUhRj9b8wCqvb7Yct/34
pXv7B+jIAHhrNerZMa/zpSOY/u0Nx8rmO7tW0fsawo8DX3DIaO5998jDyqhVcdEiDoIolQFBGfAo
SKGBhrHUFsa9NCExWhtWQelfmx0ioo8BQzAmsUoh3aw9EeYLXzutL0Mg22W+kL36zv21+7du6DkE
hEAuIdptJKlk/RBOqNsNjcpvSdo5pYAJJ1MVXQqiZsnzTOYcPWQL4pHgcS7gnOEW8d/qsvemYZ62
DQwlctBulFzYi/GI49uf51VXNSv2FDvfu4LqsOtq3Uhmhi5d5P1H5v/sVQxUoqXj4Tb6CWsQdJdw
mM03fo7TZraUjhSOGrIu92lih2gU0aTUdFA1yxKuL3E07fzbzXXdjUBVFUS/ZDveUAEkQPkm4GtU
8Gh/ksduKy7pyIkmq3oqLd7AmWC3nrRqjQ8bZ+IwDs+WncV24clppk3QnMLZvHHpVuQGzJVEYYT6
4QDypmTcT15YEUWlDo8QK1lm4UiDHHYNsqXYzscefiJKEGUR0W3+9WyKSLAVuGWwjOzqUbBxGqLt
I8wdjbkiYWxE1JWUr1wSi/PtxR7Dsvm+xiQ4BqY1177Irb+zjz/kTbtAp+vUc1gSv9Oe3dwecQQy
o5BP34hhlP7ofGVhCf+++NwYZi0wo4uSHUh2ln3qIFXd4DSpT6Lxs6XJYKPk7Ezr9fphzgswvA+p
iPr8RO+3exFqaUdfOBIl+oBGBpZZsqlbb5jHZi2vDrKlMJ5nvIE8TEK/3DTD/p1wv3gvNSmQ343k
cDDXI+OreiXKLiUBsZJV/J9Of7PgogmLjJlJ/EnNS21LYuq/8entp1PghaEOLSRbiYEmzFvk9CQc
TIiv50U0AInRmmiMlxsFR1RQqZJRwE+CSY4yKS8T8nx51bKIirvSSLbU8Z5hyaaE5qiHkCaLTsja
C82WOkiOs8MwjjDE6Zepg2FHaOFUZVBCvRFCw4+tU/8EdgEfCUyiEEFxXF+coilylBOt/imGn4De
Qx/F1/wo1hBmxBKnBV9rRx8BALoUgE1pFcbA5gfUKV+LxEMYa6RpCuZbUAFrMUxXcVzYWN4E7ZRg
L7NPrq5RsF5JzJU2XJxEMlD0tRt19f8C+6BkNKp38JFc7MqLGg/LrR5qMOjWhCsRznEX5W/78wrM
cCw7hALxObtCyl/0brH9qqIiI143tj0X3unYT2lqt00w7vSxF7jkGOxKEdepZkix9Qj/L2JUE9Yi
xXW6L3opyoPN5RwKB2MEg4NgfmTacmorLvoGsM7+5YE1mUSir3v5JJGY3zhz1+s3Jpqxb1UL62fz
ccXpTLkC0nUAXVTmZHxGPONjXd2jvSEF/I/nMxa/sT5WsciEeGd2YmVV1QO9uPK/Qc4gSVetmgYG
R09aTX19EKwXf3m7bNsCIrnagpdib2BtOoPH6bJPXZhx9wkRJSu9IpGiPC+dYf2X1NQVK2rsWw21
9F92cEYYtd0D9JROMMOp8a4O+bqr1scUx78mCNYtyR5lZh30bJinoWhxGLB2eWzq9RcjbOvuAMD/
XRTmyrzUmlK1dCbBkAMdC0UPflkcSvFjliWgWPJTAaOP0n1f+XbQ0gYXmb09HB6HxCsrmn8E3wIU
wj2jmFuTfVzizcz+Y/Y1dJuuVfaX9ixs5t0R9BqIhyLtxkvlbBJYK1SBO4RfP6ZtVaMbyACMdok9
wP+9nzAsYWtknIBioWPqqLuFn66VFyFJF4gy1PypTJd3FBrn7FWVJa7G/DMSr2jvMlMv/ZEVYCEH
6/lMuNKH3W/vVqg60HcMYa716MYRx/B6nU5kASCSg92BsJwbLTUkueUN7hWAB43FV/yxaR3I6aX8
5JWAQcIrdR/yJgFWo0/Ghtl6tiz/ZhmX6fyprZMF0XDlMEc0PcMH3HVabUxNETVGAVG7Mxzu7FWX
EmiGuFie5jj7A/f7PLk8nOkD6DbE1KMqM290Ose8t3rmuaNDSLnmkZ/W2atE8yOj7EYRpZVMzb0g
+WbJ5/ixNcbBMzKMQSSwVU6b5MmsFb3ZpRTWfnaUA4OR/UPfMmavP83D7862Uiu120QmYUNYQTvm
BOGSe8FS1fKNJiW/xTUwvtQMjD5LTtirCvdXW4UR8Ekn4OAAJ9KoZse2ugP+3mpSOGJ+DXm689gJ
hVcz0VTko3reR07FsbxGIPxCvl8j0IN0an8ks9NZTqJRKhsV6mGMAgv5yzY0OCq2E+OsyKwX6uKR
yRKkj2y5FkUIVwOvzeX/7YzvNuYrT3Z6V+Gasd50CUe9/Ob2pyvGf4Q3LMC15jcImGkbTQJolaPo
SXCQoDKMC9kEJHENNgHdWDOdsC0ozRDrN7YVDzK0Scj75n+J0GpxOmpFBjWIA91NEOD5wFXtV73o
om7wR3cn0h+oNvwj32WACId3aT6FJvuaShGyz9DQVkLnlbNtVaDJqYL/H1XmiqoDaouDJLkZdhlu
1MaEIPIoADkz3XGJ+pR0kAiGag32xMtS77PLqcyPKQNZReB6MxHVr0Qw80JDhWAVl55WOZVJ19uO
Llz+E50w+k8ZQxa4cTfI93IUZp9BxqUQhcrpHNZ0bFqcO+duYERjamUAC3tqGQ+uwJirhoWgi6ai
1DkOldJOyzqwzLJMZ4LTbiN5tfy5QglBxTyzmARBfnZIlsINq8LJekGlQprw5MlNUBuiiLjeLcDi
yPWbR5czKkeeBqhCgyPH9sqX7YuJTXLZ9V177QGTaqdyn9GzPgBXd6KgloIz4/iPLbI8BND4fbFk
iyYlqUezhvChoppLOvk2KCDkQm9UiTcy0l4z2DGS9yaghsShXCYDIQ7G4n8CVwT7v2LgsdCLaX5X
MrWcfV++2iz5IOjO38G0aWP7vYanoSaMRyaT7dCMMD72NCbITmCqR1DSiwiJPTAU0HsVV7m6OazU
60zqsciawZRFjESOwMWr6rMhDM/ZTQyxaRNzBcobn15vcDHyF7ZabfcziRFgQb/a+9MMP5ab6qDm
+29QnG+Gzb59X9IszpruSeU2h0v6smX2xpq25SfDOvWyFTSIk4l6GkIeDw32A1gPFTZtY7mdhH40
4FZExbebi4rO7oo3koox5WgjkH4sY16eWSCGyjvIZRp0gI12XKX7owapzUz6WEveQofpOdoGUBPD
lwo1snUhWsLbXd3lkpulumaw+u4fPDaYH376mjpVQJlQCx68QjWyYM6K7AfemHseEWtWyNE/fL73
f32KV7n0hakLh/+aMAb1QpNV8koQ0Ovs0M/PkRs6bUITAcTuEApwBJIbUtd4LmmNuBEx5Slqu2YK
+jlcqwsREy79iJnKirJXaDn8p4IWQkrN5krQxDlli/5nmrMMA526REzfAWj/rjYUNz7Xyz72BN7q
ZkITFSbhplAi62qsMUVuOD1gxOCw37XHRXa30NCUu4EB6fFzowRPRTmnbV+eXcPmR84lI+bzlQls
QNXmjYDDaZ3LmLv6bwoi60fea0lLN8WvA46y6d5/pPWTDdhrt3VnhZyNdls5oKi0eC6cNrK1SGal
Z/KDyRqaghcvhzMG3+z3Abh3aY2txEb3q/lM86J9zwJ50BTLnOACKAQ074fQfubEU4qufhSpYLkr
fFXLiuF0JOec9RKdMkdnpbjko9vdY3iNRY69AK2WXjHNA9ZkW83IfjVoRW8uHGZXqOmWMQ+RixQS
iinNhP1IVS2Zxz1G3wYQBG5/AgRp94uEryviooX04/W5YipACRqORbmqoUmCvecuejCG2Kf3CmMz
bQ9P2CaoasZUiEvUyrZx9j3u/5dQQKcC7YR/NR02c17R5PGehZnUmvgxb9YnkF7yh6L54rZshCHy
IpD1rtyXp0io0tvRTb4HIDObghNkW8CkXaCLkcat6BGMaYQx3vvy0TYBRS9b70dgsQY2P0OYcOaJ
iqY7B9w6XsqSMXyEcfDm7azUjoiSQAROqKeAphW2NpRiMwSmrNyNlneLBCWAFHQ/Wb9nXgeKzesl
2YJgRHEbfdPK/le8vT5wVCQz16tC//zNUUE+7laQqf59MhUMb/s3kcmGO/U0JnFH9UbB5Ze/8DmF
Nrm073973ELKnigdhZWtj6AsCxl41K8uAWZrZ+ZJhNXk+YikvTgSpTQg69yhbHFTcUYpLZIHFArS
4b//ojFDvPpaLSiHc0qNi4YoXKDSuOt67pRA/vLJMSKIaDgXCvqFOHMF5jF1sYgq+oyZH1jKlvwN
NbF+UZnEDE6b7HnKNQc+JrXrr0QoC7XKNsBawqB3SPYKXJjUXZiBOnIXPlh6tpPAG61QmhGTheku
hfDAQsD24Z7+pbLl6BAtvkJVJJNcCTH1CdRJ9EvLIXgENmZenLFnqL8tm7QkPd5AhiHGcqOsT3ZM
xuV9dSi5p/fo72/deFg2ebIGqxLQQk15pj74RD/pfT1SSU9lYqc9RCgYRA6LqfaTUZAAaVDiJ5IO
/+8YobDFXQ8HDBdUSvh8foPEvfkwoSsb1Yfs6CPlcZ2JyR9sUOXndrpz72ULMjK47Tda3HLuy1R+
hlGRn0To/Y/TaE8oAy58e6FldKSTpcYuBr1d25KOFsERDKla/XZFD4BaNd5DlRHcEjfO0tMr6V5l
Ru55t0ErySU46icUvuP5pqCn7QMeRUdG8/paxjY8Ok0USLMtXhqNJSKuTNhHgOBIkkRsiQjNk4ly
hIlwb9kYPs1Ks53B/sR3Xi4m3+QbCjCFS2oJGT/otyNzA+vWPr6iJA6Z1z6HRHnjK4NG3luWB/9h
ofPzqibN+hFaLklMRThCo22j9P34XaCcGTuznwF2fxCdD+IaB96l1L8Q1KIzmoCOmAguDVaFIwGi
LEDPg1TH6alVVqJa5wOFUP2I6So/chMB62KuDXfsS7RsfWiPBnMIn95jJtF/P2pgj2fVEujYMovl
pQxxn6PT6m6QgShUo0Rk3lOCFDTxZ5dRsc2BGvimC7RGZf0qJ7SVQUpmTaptoMPErB9clUKxi23j
2mOxZBQJZn8bLwV7tIQv3+/oRGSB94yRUlcNB0wIBbOkkh5CgsALGj62XAryu07NcXrI6uyXMHxF
FW8dXvcl54RUp7eMZKnThFKUEjxktWQsp5yqj2AWY7YILdQ66MlzY9eT2CwP3j0Xglki73LklPnj
UfuT+odVqEW3JGpdiBctehRtRt0FF9vB4iJlwwCIydDWqGdD5He+H5AlDmhGr+UFyq1QZntInlHq
5oPXeoLeKUwT0/1e8gxU0Qn3ZXuxuq2nTQ66T1QmuDTO5HI8ouLhek9rtkZuZ47xEPogfI/L4y+E
jYurg4ZMNayvjSjokNCiLy5M/WGYCdn868tCTuyVXrALXMqb54xu4knfzPbrypV4GFuQrwSiYXin
lwnk48++UK0hBbdfghaKQ3OKqHt+n2lox4wAEehKOoESfRwAzwd+soR7YWbpPne416gbaycpF1l9
tXQaknuDOViSoBY/WAxbP9wB0ilXQ3ySruQi8hNcxxklIuBZOq4D3/z3SkFyZZx0uPw4pvltDOHb
wGYwFu75U+EJdsl+j9gBKmsxMuAW+otEaWZPlJWrFMRl+CslOdgGOlvG3JGnB8i23mcdctEdlAAn
ymqYXfqEGJl0yZjBubb5cxqS/7mvmitn3SeFIbDjEtEE5Nzlakh5eUCKA64ijJoKsRshVZfKMx3O
SRkYgK6bVvi9xKaw5dElBIt2StoFypRB0+TEFZEetCavEwadWUtUZ7jO7FhbBxxNIxTlRbphPb+C
6HC9KnS4x9NcapjfvRH3Ta3Nnb1fdQxrQN0LZooZkShgEW1gFHJnvqW7w3O2X/JwAkwiCs6AtFuE
y9nCS0HJJQcDZONs5SpD+0fFMOxYtQJ2idmLWdNzFLaGajSTyKpZKc7qzgk2S8xGj3qx2cE7Tl3J
0iG+6Na1QSXlDuzslv/jY7IVdt/XRO4o/U5M3PTc2l0WkmDr52ei0zLiEek/fhsEVOdD+wNyp0gF
o2dmEC6RkeBNLm81ODgOAIm85Og2vKKAwVTJEjvLCie7AR09tU8WJHPP3UyxC+y6Q6F1lqv6M2wQ
ODcZZ+mwBCqk8W3uIMEr6/AvKSsZzOm6wIpEiijs8hApg+NeihV7DeBN8AhOs8ewNCVzEc8t3sMB
7O4/lwi84ChslnLZPM74JhqXx+3RREI5aZJ0yNE7KQwfHPK5PXH5vvHXq+LAEn1NEHx35/P+msrK
WDO/orOtLGiX8GKQvrHjyq7IrtWqNz9a+llevpszOc1Eb8NQ4SP8Vkneq9uAoAlhboHwPyLYGkT9
OLe5tZhZuRAkFaRbhwYKVwMHX7lq6nV/VbaEVDYk5sV+R/how0CAn5HfbZ+Q9IsdB+k7oonOq5/r
Lp79pcHxDPXDd/4QxVEa34uV4HhTSdGGzNC500eoXeFQ7YHFjVdYEFKvuAULAUZtxy696MBgi0jO
wGy/Ut2028BihY/kVT7oiO1l7+Isp61EG3mGeMPBGaPh6vOe79VbN8ESiJbzlAufcCPvRnTWEocL
cpokCnnh2SfE9WcA8pX8g6ap+WXcukh3eml5r7itWBIeQo7CJCZFjmpRkS06BQLVsWyy5Ra/91Yf
JTSypR0rPhLrJKBhRI0EoPykBo7G4Pg8MACyOSPU81ZsxfDmc2YQqWd0A/FaHO93ihLQcmaZxnUh
0zScJ+AooHr02Ec1I4ny2qifF5NgS4z1rwIudyNPCC+PjilguXcGq8Mwro2gac1vyNCPw+8yaL4K
UQHw8BlxCFpcTaVweuwwaA99lW2LqVOyphxp6ZzA+H4DaRizexi5OMWg2vwT5UyRqZEr8BqLv8R2
mJ+Ed77aw3slMGoZdUscJ+UNwmz0pflcxZ52PHKOxJBQTCLowJAt9fL+629MHcULkF7zzlLqYl+a
7WXB8hZztXIPQHSrp5ykWDawnpWypDOZC2kiKgMPbBVbHU3uvsvxyakU5iQ8boRsJb0uS3g2nWnt
pn7RMrFW5xiu051EU1y0xtu1nsXf6wOlFYecrC7126cPx/efs24I3SlT+3MiXMC5FE3ltw1W5crN
xOH5zjC3XUra/4daeEejmattzYbnvQoT4el/e8JnEcBG4K8Tl1NQ5ivqfuOs8YaLuAjusUgEtosA
43UsTIN25enCXk76MA4tDgouT5bFxARiM7HGLU9RSb1JoVF4wgcivLRVK8PBPag3DlHU2ADhDjKn
nk7SuWgUhtpPZZY0bCmPZQ/uunc0cvtEAZCCG2nKIZ840PAm6FJo8zusK6JC2rWHSlKPumJ/Hi35
Rgi1JgUogA2Y7vGqDoCbF0ZmAgzE6NI3VNg1gjf3pWPhFXANwvJyEX+GbUvvC3MRVbKhJbLGKIaP
U41PUxdCNroX7HaFwtVHxbk1d0v4V6gabKgBTF+FozShvrvy31aoB1QeiydMoVq1G6wEvAQemvjJ
u2huzX3snjoAEJ0jYbDHFgR6VMBreifCvHlxgOe2795xcJd/nAFrC21SNVjVRanf1MvCiorTT4o/
enQv/MQ931iuSXaCk7HpKfZqDceHdjiCVh0/NDQI1kAQ/G+9ixzkJoYc9MON3PAWGf2tOEFH5wRM
rjMDwwobXO4sHe1RoFV1l0nrIAYt3ls88Mhpw2/GESo4lAjE9PGVwRBWkw/GeK/HcRgM30C6zKxO
JQpzVi6JMFCnmb28Ve/rFS/IuROdVL+TmuOwga9so+XxdxFjYLvuMoEOnmH6jxr6orqE04Ev2rtJ
1JsSEZzrMg64fTdcj+XWUEMEp2aV0TGT+v95AmlwWN3KdGZbJBJFbX341nshPWvQBGhCCma5/Eza
HRVchR5ZEAXtke7SgJNqUaqbkc85CqmjzBWUv9D4wEI7ivPgdkXpsEJml9YjSHWCJlQ99FvkC8B4
StS467aYWxFTZKj5+CLQOTpyYKmgrsiePSx8lfRtyZz3mf60wH0BKDa4uFXf8zGEfMocZyryt4jZ
zDm5udk8ogkMbulyFfXqGdBEuXBFl+XQHmPArX3AQuhGQfVXDTK92N1fVAYxsopYCwhP/9lMkaJW
GqBG8FTF62LDuxTOOjNC7rxLyTvmra1wZIs11OYBGXeFO5cAj5yRRBWVvgSrdLFYeyI1FxnMQUx/
9UMlFk9dvmKQa6ozae2aYIT3ooJ3jY7g4OEV1EgmVTSW7bOx3HZhsMvuFpILrS0ud0zIopQt34Kx
tXtVPFGnYfO56ERz/EynyNSAOyCWJtLZ99I7zjsBUnFdhfkViuDBmwNfoijsnJ3tOopJzSWbdxqc
Gnvdi6x0xuHnByvJK9tU45QtmW4CCN1RWoGXPYNG3mGpkAyPKR+f3U4AEc//tcCWhXF1xtzFoBXk
AFW6l7rsGh75TrNWeITsfvJzhhrcbstyh1Zr4U69+mWs7CcBV29IN86z1FpHVl3Eu3YQI8Qteb49
EDi4ySRUqhVSUJLmmTDQbgBe+h1riyojiTrKRs6fk489jYLdJVIgvrMaXJ0agHL9WGoec8LzLEa3
LGF4sxIDHLNGEDfvRDeJdeSBcEh7V7licl3VGqd/ckVNfnzrbEJDWwulWnnI1mN1r1uYiAqUYqtH
Eun3KDjUP3NtlZYl68HX5kPpFzZ1S42t9x9nXDygTDvHkgS1XWKqknd6RkNZUvHeR0WyG0rdNjCX
2TfqkRZk3CxeMqx+bMqU/dq3X6Wj1g/Pj4uPviOvDCz8NbxxJgOvUZ0zsmnS1OQZgjh7vSHA7KhV
CIqVeVo+EhDCBVroQWC0L5Ox+gV6qydLyp8uvd1O7gvepRcEWYSJynqldzwgZ9qQxAHuyCLk7oVV
gFbFjdlVQWgVH4hiwsUAhlSdkXWSSb3JEF60eLNc6Z9w/HqAJK0dPQJRT49Lmd0W9bXfTIU1CFS9
DKY/bRM8hDwSV9qk2I72eA9wDPA+KSORXhYuCPr1WK3hm6OYM5nV05bR82CzCLPmStzf1gIsO1lQ
+puvZfbrk2W1wKztbUEtp6/DcF3XDUWL5AnPMyP3/uXw64wZfA6AJIwTuMsIjZ7FoaivKMW/V0Xj
+pXtEYwXTxJs9TMCSXMPaQAuSXvjlcIZPnMv3dIbtO9TtJ/qkbSAIqZwvgQiCLRS3mJ/gQ9PakiK
/2Lm9GAMSFso4nI0w+nnjuwqWDgfhYRFPg6kkD8Kp038ceevCW9K4USf2hc+43K6p+xSJIER1skZ
08kRrYfxEFq5dopa4kFIR1eJ520/IHyHdTFQ/IldgnW+lVnsfb1EUj4u3l1/JaHNty9MYww29ElU
SFT3NFdpHFbmq3A0nSkI/VfG9HAz//hX9aYAZmWstg4gmi1fUwpCYjECHjomq6WOofmIVBfEodSc
8Iju5zKs0xNaKKZ2OS40NSkSOnt1bGNUl5ntPTFkx+nYn8Y72WwKNroQZCYC3WqQapyjogRLDalm
7ieaWv4StywNmV6zyiRzgF2WVrK7ypAE6OkmSkj5VxTfV+xeMQbWZERjN7cL5iPYnJx2haXXi1XN
YlbtVja14zGriUFREnIXzxnk0/SjUB4U82yBrjaOmtj+334YSYujDAHRk9QUS60sBWMS3GFUEYNf
4s8om3HTGGZuyMa2TyGQ1yd8UEAG9Xhs+a8jICrKmXwa8u30dp91m16WzFRZjCbCQM4xFQEkBXvQ
JqgHSF8/tUDHzpJURmh5Ijmq2Y0T9i5cEV6ZgkmMUYSOh75gJPLebK13aK0Z5lh5qLGk1eQWVgx0
OInk9X57qd+SfaLWUl1ehxwsT+H+AlksgIlBrE1V48NWzt/Pb4Q+K2+W1uUgfMlG46x+iykTqxo0
705rcowMXcgEIQkV+miCwS4TaurxHtRN3pc5U29hj0NVLRON0wVsKMVkS9N+BMRYhJV9crgwcyzh
6/pBpWNOolkJDcuwXYX3ipbea0rP7MU5gSfRGSURoudpFPZ4opyOIkfbsm7y6nmE2UWrSbStlTRE
Bw7Jp1y8ZjzhrK2GztgHiiGGP4ATKEokp5jrTnmhhV/6+y6GrulLDruGtlm4UpNzrwkL5QIIYEVp
FpCRsZzehNFaRx1BHOQoSmZDRe1meK18SZYoAo++d/nbHqYz60AvTrp5QCe9vLaFJ6psSOi6FjGV
iBr94DmwR2QAUvi4pI0UXykAeCRenoVW8+a6OVA8F1QIa5XLMCNLTgI/cDvhI2CmLjdMPeFPmzcn
Z0svzp/ZDuaohmfSShFUgISHuSsHvQtaBDnym9mNP9f/XM86gdC3TEz6gpAiKNgH34R/91Jem3om
jrHvCNsyJSZsEWSYjpJaYBGnhRIhAAtdCdPgJ0WFzdFbN042RnKWHx12gccodLKujqcYpJRSZfSR
unBP5iHMTbT8Qxr0GNCDHFQJ7JunJ1LHd+hZWfBBWFGwVWymqcVIUTlobFJ6mB181ukkW5bzgv4H
GIHs6QUyarTOdfxEWSPHI/hBzoYwX5frUdgPxsuqrn+Iy2XfY4QF8c/lofqGVMWcCafDcqV9z/t9
XpqXMiQmJO/0QaJqc2d5bWGKgwTWf8rmO4Tbd5jNWcLpGLXamy+1adZ8yup7pXvkZaBFotL3lTaL
cynXDFI0Y6IyMP50Voom1O0CYP+D9Dy9yL/NlnfFc3VE1y9SezyJunxIZNBRrS6TzOm13uPgWpip
0Oajej6j1k1FT4vS0lLH7us0qZdhX4/oFIp5qacvdMVC4CEwagHxXe0PZLp+aXXhBH7loroCyyTB
FSzXL1WHHGcK+LAdMMgAAzrLo7/AvEp0SnmiZak9Q3xxrNY6BNYgoc+rmVyH+ywC3Tuyp+uTMW+f
QL9/AvEd5CHNjvGRGLs7pBXecuFtIybywkyFAR+nmkKVPIrDNpsJ/cQcEv8ifPC4gQfWlpGRow9G
cHfm9vQ+Ct0EQ9wUjppTZC7v8rubO/H5PCzzqdblLLb8j9mZQNt9W7Rd9P8EQ1lKTQ5FNjCj8fMt
msIqOpdSMFiR1De2cpSU74FaF18rZxxCCwW3NDeO7mgPJmMK9t0KfaTAXjYCRwWZPJ/BzLqWENkX
XbILNRIr0O6GLSSOa30PFI5W/Ic5zALynR1m76+XHfr/Q4GKPlH87djU0jxvA3oK/4qdpAiB8vDv
tvfHAX93lyCHdV4HiI7Ubo1XEaPALPx4ZZn0UpO85O0ZofSqA9lQJEH15dVQiOFlshdUbSmC8g++
+bc4DSwNGETxDGuPU3YVC05Aa8eN07MjACaTlRvIDeBvCtu5mM9XVjgegDkNk4efXqz5T2isehN6
emhVWibI9pK1rICevXgJbQigzQmaFXQTlOzhapmAoBNAZh06Ii8sYHQceDb4yBxsMLJ4uC18Uv9x
ywsijOS7WRYUm80GgMxWo2+/Zft3We0i7LqQET94geWUIqs8fxx5tHWERTffddOV0JWRMQTUUgeu
CFnubHoJ8B82vpZDQkN6YlQqugj6jmHrlQksPLO653L72O5wc8YmVzkmnwmt1Ujq0d1t7efsQ9Ee
2i5tUivXnYreYhSInBO2/K0i6+dVZPB0eOBy4k9d1FMsarq++ApGgXOQr4OAYw7aaV1/RNTB5Twd
hvLN+Go8cbgJdCXhjEOOpqMClCaL5OhWnPuHy0xdYviQS1OnQdb8OwsvOZMnEJ/jtOXKirH8YoYJ
akl0n+FPqwtivuTS1yxK8jbhiT3NiMOhhLaptV8LU3NCVO2oiZIvswTrETO1C+go8fllXYN/5XPU
I+/3nTy1EqWrGt+ALEe4ztpQuwjc9N9T3iDtotwHNconHo/DBJQWXojnKj6gVo8U0IAgGxofBgZz
MU4VaiJB8/cyKonuQsAf5/jQ77GgEUoSQPoVw/NSb2hdwxJYytEvfChKyU099pojRFOQ5CW/c3fC
0DaH59FpGlceqy1qIaDXdYLVLzepzJNhniM30wGDZhOtuVP4ijcYZHYS/U7xli9LLWwjq63cQWZG
7FWdh8G4qIpik+J/ntsyMFwdRqLaK19W0B61XyG9CAyAVxozMhgfjsnJibI7fw4323wnyjg/CceZ
Y2TRwTaFpPUQWPox1ps+Wpds8j8B1TX/O2e8HHcOEMq2QaUOjalUTZQ8tY5Wd3LM5I+1ERPEm5qZ
HVjykssqpwoGqXlX/dAOFoV8wMQaT9gFOrLuYgDjk++iEwW1ENp1WfGtzbT7PM/A1+ve/NH+F7Nx
/PXEui0wJhqJcHnRj4fxCSTUEzfIbktL8I3LqHZvVRJX+saab48wDXc4ASXGU2Sv7pyGI4ZasxbB
ennoKdNyz5xTCF8hqk0a/4XVeXdVUV+uKEmOZIAGxfY+OFyYj4JI2Hve1OI7jmRbxGyFatkFMsf4
OMI1G1QmzuqwmWrEsLho8kHotZJyJT/AcjiPoafMVJcek9jHlP4SKIXhGnzRXGByeSfJolRplAqz
OJdq/JguPMR9xirwVCswUp3BUzSIt//BpOSt1jiCaIRY4nbHjOERJd8GeQZzasGBlW3/n3gXkwCp
8vmFwdLneJphxYqKridz39+3V8kiNSsLjQHV04oy00+iq5fI+fclLTaXXRTUgVcAu4aF2lWzpH/R
jNbVioRi8TGG9xgh0wDfmNLo8xwft0cnJ+DKxQCstp24WIfJ5Cv/VRxctB+GzqHBpSoWmpDAMQFn
GoSypz4U1vp3NmgmMzWiBshURldjgwCSSRqbBHXXNCbdjyg8WoBw+0s0OnfadFPXY3Y0CCspfMKm
MvsaLH07s0vKriMauVSujtkgh+v6GJ0aqJG1qk8mvn69yQIoIBUhCKL1bu4SWxX3lacN+VIzw3f8
ibdmPRup1OIPUTCgtqXzpIJ4Vgw6To1LLiY9GhSpV0H5LDj5ThawsXlPdhKiJLcim0hvSdyHDI/Y
lM6EHi4AdLmq3zgewrfQFWYWLRnq3yaimQwKZwQE5UOLLbjLLaXN8AFs8bwWM+WxvIoNuLdDm837
LAT8Jt6wp0yLV4zxfhshGCdEC5QSmiNjnAVzl9LJq2Q6QpXRdeFwApez2q63WeN4RvK2S8gqF+xE
jt8FtY9NuieLHieKuokrfDdjJJshCbwwcqQIgYCJZnXWW+YAtL9pnOvmxJqxiMpySuGwJACf0nds
Tb/Rph+xhRH1+IOaITPch2MbsHMQ7Se9xHQ93+8vdAcA/BcIJXaejUKxtFgw5KZq/FetLVwUKPG9
ozd9ghjOUgWSWwsX2OMD4eslQZ8+5QsODikmZOWvSIZO0teMg67qCfYo8pw2WhDidt9QXr6rRcWJ
5WdCZh85Soua9qg813XyNSHG5Q/vE4c0MWabc6eMzpQZ4WpZBvDBXKYt7dQQ0D7bZfLLjWZzQY/6
EU500GX8rHye1zEnOhZtWmGfNRsXKpITsYG9l7HemjkjyeG2ZJyqQ9b7uvieoeU4oVND//SseVZZ
Nvm06gvu9IuWJy3HifCXAV25jP+jHLWYkv35IuUORDdsdsSeDlN0ZlQs0nXY4A5PMiklzgAXsf5f
xtsxv5RhVBfg74x1996TKf18fdhlE2eaNI493I63JuQOQNZyD6nqWughpUTtTimusnZCutuE/zxu
xxd/fK02aeENOdsUS6VttFKKVXsHx3NTmUlxbkg4pq2UsxJ04+oTwQJ14Tk4ZL+U2asGENKh3tJC
KwSGm152Q8s4JoDdsiYJYgv8A2zDCxxWJLpE0xQaUNhsajF4GL5ww2PDM/+tdZYtyhyLwGcH3o/k
hP0OqhdrhJ3EV6BnWBJN5p7C73RC1/0FMNehxNxF31NUQ7PDDNBc5VWhtQ8z9BA/enmHGMybwVuU
Jv389+A9hz4CgMFWsAjEjEXA1XgP09IXwyIThhkvdRthV1GUEJcxTz2Tvfny1dPqWYUpy3yoJdLU
nIEGZ9tGVIgzIJ6tPrcbQMLIk/hIrigm6hvei3RsgZfgkQS/QJJGqMccMXt7J3lQlwYn/3xIVLxH
rwCqGWumhbrcdrhjUMxmkmHVK+3F2m4DujqEX3qw1J9XsqktPC2ogeAZsbHGqyMpZnLF6LLm3hbm
qKH/lKsWsX5nwSwnNSPfuJha+Q8HgVtxmTpofJjFgwVWxebTMsqhFO4QpJnCNHyMmC+v9xZhm+ET
iEZAJASgcqxeMewaG8vT24xmXIcKJBHqnrcRiKbCtJkMZi4wEyWyQ5NYacp9yweRtEBz07cO84UY
ZBoWk/kKbxIfbCU62gSrj74ZqfH5BXoSj5qN0B5j99SEQE5HBMFWGBDGy6reoL1jGh97wdI9rKYR
yw+FdP0yBGD0Cq7JOGEtPNkqyZn1/KLJy+qBxx1K4GwhSCoGlmqdJnD45OwDIh63ewGTzfQ4DKrk
ecuCS/Vt0G9rQD1xVAI7VaBwo5RmbtAX4zdmI3k2O2oihF0WqelJHqtppOAQ18CjsMC2ldfSCIp4
JElBmtugrWnLwcaUfqQaBOfbn5ichdhQbtKIuRuWCBC0RQmuoUUpqudTNr9HIB4BdJf5iRXQjDAi
KbdgmmFe0868sL8Apn/qxmx3bxrbDL+7m3bp04pEOQ8cA0wEqEAeyRFRFu6dETE7VHLHQt/4wOWz
Z2wuXhnG/bBU85JK/7ydtB49c0Q2IEVv6ZXdM31r1IoaQvYTSA1GWONHS0wBv6cBqCyCQNMfOO4O
QqjhWGZUrroWeKvM/zEK2jvP/TBupR8rDgixX/vargrsA+vRn5H93+DEoGpg+SprlGlysfr7/tuR
d3ggqc5PS8MJm5ccEpH6Aka/yyCqqObhkgv3gBzxAQRXfxKaBHNal31TylWUNyL+tpt4CqzQv3ec
cK5FM5sRjajR1ddTme3ixl2ks+sZKJ0MMk438B3wBpTMb5RpXAZoC20OuvgzgjU1xJOEvycfPgmh
nFpr86I8yaXIWY8jt+VOTO2/uAIOeNITjwb/xXTdmNuC2gH172KaXbBhDsMlqeBJ/ZKo4NWhWYVr
kJ8E9lb6OkLQ0AV2+3MKQOGeN7iqAWiK8QGi8kBpx3oVTRGZc8p1T/0IaQvRgj8caBpJx8prhvh0
PZzuGC47ke+3PgePyocI0lQnv3BmIHriR15hITxzNPq+0Yf8DALM61roMhccXbUW7KpCUhVEsEA8
uI7Sqn8si+uPOJn7ffDaJYT7x10O5Lpu0wi56PR6kF3vXhjkSY1nI6ao+qCfFBj0VnfKNWxuMCPI
PjRwjETEKsQRiY4wsANkhDYz7dnCBBroVtvBI3NmAyxTuyUZ3pmZa30PIYlh8EnUMiFKk/wUv+U0
pa54JuILCDUg4Kw+qB4SVhxkmByGfNRvHWLQacTHVtPwcbmy2vXNeQ/+aejtlGYM1W2VT8abvls0
3FBK82HgzQBzwa1dBhIGTYkkCvNfbnzfzRt18G/Mazs/jPEWXX+3YLRbt6LxgpC9WopQfxx24q83
EhSAtItdz21IRk51/4J9emumxmV3lqJvO7zUwdh8vHYZChuNMNgRyufEWNsnQw9C9OwqUuz4ZwVZ
1fZTVUB+jSE3TJbBE6M5hlGvg+rNpjmRHm6tUJPX0lzKvSK/3uzL1nzwLhs399YiJ4cTiAD0lxxM
bt3WnmuxahYgGyZAmK33+p8pcpaDtTuWAXOd1P4c0+u7TERATA+IgzeYHZSJEgbS85iP5lrWMqWN
2PueSXDD5KmOeK4uly7Yt09Ik5//i5X6wBhUrpG2GEg3YLHiUEVSLmIUme3xLIiSdS7V1LGw8g3o
h/ez8m6LcD7d5ZUA1VzYTfTzoJ1LUIjcsdkpi5kE8KHrMR2uaDWkVLEvMO2LdnmJX4ccM3L6CSRc
+pFdp3NIDz+Fi2MNk8MUItHl4sjBNShxGVEXVjcYl9znx8npHjIxK4IgPgEp1r9pT5tH427Fm/UC
veobW/LSTfDtPfTYH55j7LSVyLNf6ZN6jloWPXgbxqWGeKVqolGiVNsPKOjZSoJVSNJbxa6lRCof
c5XcwUCKT3G3nSxiMPmT6C0Qj0Qggct/iVGlH2E1EUHhUV3y9syOnWUKvC0BeEJoJeNUK0NSLmKv
T9L/8HM+godtroWfxU9LvlNz+i9x2FjNwYaI+PuqMOmxgKRmFiDApZJWOPlRm/zwyNNXkYWSqhqs
G3YgM0OCId40K2usQaCK+fpMbadteDK4xYj7/B6Jl23g1fD8PMyCUqFWqxA6GfT3Fw8u1BSfc8ap
DcC2eJ1Fq345/wqSJkW27bJhgm5ismM1tTtv5RKkiN2MBPvvV2r7rdG0fKmUCHHj12Ku6L8alL4R
K20dwvZxXp+0O1qfXbVKpIaDyZPnK3+LPzWgvak1zVam/30J0XnczHknuqg69WoV90mS0Ogr79p1
5i/fkJ+WVDCRMRPw7I5g4f/z3Y+RSmyj3wC2JIPDaV7OVKtgT8Smrp0wB6+N3Qpb8oY0o6CZ5gG+
aClACa5v3vf89mHBsLoKzpxzUXAqVTxfQxxa3k7zTe5zl2E1OSpEg2NwgJbrVRQGdBAizUtPuzjC
f/DDLI2NWpYYqWB4OYqCPE+cVa6pVLZgAcH/p3p0WCjdxqRFHCvPK0Lx8nboAg84Y10ciB0M+7wX
h7QO6+SBcNmMyBIAYVJT2ChoWajFUS3eQsXOQLmYZktvI6//ZaP2rxRVtFShjKP4gbDd0qjMBzkZ
2tvDsFR5HfBEKAEhdAiz2n4JdGj2DwM7HW3ovxkWwwSsV8c/YQMems4aa0Ei+Ybo/xsdEmvBhIHy
Z4TnGU8WbmTuYD7A5xsCx/kChNGz6AMUw2i7YOrKi4vDg2dRaT0dTBHf9ZJGxlko2r+2yZr3Eh7f
MCp6cuQolT/dseaBlpey/Dy6SgKc5qqbTCoJYPwti+D+UQt550AKulZwNo++/xccHbDXDz7J/b79
H4q9IKUh9Vl0l5ixqvnqXRehdC3JZ0E0iJFqJVJTX34HR4ZVPRiChpkd0PWX8ZPEdTxwq3y7FiQL
3W7+VvUSQTDcH5UvCWUxzl/b1XM5cbMaA4d6j3neOM2viqdBEyqW8aWu6l1znKvUaS7gWQJ+/Ny7
IbohZUtyFlcunmowkUPB7kpe06FX0R+2Vqca8MrghFj5lUThFFfMYNYE7pzccEHUae8eFMAlfec0
oSb02AxfFcSKHOs5//q2bcKVY2JaVznOGr9OCpSV/MSyhTehz7wowTk3UCyMWg27fBRXZJnmbfDZ
B5y+DIRAVyBHg8T91Nci/ofJDFJ97OT+Hhl6GRHcP7F6ookVjdijwvUMxJpikjRL6xTn/LaF13UI
JGBNAUa0Wu2voPMud2uq853wWO/MzgLZmZyRbW/tLPtxw9TOptCV6VMSVDZDlzQJn0WJcnIRQXg0
N4Y67YDlPbswHtTS4FoOqKgauFnM/h5BOIj953+exbys1ntiLdmsDAzGXbwPfsZAoAfILaCdsu/S
5qRkl8c7xcW1wmwLq62KdCywqmMt3HGYbSOZV7xy7dTS9s+kXKzZbL6RMbd2obqGLub92uOoCYen
zRVsjVH/UNDEacP7Ymc8f3JBhporRVKLbLM9gqr+NK/xJLiQUqiRPZpjWiafCjt/+lj5qWCDziPH
BedLq14adrv8Xcc1JcT2zUbNLIhG9h8Lsl+0woO9GOCc9vkq75Lks/YSXLzZxF2SoJOAiIDAF0po
p7jglSR/GHK7RDpIlywA7mpQwCQMfA10mpdt1+Q8h5ayZNYnahRxcfF3/ULUqFyNoxIHa1juv07c
0nARSILRFsGcoySg7WJlYD/+gfZi4DEujL3dF4M8zv4uzZb6upxt+z/oyqfIsw3TYhQUPq6wX5hF
h43MUac15Gi49YA3LCUqX/kFavNqb91aL7hJvoKTcaDa+Zr3cJx9LVCXdgomXigbso3Hb3ehIHNg
45LUiHZAS2/S06Z69Wol4JEswZo6bp9Zho4b+U37cgzvxXwtwVXKZjdTmnqjNYb7ovJ3BEYc9f7b
gOdmaZXQZehFqPUxFsj7kjrWPbiTgXdsdRYluekivQ25fu1iy/GokH1lxpD54zXyfFsN2klMFrNh
aIGPKlA5+4q8tQrjIITqUwiV94hougtEERwfwXqwRSDVOoN/o3vW1PWYfDffqVaCZZOWSBnmnNnD
5h7lTSNwg5t/LTElzO3YEsqoJ12gzSqzR0KLhwRRLCBZZ2HU1lS/LzfudzrNuMd2J9bXwNLwPc/0
dytZlXuzS08TPlUGoqYHNBoRa5W5ctJGrDa4XW0blQ8Zn9RAGlDCZ8rbE7ooS0LNLGnzBZOwbM7p
Wsk2IDR9f5I5ht8AygF7+hs6wj93jdkjpsoN9sj8RThNfgvuyJm6CLtH2+HCOOl9bAK9qF6PQvou
fhUQo9/D6VXvxN/XXP6HXCMdsonz2wuB71Z0zUtK6RrxZQsv44UtcakfP1oGMhfC6fSBR9a6r2cA
5hCM/kXdbiC23ZVM4Z01ypA1t/wGsvTHpuhn6Owwn5N+lzed/UX7pkM3dujDsUUEG6XlAdVUKgH9
rZWXZl6B3MqbjkShswnyy35m/y+2235tZEY8M59paGAk8OwlLjK92cYemVOcOZuocFqez8yobX3e
nUxCCIzYlC56hKcROddB/vjjycxLJt1MS0mxmF1bUo7X7TZHXkQcf4vLBPzGiRuIlqghwulv3meP
cewvtSjnljBRVnWvfC12SK8uo+RzCIlSjrAhdZDUR1nIDEKgrWDNpeD3452NArRu28+OGkFxuye6
DSsUu5ooPiDdj7xGSc3ZPEzDYkg8XWjmMIR5E3j8dgrtWv4Rk31E0MTf0MQS2Nd9TFt2ET0pL0i7
ZgRosKLPlSAEvemUV1pFCBxpQdblPbdaSDQFkvxkt/nEMx0kfCMQUbZcZi8Gkw8Trj3wVcsEJp39
9OM0q+qs9BkVa7/UPQjDa0KLZEuj6BZEgT2xmky6Cx6CxMPuO1pqLrBOnJiYC9BIlKQYNHcnNg3P
Kt3yJ3hVS1q2dLF7eDtKJeLBthmiFu2s9ALUJRaUyXqt7slgy5L4d9M7NCClb7of39kvC9QTtXas
ZIgDu7mn2+qQu38aIXWWFdKdkOzIEz0KsMADEYOlUi2Rev86QsXq9Po1RGatn4Nc0qvwXIYYY4bq
XInJrGL5znUNNunFnyLahEJluOifq4OLCGx9bO+p+PD0k9OX0+MCkCYOivA6s9IwGfGRjtWv1HSj
1S1Euu1V73IYAhRBOFFlWNfxFGyxSXThYvN9tgV/u2vCSblH+5SJoDpVc4dtoTcVvzRL0v+yEldq
bR+w87oRtJW9O5q7V7f16oDxIVdPnPzYB5yxArZIf0wOKEMxOF7m4j7h74VSXnCD31+Xxp2mXYFQ
yvRnpdLTUT7txrJqqrba+YeDmziGgEGCGADnNRdfUut5B9Il1KRCmAkQ6yQbIP2d3qKv9BYwFpxR
343PxyMK8etHBctbaGDzOgPUmQ9KZM+8WOYMZZ58PmhfKRHU2v7dzAfnlssz5Or4AmAZ6Yz1bvjn
kvWr6oo21O+LwzHnzqcl0bwHPg+j1CunjEYjbn8fA8rhe8ZyO1sGIUmkn/5KHFRr2O1MBFWLmiVc
u/JlEtnQi0Pg514hbadyQoonR1qp+lJppkVdxMkTBV14ZfTNorD0uLPIGJQRsXL47Zi8M85HYQ6f
bthhZiVRgVnP2b7hBsy7Cw/VUc8LRgjEpE/0rTMZ3e/5p9+ckJg1ILoiCynw+RUv4lviSqk2FCBV
i4R8arL6tmtYcPXgcnic5JdLxwljuiT2Na4EGlNJYdhwPxtuNXJMNh/vZLZIR3F0w4v4pmy2EDGw
ExQy2BmBiBlSt8fl/nrmHBlxPZSaam6tDL4xBhcDv82UWLlv+qiCQPjfSPxkndJ01gQ/Vn21SH/Y
6c+OtFpb44itElBJ6Hki/zVD45LdgcEsSyS4TOizyxvDgK2h+FGSjFff6MxRgx5K1OJWilLUrYT9
TR2BG5ZUXgUjybAy8FhZ+oJvsZoPgsLDx5kvxTZug7pF2eaCCXPX8bopEA4ep/yIivl7mbJd5Yoj
lC5hy6hzsGDTGDGSmGTFTRQ0DkVKuVpqTo+pXjkuFJmRT0Ys+dTdmPubvrgXfI7dnj7NN06gT3ue
DcpVOry1C/3C9ECR3fco8cIx1Ljf7IpYwE/5m8py7L/2bM9C+JaVTScEkQL6Lpz2wvRSv+SdzIvQ
Mo5xaedgBcj3X+SeUGc5Gtvxj0VdbFCTvcqnxXa/X1fplF0N+rjma3azJtHmbv5l0zzV3B7a+sXt
mhkidu5On0vuT9hbITGtn6XRgnvuN3JuY0Ts96BlIHCpbcRSqktAhPDE/8456+yuCQTS3b2ZUF3e
9LRcxpAZ97mFPi14hcXuCIJ+jkg/r+0Pgkj3f9bPW9kLmqYvW8q08gNG94PZt5s6xH+R9bTGL3XP
dhtP0dJxz5iH6hp5Pu1mmYMDaD4dYaamhSZ4K0U//NtAyV5v4LDJdoeVDlj50ALlQnHqVjh3mUgq
/iK+sHstUaQIm/eaDrCMrwWv0g4m4rgMq+YtoH+PUeL7XbzKTgcK0zgNdxQNkI/Y3r686R+kGZyK
r7GL2N5VAgcI22BaFeYqsUzc+ojREAcKXCemeQ40PA1FCTUJoEwslTrFyZkCcWhdf2vzrMfk5DgO
lQzc2iVlsfA/hOPkNLlmw1t6BoH3cV4HCgljbkzYgQxdA2N5N06XmqXAeItRUHhKgdkYm0fZD0lz
xpEeb0AR9L2EtrreRhfLqp4tO1wpZWwflLUSWP81dCjPtzGbiBcgCjALQJyo5PoqixRWBKV4NnF5
RSOh//O+u6K9/pMzuDl9y4QFV8M9mpa4ors1tGh1u/9uu7Cpr5kVGWb2NH3prOJFg1hFYUArfY+w
DeXGaSCaSmRww0IdBkNjsQI1WpRS5glXx2+Fmidtsa2Rv+LOuOvZEyySxmZuiAqTIwoAw8F3X/S6
UvN7QQifkMtOF3jqYWBzvAjvEHTxUgJnsnOGQSiTCXKiHaNb5gRtIbfn19ekciTMGbAJlTuqJ2wU
eB/Tn85y0Gz/fk5OtyYWlt2HO1eZj4LWW8Lp6zPRlBm2N4jYGJfeeaFiuDLddUbpQqqTlqz0vj7r
AtgsDC/WBNw/Sxg4EdZjenm03Y3k/H9oyaerX0k7Qga3nuOuDnPuUPNg05qJy5i6or1S0sTzbAsp
0BsvlvoBMaeNvgrIKOard5T+8v8YgekeLBhK1k7oP4mG1F90LK2jDeZv2ny5ox7AWllTLF0eMY9i
TSf2VWij2qWRdufAN5Yv14Tpgr8Bz1/BSas1YGwYQCbF9H54UAMnN3otQxuBmhMdoRQH586xPvOc
zMEWGIr0Zo1do6C1YjII6NJYIi5sweQPyUawRXytIp3EIAS/Juq24WHheyKTcp7QmsG9kFF4uXCn
FMPYjryXhezFVY2CeVg2Vh7dmfjYdND9XZjY4AupJzAlIbJm/fgjfDbBxpC0p8ZGgva6cFKuoBuo
oYxzcpXzrT1JC2DA0I6l+/uSLUE2bS34MN0nQfZWGjZMXR7w+L6vM+C7A1Bb5b7Kci6jdAiJmf8S
1OsZ/jqNVns2/Q813Y7bw5UnBj7FvcyfXvMcqFvbnHSRKVw5HhKCNWROMBlp/sOmsVboRYs02JGa
6BALqHpc/qg9zVQfqfgzul+9tTSl+FsnuIZCoVOHcHygftguWOVYAwaAJq3lBDFS/sgrjwDHc9En
E5a8N8PGdqjctpcjve9oBW60N9VVQutUfw/tHS7vkgatMd6AT20bGR+CZvppH+N7wBQx8oJg/e0N
17WYzxxoFhyTBBG8pIfa73ilqzDgQvt/db7RZkZih/oWjQU8ufjEpIqMChpK73/UVmnhanaR7AxH
VvLVuz7g30SxQFP+Pc9G80xFl9K5oWuwaC2m5ArU+86zVI2N7JriSXooPjUl7f8jXoO5oR0MJn+X
mvcJm5KYL0MmNp4m/vn4rWQzmiA/3WLGZF+sfR7ahk0VFZfh1MIPTrtwvw5xkLKVvYW0Iv4MnDtG
LxglbYZYsL/RJWzqS4B9qaeyhmh6bZNOaexD6ZsgaSlkgOXTWZZHb4gQfu50olSRPYc5YkG5oZAQ
GPCEVyaRv58Ozchujk1xWY6THbXZeo8dL5LIpBJDgo+PDvmSczgtQON0Zor2MbVJJt71D+lY0TEB
7aV9sFtYlxEBU70/ABYXfioQraYA7SJcDSUEocpz5ZWiuxt9zPc8WzoeGjWM/RwJY2Xg600U7SeG
tnhXjLqCA+4yc+DQW8p1snid2py/krI4tuab2cIIiYzLDmJaJ1WzkrouVO+XuNVQMF4AP91rZMWg
yxdz+t+JzIdR9yE6EzhgSQahXcPdedR7glpWgLyWrjCl3nnqTWkYafRskA5cM/ga+VUjQSefbPpw
t6sErJaFKYN0ruwJRjS1CeXq9R79q1wiqUgULFVMU6J1/dG02KpHn7jyNFGkDlalil5Ozvehcq62
HmL0FFPZfO6IBmGk0NU9SlWd8M8YZCUBr3MBO63NFs0QmFIT92N6tMaoCZlGwQMCRlT+6BaoZLDw
aUq8t2STRqYRHCl6dng10B6Q4z5FcJ6SYPwyjDtE69xsWFXuYLdYnA5VcDwqHQCu6ag1NTh7p29v
RNBcewRz4AruM5HXJvzBcWOxJV+6pMHq83sMZ5fZqFEnjCbU+xvBNzuqrGNgDZ6XoU0wmLYpgosv
iGxPWEdZ4QL378DsFw0kTU5WRD1FpLC90N7SlIEOXX9t1Ngs2IFwoe6cOM/awvn0bP9hpPMdtiXa
d4Jt04gs++vmxS4Fqt7OY6hCGCbTs2JwDA9Awr1mV31qUTr5DhrLqssjWwnqmslbWB69GKHdecqU
LM44njUZvAYV0i26I8hvxu3Iwi0kk1zEXGbRkA1XtgUJ8zQ0xbKBgI5Gnzdthn7Z3OBovOzqG/M+
ZrWbZLzVZ3KpLmlUlGhlP2o+KwyDlwnvsfBG5LjhI62mbvf3l4NGsP1JYKdvQ2dM/Kc/gT2i+wiI
o2dCgm0/fIyvI89eX2ScioM291QEmKg6lJRKSRsp4ev+c3PvYAF6tG4W599rUTAi7He91Vf02Mnm
h8DVFQuaSshR/QwV07GSFNNS/VyuOD+Nb8NfhCkhVhF2d8rentuLKq0EmZtg3iyrqTogt2vhUkw5
J05buG/50/VVqZDHWpzEwYeUWif9GXHJKegw3mUmC5hI1bzVw2BvZxtoXvYfcRfVPU+1wIQKDUuV
OpmgbHbFEsPLlglsiZ2egfwQbs1ugrFu54QJpiWWI9DHJaBC0q3Rw3ZgXSgtsGpvKFvB5ViefZvN
CjUUMkKNB3VVOyISN4pZENXgn2v2T5SWd/3L8HB8SFn/5F1wsMf/gfaErLHXYIcKxGvUSDrfQzp4
mbLm7gmq5wH5B6uIMydXOyNHAkXh0iLy4vyRwIBJZgLMKcVcHJh44Sa3UG/jIFT9zNvU1fpstgiV
WnwpJZqdVkrzDkuPyCkszVNDDePDBZ04PurFk+Zo/+kfGLj0RBZz1kBj+uEigNKSEJY1nysv5L3b
bFPdInZYpThSN1c6XluxrcxZ5YV6nDyz4avMUJ4as9ne/rJswdO8MJFxsudZzTwH4FNHO1jg5Znt
xeMcWUrjVkEnU3AGBAt87FPRx6c7wjizc1yOnl1wSGgXXNM9vd8BKwqznjjtNpr0j0UBLRFV1ukj
J7NWT3aT7M/FCtyw3ZwkfPQUdi6h6HcW1zAhW1B//oLn2dkkNVdn29doqZnmUyyVDwmmWGdTq/4d
LsEjbGx0QB5jrB+ToRgrEKjWgjQDsWrt4Kk0NccJDyxustvf9imJGD6bFuMElFRVcBZ7zyAxaCLS
+fq0S4B4t8JCujGpNaCnTzRPiKdcgAt2d3SfF8KMblpL7BxuvLBeV62qakLKzUZKlotIocsKlUzG
nSfUuyzkDTRugbahPoOrxHjsrw9lzERYaxA+KdWotr30809J6htzmOnIF+eikGUhita7vnIA9FmQ
Bz3ZBBg0SY7VWbkBByoThxREvBQXXZWam5ZwFklcQTFDCRcQbwXeW6hBPwsx1Dvtx9E3DZTyJrd4
iFB2YwxuK3WbdEp+29gpPTswwia334n5F+zVZxg86zpaO8iAWiK3lgHBK08R8oY3L1V3qKMhSqp5
NtZD7CBuy2toj8UwMT3tP9JqaxpHqA6nVJL/Uuv/tR1209n/eWsWHiU/rR9CjRqLjWWrZH9Ij0le
Xrj6auvxILz8ct7DsELNuxM73W/7FT60zS74p/qz0ZE9B0eFQPsOUGZb9rmyS6vHkwZUpwvRE4um
9uv9Blv3g4BIxSCjdLzqsf+bE/zC/hizCc4EixnHpdS0xYRyCqCQZcH5/B07j2mvSUCTBRu9El/+
m3Loz4RvbgoIF1WissV/2ernea2mqxgIybSl6dPjyWmHCtQ7KYHofqz/oygp0fqV0rt5/DSInNGA
MLVQ5Ug02PsntkclC7+5SGtTXsjEb2BOhD9k6Cb+dMEKsPumnKG2Fyb4op9UdrSp7GLmodvcZKbS
ex8JSXpf6zC9BBGPVez6y8riFdM4J8l4rVNzPxpQ/moW04Aslh3wBTkRJ23ggO6FlWG3EuCFFc9f
pikYXHrWzMOvtlrR+u15VSE0BBkWOFC4BB1I9vBvrZLJ7FXz3A6mEFjBPizSo56aARYzG60nTY9n
qGB9zf/X0kobJ+4JJwBXjt1EcQdw7WO79//K3MQ3PYA0tmafMDgXUVJUQ/oSWKdIrCMGOOVTEniW
aPK5xXN3sh+iiwm8wC1KGyLhLOilBGJh+sQFcQ0UEHBM2dcXmDpLazKd4T9LuBw7rvYJHah5oozZ
QQ0HHScTnkBE2HbXoeFAjtIzYxReZ9f2bK0blXACabCLZQ0nRnVX8QCdF0F9AUh5jCXfooxZAnFP
vjAgqQdLvD+cgwMGei6qtYvwHXtr5koLL+qzz9Hz+l0SlT4sTgCVI4NrLLaXnIXNjzM+N7wz5lMW
WVKJGMapEOHZQnNSzII1yNaRYLCvy0zo5q6G4+xzbauqQ9mO2WvjZT/dhiRM8zP+GaeSvpIwUUwP
JJh6F0un51vnBaealUvAxKjyv5HVdSb1fIahriITP0cdClt5pA0H84d/l8Tx05/RUC2gyLoV7Ae8
KOwKzv9DR5X7uYwl70WXnWcXrZVuXKWGWiN73MLpA3dLCZruwgccB3xmbo44rYWuDfZWQPAO12Qm
ZPUmelLNe6ZvNybZNaQQNwrtHKfRzxuPW5ZhCA/ZVuTE1eJIVB2lji+QG7GvopGj4DJ+eAnX9I2u
6uaiq5a03xAa+E2esMHyQAIY00eD3C61qkaY5oBTVzKF+F4+7Iff/XzuKZFOJj/Z6Zz+XuT2GBJF
xE+YDrgNdqxqz3XhQKEs+jmMDuc9B8PLs1eVyb6IKyf+/rOwA7yMp1aCCflZAgZbXJRVWD0mox9u
MuvdY6AxKu+Ihk3BtDtutAgyE6wgsYIUcV4YdHMpst3iQ40Dpji/5o8b2La2LoA20J7Ru+hfnm08
AEuFT50kT3XvB842IeAOba6j9XRRGMGGoInuO+HltWYOWTo+7oyeX/eB9vAW42JYs4KvWB1ePY32
6eJED0Vblf+uWUY9T8DhSrKxYL9jAGNEw+/tvSG+2SMQ4lGFxmyrDOw6MjHeT6Z3lWW7T8bQL0TN
tvlQrHdcejPY0xJxcGXnnV+9rDxjXcKV2tDtsqhGi6gabu7ychybtL+pwDIb3eeyLJmLlvgfEcG/
czm+DHk0uYotsl5E5SNneU7Egm8l9sI9SpKTY6L9UIFirs6/E5UJOKSl2MCpAJMW8Fmx5PLGaGfA
FuAX/kbUzjR4+EARupRjngTlX0XlyqGAQro8fvqmvMunrv2D0S68VeLEeenkH7gAMoMH6Evl38O4
n+ssj5x9qgNBeBKb9H4CRwKJkVxmFgKzu4oNsfFaYfLdWMj7Yf0ME2QllMpn1Kc8SSuhp5SuSDHK
EkG7GXeVVu/Y2jkYk/+ZdVJmryNPozYIfMeUpoFgx1vt7MGa0OxnZd72c6I9iIRTYYhHjZMU3Pmk
FER+4cEfUBatUZspfW78x0Af0kEOHuf4tF8BJLDn8hgm1ehkx1tcBZau0oCBHHx66Gsgx1PHEOAO
WqTMWmla8vSppc9fyAa5/JE9kMLv/fCZL9BxoOtUePWro3eJioz83lesrakhNJy721CNUSxSVyK9
Z2tV6Qr7SoNx+MbDRJqLgZKScQ9biDw2xtHKRqnnc6JuctMPjxz66dn3/TLwzDVepJOBFeBJ/r88
4UWAObDaORjHHljh9AH/gWJe8cVBSMezWmlTXbSngsOwQha9LofIRP42NTvYK+3q5EXh9QdrUw2T
HT9TX9sDuUTKX+UK3dJQCKWm/HpvvW4dOOsd7sJM7m5QV2W6VyCWErQjnfOINJSM7blduL76iKDL
Gsm40gi7HAMt1G8D5lsV6cLY4sxcuqHUf3Xj4G42CQkIJrninERIr3YDNBKRobXAYegdYelyUSr3
Aqi9Yx+EKZgOdbEUbBVU77wxECfWw+Zyr2DqPZ0DJogXIBuSxFKiRy4lM9QmwTvt8Y3VHKKrJAuP
+ZzlcyXiz40nDj21o6OvPcejv7usv1tXCs09OJaE0g9kqZ+hWcG11zt551YaJ8xdHJmVtUnbJXTG
BgnGAhwi+LxdCCE7lC4imZcBQbbdAkS/sNcDXjEhL9XvGPefSNyhPlGdCmIpuD/jbH1f3U3She3v
Ml7x0bdc+sFyuss/K6x2BMaHjUpMKvQlmVjv9uDBLQplUUcWhqey6lAMztAH0WvCri1UrVnA1DuW
mEyo2HS7pN5Twz0FSOYzO5ZRSczeRkbTNF1EyjlnSA77BY3WwJrI6vk+pmjQGTjLZveOaOH9a3vk
F3sHt1Pu17m5/GdwEDE1y/YX/rKVxMpTodVBvxfAn2v3L3h3Jl3cFP5bdwPvui7DCQdi7JjfQLpe
HhlHwLsZjrFpTuYoawt7uj3fRhdxF6kSraMu+JTJ0dTwTzuu+ZNmJ9WPoTOjKTIdKgQSTzXVERAK
2dzfu0y98DHyApuK5azTDOw+zvV3k5/MjKZjfgBtuN/AOp3K8XTOC7qnI8w55zZpvFaHJjFz9HUv
YfajfaDFgY/qwm7SZcAFMXT2Xahpg4nLKXMsOO/sEXsy7hUQ272Wed+CdCdN888jGnki6f2sThZ0
6uYzTaEHYSpj7pUIrm/u1izrd9mzSGp7RmaybyTUeDYD5kufx9GRXZzmuukYoDzuVgLbjQLO9O3Q
9jBUBuTzeW21ZOjIuyfn/L70kWJWzMjpmGaSi6APBYRSG03zFrzXF6x6a6tYuoDODYi4QZOWeFJc
cdPFHla4YZg6vDuZ6hKOVUhrWOSww/A3ko8EMH3Sw5D3Gz0YG9a0gvvFBudXaEbxYrjO0M6T/UKy
wS6yiPPo3u2Rkh/3fPchqhegBa21TzWk0o2cqtI7MTNE/vjUSKCzjCU7G8Rv2R5tJkliZ33/31LQ
Yz5/ur7UUpWyboGKNsER/fOc5JtVQZxLPmx2sfg4N1JXHho6zztxe8BZG0Ct7uPO2dx6su0QN+F2
+MMoHEBoAfobi34KV3Ll8x7lUwUvxqqvM6mHAK0EJaUHxFbW0f9uqhVFk6jWBsNGgVfxoYafSn1H
+W0QDTeuuab0fuoGB2q1TpcBMCh0zsS+i2Z7hk6mlvnJlurpxomhjSW7+7NvTzmDuZv7i9AebwOi
BUDeUVSaD+W9gg5YtogA4pWG7Hh+PG/55G8S+QoaU0Qsi6+fbiVD1SuealWxPlWKG4h6YZguw3RM
lsL+CdnhwrMn7aAHLIB69bOWKbPd3P62lZ/1wQnJ27jrZMBc7Hp3fjH47kAKy+KdieXuvI2/HZXu
uEUoaK07knejSggykIKDvlyN5x3tqmKeRwqiQvHY32uzLDyCPRqPFh/7KuZtfocWJUyht8d2v6a9
f6CdyCM9aAW56PYYnySUqjIgjxszhuFsdmMdsDjW/dIiClEI6v3ZHGCejGNGuDLZqVlTX5kSaEip
U5OnBT/c0rJ8IprZJgPSK8isfW4O0RNf3e57seaeAhkrowwyHiQ1rSq8r3CGPyw7/WGi6qlYYYR2
FlXS+sFrzmcc/eVa9gzyBeA3hGiJAWxUOLJa5PFhIqPcF7DL7R80shDjJJRre+pgSYs96va4VQOF
lAEOMtvmugcpbXQQFePCgojfYcBBGKZ7XvTXAhs9LPaNh+LIv9PhDtzPti7buWc38/Q5BuP5x4Cq
+bCXYjRLY8599B6t4S7poY+D5dixU5KLFCUPDxihBe0G9r+4ufHSDDq79g9ZC5YIT8EPgrHLc5ys
I5a4z2lIzzXibvyq5NHY6dfeCksjYSDMsDpTFo+RR6vf1yeUUNnEYXpeEh7DVC5+6AIte2jqSYVu
SKiVXvBLm3TYisvxbe+TwPjBTVUua9m6685td3Nlbznq+jeORqKUqc6cAygqBw/v7d51Fxbk5Myb
I/Ra1tbYaH3E8EhnAg4E+7cZUxQGSj/REzvufWmznrvNvQe28n65T//vvojtUL02dlMyoadCApYP
JsjfrmxbOAfs0pHwNcsdMDdEfgMMBWn9h4jC/5gyPxwtSKR4HgWiW9I30JYlSDwkAINF7GdTJWrr
yDKPWqKH4p6lJ/7f+B6voaGWp3/lfniKo5uOX5ugIRWkYl/acPRzO3bQcYi3BRv3h2cFSdcz/f9f
RvW5blEV5qV/6fqMaVze5Ij6EYuIKJZ/1cxt8QrVImcWfa4LDJkXqGYiZXxfEjmtyVeK4XdwDcH6
EkbtqM4biZxx0pRGla30FjtZNs6Kh57ryy0+AUm4iQtxHYd2ZGCAptz8alb3FoEQqQAL7YDKEbOB
N0PIQgRWMAfknxdJVlOCVRu3DJy8I0uilFFn88PCdpc8tisNre/rG+/ftXFD1fukuYtoSvxyTKrt
h/Wb1hBBnJPQ1BtKJsfB+9s9giBKnFnLfIq9DqwemqGsCGE09XSaAR4UhZIAVkG38eM/9ZjYgnsY
3eDacdGHUrGsX/hfXwTKICtECun/+W0iNN17bqGX3bNlBjQ84X6m/+Y91ebl54D6sFfSouqCJQSg
0iCBpisLtZdThZSihdywhWkfKpeUgi0UDZSE7AsO0OlQ2Hv5N5Czh/C+3puyutl+w3B6X2exXkbf
mDqQFUR45Tyh5OGQKPNRnjKxcQh3KDBACFeX/PKx1rPomYXhzSVmZ8xvhhv98Iv9KaXIEr6e89SH
wPl5rw3X0FLUrdqbvERUa0OHapt33FutmfuD+JmzsbWivPBl+535whrhdUHKC10Yr12gJRQHhBFi
aQ1T8Jt8lAPlwy03arSQkrME3bgc9vzYrwVMOpF880z5oD5QrQcG7RADd30aGp+/kblfOVP77ZIW
zZGjYwmcURHJtFMoSRvNZ1K1Ir2G8OSTEanzDR9rCRKzwEO9hzdS2UZ3ZYuAH7Egbt1Eno+lwFxI
1PCAr0s4is55i3uiEGWYRxmlvmwndpua0qR/So+Or6Hv1lNxKu2Ci0yowJ1igMRyFjpnw9d4MU1R
gziMwuuhtLVD3zZPBHcwxj9dEGMlAAPCLRy3wpTKa4/oDSRkN0KLlltx0S4BJ4fts48a5Lr3PKlF
GDOGHT+NmXRRxYaDA+1vSSHH+S7VXwcdJvLI7I/+myY6eDVbTEhKbdKoyomzjt9tbuRlETWwZ67A
j2a4glJly3qiUCrSm5c0Q0oN9jxisVJkzk8PPeyHDbmULVRbWwYQDcm0Tr21zp/U4rDBYzzgNE4s
YmvYZIG3K2+dpM+dvfXxiIH4quFgDBUx0eipPSfNnhCLCcgzmwwbboJbOp47VgRkJe1U4BSArdmF
NfJCuicMwRqbsO6juAigVbuVknEOOuMst6h9oNk+MUkfjdP6Irrk7VvubwQJLnjr7AsvL7emXnMP
p8doeM+B6KZFpwZV3q/vdDhJS2wfALkbT/sipCGerV3jYpUzP3vXX/LYUVkABRu270ac9Nf8IGQG
XDXpXbxY9sGlGGvKsakMgupyFdKd7xGmO5+T8YtXEu3nOJryPqdIug8v1o56wRrzMrusBh0EWya2
jm4uf0NAobK1r+Ui2HzM3JrMLDZGVHmpn9T3hfk3fTqodwYXsjGPXwYW1vIBc1Nx94BfcIbuMNbN
5jeU0dcUNWsWpOc20LDCfxiCA5GSS/U5SP7muDIkWYG00s+jZXqjXAblvDhEOzeC/C+7kfcvy1r0
qSos4hthPvC1PIGfSsWDqX8CavFbynoseiT4GIgvFneQrT902BlK5+XWbIILaXG8mOArof7JcVNX
XaL302WY9p906Qggoc576c8ImokNLVRZzjVlk4t6QMAc+Ua+J1m9Dfas4erfKSlCvE/qvz1816We
unLD6Ztg5s+4uls07UOxjjaWlKzY84GjC0UpmM0gaHWyZn0qQjCOvQD/4zyGtsxJcCVaDumIiFtI
JCb7fmZUKNjchg/cRaYj3g6w9dKDiNM/UPQsHKoUmoL1cL2HZZs3gsL4YzEbOcFLz+IPv8wdFrJe
2qbQQOhNyxmvohEskTyH4CDadKNbrLWvGpmIEOQMzGWv9RJVqBXm5qOMQZcBmAOhDJ+x6FmUpL1X
H6NOGT5lo5p5qB3nrdDCoW63QOFTts+5JuLgylYeBE/X52L8sGDAoxBWalxV9Sdz1sGFU9B6xm+X
s0MgefD9FKhpeUBxmKRp4MuRW3GAQUb0moAPObjuaQ8rz/5srgNrpnMY+erXxMn0+Z/MUG8II6M1
vdKWaWWJB713pO0VpHs8QhEJzevXdgC+a+iJ0zcQ2/pRhKkRB2BP6btOxYF3x+7DQundSTY8AMpp
uHRk9kq1LhXa2G+iy0X50cA/gt8jaxtt5Hn3ycWlmcr512p8ziboD6oktVlH7XlgqY+xCPc2NhfH
WwRxmFPXelrYgrT8cvhS9Mwi4YpHYiUxThfegTkLh4pcrTpXYVIjjxzV4t87Fj95TdfBJeskUpuR
d52hEvIXk+QCLF/zpwQuXn3KKxTykpePqhe0q3dat2hU6vqPkXxWbViyHuielH6+SpDhWA9uRRlj
W2MAigh+Tg5h8PiH1LBNbUUJne2lUFlsk6CWC8i6jIa5GTReDE/U2WbDmFcaK/kzG27zu+r1ChDC
lr+S+FHwtf65TpMpzPR2KkDhw08HQDLp9MHBjeW0P9DyVSBkuiSGxykxfp3FgsXedQGINOPwGg+8
nx8142PXvnYb6XtNpW30jSZHBzYucSf4m3uthnFpwWuHs53fjJj8tSPXMFXDnqQGGIIVY1ypznVE
1oImeXkzb66B8M1vBZcICx9CQtFiWR2ywLjqk1xjI2U1NkZPWI2KF8FcB4SyYM2ps70uDml13rD4
FutV1/QIN5A/qVt4/Vw3jkFtECklGO4rS6auRY558dTzatdExmwcno3tZL22KbI3mvQXP2RDLxq4
GNymyQ6ekmycSmWS5qQWzphjpPlHUQbkinL5qUIwWQyXzetOWdClZ6M9tf7SXOcWWlHzEpxIQ09V
r+7aDmNjm/z7+I0Gpy2omt5aFrLzgqnCa/3qwgQepFe0h5ddJi+zL3ss9Rvyv9H+heO6cXE/ru/G
RpRkoNfwPTBycdJxnHvoCCMDS1hB+mOa9ajUpglaAWiXcmoaRaYGGy3PHK5cIRWlWW0YemojfbbB
xcDLzTtCTHoaOX5T7id0dFTLfSTivz5TOuuFPyiEmgUl5wvtMCs6X8hf2DQKyTA79yqM2ZL8FBsX
EFMghOtLZ2Qj3RRLAN8lvY8AR8n1/GYlmQ8yO28rCeHuwRlIlchGAQIc/T3/fRN4hICT9oB4o5H4
mO8fXlEPwUUboZQZRYV1yjDKNxUTemR93HWc7IhGLcJSeda2fK9ZW3+T8ijN2SlmpnQsC09KPrFj
WVmXY6lzI/wbDwsJ7Z4+HaTASzMQrmfIjnZRcR4Hc0jY1Ygcbc6r59QnaIl/eMyhs+jcep9Waa3e
mifU0sxoeMjqG08W78RHAWDcnIt+hmwgV8ymwCp6pZbviKGEjilJ02V7J+w8e+e1AT7i3v1CNFpy
7KokqmWtC7H/rGimGDhsTs2qE/5tiTtlU6PlIDEx/4Yapy8CfbbBq5MMPwcLT5OX+d4q0Sh0p5G7
/skfiyyBWB8whzI3WvG7uOSLrXeeXEIUMCKXw//9f1cOIpqyuN0OufBY8Oa+jRhBAhRMA5F2p4K3
ne9Cgmt5uWIKF22tTe/YL7PO0z02G/gXe5E9mcqg8YQI0dWcchncMg/VzZvYXvPT6DmIIJHQIGxn
y7/Ku4gFYNNijXFgPuEAPukc/GaZ6Y8eDRBeacKzOXgYuoG1mcj99S8er89tx7mDlUDcmrO0kTxD
uCYpFU22ynaVxroE2Xl2FiLvzSbZn9x3x686Hyo32iQONxngWCbMKRIgf0MQcq3BVtL0TbcAktn8
p2r+K/6GiHHkgvb+bXnnfQ2UOdJZXhsXAfL7KzwjVhTdzXLkjconbundkcsmo/x/8GD+86XdMvfJ
wuM5b2PiLAwq4/YPKSGleg/G9Xc3B7uH5F1OsfzD6mJ9wPSs5e/n0b+J4fOwwqdRY0mC5QE8txdc
MVPGQmv2XkCmuauHt2k1n7wbg2osf1sovw4v99No811xv2ib1yt9XGIYDCNQPhN80aJGUzrCuZyE
mi3K/nd2pnXaGJ7hc0U9nckmckQC02LSdFR4pc7SUOuIs4BK2w+UwT/JMkN/pd3jzedaSuUE0Ped
plceRgsIOrNZgjF8GCRk1ohvAE7OTBPusgWkeF3OP7rCmqZ3uCqIFx1aSx5/K2u2gAgeGw7QGT0W
14Zb4MfGrGpF3nyMMpyHyrdS+54hoblynapnSIXfYvzgmkSKzA632N7LWqpdlZ38BjgT/FYDTq5U
fG+ZQyKSYZX+XNztGGcIF+xIlVQeJqtyvnLpumBPFtvVbzDvJBK9idaEU8h9Kgiv18BixDsQpqg2
5G4OZg2HjvJr30wHlR3bIu0dkI2Q3pSvMmFGmt2K6ik6kqQpRkHYbaypAnm1lbOvKQM8pX5sFvP4
4A1pCBMf6A9auENqMuDcnkjKmqmAcuGcK/MLJSVxHmdmBiXHDfTJNfmt/ircLCVjwyvyKg32gRMI
bsy93kjxI6qQPGCPvv6lWe87FMKJ/QZbPMdYwaKnF27rcxFol2or0xV/rCsy+oHrrqElzcAbJIT+
s7NFymbOwjpD4H/fORE6Tp8KCspZSWkwZ3ZkDfHWp7YZBrlJymMCJaILs9sSst2QQpYi3LIti1Ai
+cZgbziO8B0JM+GHKn06dL+n3xt+iQcQeNRHZ+QTkSGGw1QBcUXQt5VrJ21XDacbAgC+kj5PjTml
2ueKs3dESlMaAv6Ry0QS8jV2wR8noGO6Wvlubjc0U9gsn0ECD1dCFcDqEcA5H1nCgwNGLaQNFQgc
J8bGtxDiAvBCCWmVxEbvbH6c28/UjBFABHGZWgFHwVgGsATXBR1L1zfmzKQ0Zu/MswAmkDiIN4IF
ZKBlBPwO07lk2WKualt8GVP+rJ2MNf1/nNcHaQs6qnCAxxFTzy9G/svVVGgiSp4jqvJFHmZ/T2+s
zvNGpldP/yJq+pJn5I4e3qIsfZZWjweDfVGi5WJ62OsxJkclDFtHq7DkmsAxnNlVl3eBn+K3xC8B
I0KqYtMuqVFCVlscVZKLlUVsM6+aTOSDCPpXTlcLc0hmDMy3JhNejHgc2SA012ziBNt3vleiRpwj
hbBsrPguA8nOk/8IqmTE1B9//Cu9MGRng/E8OoVXyvEzj9tAYmiGrF+FKntmRJXJHn1uPnFb+8WI
F2ha7qIx2puo04V2JqVGfZGXHgpm9jtts7ddMcBuFlYkLV9m3dMRtsGVIkFteDGUgJoCYtyTm33g
Ufz21LlchXEO6bYwwVoYidIEIlC5LNnL6IlpdoLh1pqYm3Jm9iPgNZ6/6ORBmn45C2tfFdZtXARu
MCxzqCIRI5IHAtR7/SIDBuT8vKxpFqeldw1CUl5R+KaaHXy+i9HoWaNqFgyrXjKu1Eww3F4JZ9Aj
HlU9oOjQSKQ6X+6NT177xfR8E3sI3o0tbDAoNnJVReVLCbRZcnURkQDay75lYqCjEg51NzinNSPT
wcciwFRz6TKzhodRiZNtawRE84/fZBPPEIy0d8/ZrJsjtM564BvxUhOVaQynp9wvZz8DsiaItRhV
5JuDFGz/Xx2sfdy+8hxQffAOHQO9UyIgRbOEVZPisUpbZGi32XzWtSXrDVwAn63VQ3Hk2fzkAPoc
Qw66Q5cL2ZfiIiHjFlCmZVmNXdsHRHhTuEILVbequuqy4m5DWwlv6QLStNp7CjLY1m/5tAuSR7fa
0txMAKOFnzPTdEzjN+Cvt++Onh/aLAEz9RM2+EzmGmK6V53Qv9EmNDU+mWkSf4BQUN7WsdXile39
Xr8xpWI4efSplKxIhJRHjKKFqc2qh13UBUrCe/Cq2p4v9KmCYV1KGLdyu0twvsv6qNEjrNCHuC5E
372mgjZg+rKXawU0QkLrqg1ydeq56HOKfmA2vv5YuQ5sQQmfjmfLQIDYuyeHQjQH4u7rMhelTJqH
nzlbQ4DrGx+GauJj8hW/sriBB2lchORGwoC9MzudRzTN52cVmZEEpYWmLepkvvJnH6FlCf7X88CC
aYfMO2dM1yFGwspJH1Sd5xs4JM7wT3IvOAPEFJ1enmzdmPPa4Oec1oTv+n2GXfkRU6Duh4b2OTjN
K66kZMCMLYoeCxzc+ykHbJJhb/Xhg4nuLGRFwcioXivaaaim+qUEaadqGUG1AYXNcHBmsMsVZ7PD
c/weCI2du/zxs2+4aK/oxJRh9o6tGggefBN3fOfh2EW0APtH5RgiLFJuoivwfuloOktHzk+5FBMU
cka3v8A1xfArE24p9PEDIA36SWttvoQ/nY7QRUd3eOQ4XARzW8+AAQwhApfrZ0uXOtwPdjqSr8ZK
7z8lCm+XNTV7xCnhPy7hhrU0b+aeHy5Go1xcOpJpF/UA/ABiMrMsFoSdWndNRkY2Oq4ewdybsu83
49DtK0fNZ8Ko+zb1Sh6KMrh5SEdyVAzKfJBL1MY0f5x6qBzoiBoaNfqg3MXCtZO1dm9Uc+dgEk/W
hw+qOtlEG/1RCuWTvU+J1sHj3DO3ZKiSjJtJzeE3pE5jkpnT+UFSt8k0Kr7lY+LvCNfr+dR6yKnO
4ohVJg7xXFdb0TNSXj8NAMbefccSoohf8wHPlVugmaPzBF7v0lSlmmnOgOYBPrObnyX399A2mFbp
w7K1sBq6rUWMApV/pzPczYVFm3EcgCr4ke4zuSdpZp0A0Bx6i8K0QKrML/I7d0b+Ec/h7Tqu+QIe
GU5yHZb8QZ+rMG8cWJMG2uzj6uiZ/XZCd+BjGsSqsFnekRG6BD0c3/cQf1YmfF3cWNeGl+xeMUS6
b+BilU306+L8clEhyALfaqYrfHru5pU/pJwNU4ORVCjIlIrVMmhcLP+8FRxE9CfObDmvtTk7fBLo
NXw44OrMsmRpf1gkGEeOQtcvmpuH7+h/X5UvEvaATHC341AmJ63HJlJBjqNOsMZSEtkwaFkObOHs
/lvUpWALGRXqQVjuYxN5a/89hdDC9xVQ7vsqXTNzc6OvovvoXQ22VaWF8u1Tz3qzCqvbS4XMprNB
TRRuMSaqssWY/szT+8DxkFu06HkjFG5EtRkujKoORajeX/P7Xuo8ZGQueFIP8+Jri3FtlkpdmMyC
q4z/BpFqfSpoW4oSEm8e5p7vLVVCZhZdetbs+6+0I6qOZjw+2CmHbHG1E8P44sG87ttQ//pylE65
L92uKEHRxF/YupAaA/KaBExylUhwlxCGLYcaYCsgw2J58rGGX7EozlVhk+WQIPQyzorToCycukRw
+9iJ8EQDoUyOzgWogL4DWeryADIjQQPxjKr8YOPPHk2nzu1PR7Zx/HwJnORgX1zZLbVKWm9nmaqY
TzQXMlW84RTJxv+ouiXxsXeHV1sM9j9KkalL7z+JsvEeP38LrOMkYVFtyJ/eR5A8+JaO372d8CuD
uNsnG86VHpCvkxR1HDsXEFasVVGwdYXQxITXA4NybK2f+aIU3ll+ax5borqnS0lqZ/raLSez5Ym1
grlIRUWZ/w9YFtLjXD1eGCi3ULF7ERC+Rf6XOcQUV5GA0PuS4Ab4w3eyimk2+15wy9SBJ5/79+LN
rqn9hUyodq6HBTpahCeICRDp511NCsmy4WOsr7sjyo2x0TpF19goxDDnCVDK8T4URVO1RPImXIrZ
32PJ9NPzFnVX03NXUPluLrmabMtpOWSm4EjWHT1t5o9Fipp2UqnG6gXZEoE2tff/Db3psp0q8gmG
tcWEcEoVOx+HA+mj1H5mqPIJKS3OfgeTDZoUEFE4JrJTahTUbhf2wzacXNhHkLzzpniRv/Ji5x1y
vo1ukL5LOYUnfYkHpHN3M0q3MWGgmKy4do1G9ZAbMM3CSUdszR7YRGFJH2yXbyHnLs8OzWZ1elrx
b/W5MY9HcIo4a4Q6ab/d5IgSqy++qNL9xcB2paviJUdAmdVfv2yIP+VCw1BcxiTntxQS+DPP+BXO
tk4MqahaV0lqCH+f3vo1kymVE9EYWmw2LkCre9pYH56wvEhzWrR7oHzpVnfRejMDJMVPAh65kQW0
5nZ++H0jbbjaiACguUm/WcIV3H/1h1X2uG7JYlV7kK9oBYfDQ6emStrHCsIgHSbXlKcZ1O4DneZK
EBG/JxabJAZ9nAKYG8hj3vHYIpezY+JX4U/UkRh/qQcIZBdAv3eOfEq2gpXNACzCf847GcR7fvXc
5ANuA7kOWMF2kzJc12fdgVzzJOmTUCgWjqcFjL3pTiMGaF0IWTWzwN33zDjnFquX2+RPjZIsfiop
wdNpLMs83kKSyVLJjKAkmwn0PBNN2N92CUpmawSAnKzgdfutQYEt37xxg5+iJ94yM059D7WxSENS
JNfgldYnDmFopYEKp8W5nT517JlHRWHjzOWGzm/LLIZ+y6wGRhvJH8cZKr+pIKobKCjAMPdL9mTq
1xFCx/+o8jxFZ4r74IE+DAS5E85B9jaH49f+4IZ1vtgyVSlCtRv/ZzfM8mS6pkjC3aVWO/yJu3AS
9e7QUWZIpyJwycQ4A1Fzv3L27clPTcebPCDKurUuR0CHyipTKlV4f0Eiu7aqpJH5oHEw8GxB2cLx
zjBPOTutMIEXvWoAcC/8Wf76fBgiKIGMbmcwmAmwIcaW6igZFN+WbGDSI5/fLiDWnogGFb2Jl/NN
YeOM/UzC7+6vXHluPs8G/NXTamUGVmrqSLdeghvFQf67fVNSwPcEsJosO/xCf/jXeHKIaspm0YRr
gUc5BlgGzZnzJm4n2qJhM0/sVPkZKUTefdz+abVJOJTuidziXLTmADosOqS84JfwWWJZPSSxbmwi
Dp7HnDp7Ljaz3Wh9v1rjI7rW7eLbpHHv9ZKvVkDjEfiohQ/aAFdmJd8PIoRgX00aEBi6ZHaicLSZ
MwxEDPc16SZYxvkzX/UTd8BypHgxrkDTiqnOW3vF+Yk6hX4WHeR7lVhr4yMh9NiC4ImeWrNYlM0n
GHeRe9RUUnbjFytxQcIl8ZR8rkC6ZVzIutAbn0chgxm8tm0dSscA3FFy4OFXAxUJpcLnMmYpcqtT
FyW5cU2jNilSrjEyBrGoK2nmF5UNX1E6z7grdfwm5D+Jq3y5YTxvootP4H0bv6u+rU8uqbNLyKgD
+wZPHgUfq3YSjzRv9ieIea6BSDmRYNFeSuUUbSz3aagjYTKSYdouiiE9TaWHnBgCkf1ezX7kps33
ui/ZXWPOkO6FGvxNOanovG6SegmeW43gkA5Zs5NkYl5F5m3Aw4kvhtDfd+rFffT5JGL24b4LWyMK
zuhw3hvLp3DfXPXMm2Ku2hnAdkekGzpFAskJJ5uPnso5NAGeZsRHlgWfULzWDBwPmZCJQeXHu939
b08OMT6WW6GGZAx4z/pBZ02DDZ2wRav0yshr9oEI8KZ0aEgaGjCooxC4YCIyp51EaxpO2Z4ytmqp
HVFE7VMx79vWnjYtGkIMkDJdbPp8EfAlhwvpH78V5nswCrxA7FqwE7ah4ERzrKMLHMb7o8+Rcm/K
jCEfiR7aJITJ+KOYywSf7icWLrBIj5o/id78CqSNzH6iEJw+Qx8HMUyG1WwiBy5A6MgKTpFI+vz5
RDXWpKzDg86agNJbwiUB319pPkY1MZLirSLSwZMRJfGySmP9CfVy9/qZqKU8a4jVQvpAFJkdrkzf
O/IfMNH/kb38agd4krsl5asmn2A8sCUHR67kpw4UorcD4MEz5QbQztAQ3ZrH2utDN5W+smSFdGO8
Fgl68eIieMvOCx1S72A/cC8yit+H3FXGzXDYSNYKDnehBRVPuv0MeXUTBCMW7r4APE0iNaeCT65D
tmb+jdzpmQcKXIy+gt43I28KfFIfMwWaLbMtN77QL5Gg8rGNp2zddenmWJS3MrrM6mH/V5+Ckuoi
tUv9GxL7H79kTZE4WH0saqSd2nABs+KT0N5wnQ0drE3qSSvbv9cykUc0sk3ozrQlMkeYC8C46KBx
hlljXMaJsmSSuPNfQKpTyVazAMxOvRPv0+jV/FFwjQNGSmqAmLKBLoq/K5Ubvdrp+Wi7TN/ecGft
nc5QNnTkIcn4+DdfUr42Nkl8BVOvqPKQxmyazJ59srM0ibBY+XOmuQjT3CxQOma8NcpjtDJqQyLw
UBi3I8Wmc82Uhi/3VG0+CCQkCtH+eKCm200goU51F1LM6L1yITWb0tFM0h19wgorcGU7uXY2GCf3
j//JO85NWlsw6INFb7rfGQ5+Ns/FMhTvfsnJXHRcp8c2RLNFxPKUqM0Y4xOnYxFuSRkn1TEgt7fa
4TWzf/HQ2IsKwyvLR//SeSSJvhsR366lTdMJB3nSVvxsCBG7V/Kjc/Xob7CzVcsSLH+4YX0q9Eo8
K5gGtg3HXWGh6k5IjU+7bWOjpywBgX54+mC9kGdVTn79w+A400B+uRFRlXMVX3P8e8g+NBtsz9ea
VIbp/404LVrQhVeD1TOxCYvfj/yX5cpKnTwGBSMGYUMcz+fIcT3lH8ddqkpHmSdOqUdkA+q/XKUQ
J735D/EnoZ1jcyahPXBNBN8/gcbIbyomRJIKsEXtzV6jurs0CDAImJkZtnHI5NMe2VaxtcxZSghc
9aKdEDEJ7df9fTl5Tfnpa/Ag1rMIQyeCa8ED7P9wce1BWMdqeBm1k6AQvOvNsaKHC/WADKGb153J
+S1k+FYy/Ru2P8csKyh8QcusjSgPbf+E/Y54OXt8ZoI2a2YSW37wGzTCMq0mfKoxXGf5JalBymV8
nkQV5exCVRe4ltdxyfQ9zFtZihiuPbIoD938TyzkwAS+7pObzqNLuoLkS80BvDkajO58Dewqpzfz
APBKBN+TX8PiGWqQghv43cGi57omRwrBuKFDlRjP+Ryyhe/B3VgAY327pBkHYjCeRxyudxM7ld0c
7D/Voqi1yNqnVhuPI18dx3J4Lc4Fj+jI3hvlqh8agW8/UmQt4MVQyjUab/TXcCOtM5iI4hsSeLmC
HtGMfxzDGD3oCedWv65xsZKlDnGRsBYmMOu8Uue98Qxs3nJI6elNELQ98+MW1p88aWsHV//3my5e
G+80ENkeVKGo7xvfC28qpT2EW2PI8vh4G5uS1+87G9ZFSkv7PQtWbLBtKrolCr5NBvqyMZF9ReQN
Umh8Xz9Ws0npLfeZ6Bour3eFCPN8pqJ4aihUwGWefWcOU2lBpAPd9ZQ+UwEzg2mBRluGAupZxxXc
/aY2WNzf140FCbthgc76+sZWwShpzpnmcb7pvbhHOUUpTrSPCAMj6uAiqVFDNK1JR3yA2CbUXblk
xsSXdY2PwXYOiNjF3GBOtC2c+bFsWhB9jT2hoiFSBMQrdEVT4j696o7WUVmQnzHQzLWGiPJ7DtY+
LIcWLyK98+C+2xGctyKu/8Jv9r5p0arfRejieG48DNixSmpZuAD6TEVd3qDpP6UoTl+dxhphG08e
6geCHrGj5gnyMAF3CC28YR7SD2DeTGM1o1vGPIVUdHjGwglENVQ3WXpm1ELiAXLnLchPydVGLA0Z
QAbh9aeJjGsYvPuj3bTgjWMljPxPlraJ0GJPnpIia/rNG0vq/cc2URY30AFvjbsdIULYD8EEG0oZ
nFciJBPGQk0TPLfPU04AJ8Y9npcaFQFAmj8yc7B+Smrictg1pCP+ylWtGL/mK0BuyCa564dYpykT
sbGpC7H46A6kHcDyNVlhqhETW9iTpSnnNDCAF6cTQrL0kOCC0xlp71YjWzN2ofNR5V8vDM7FL05p
2hVD/xHqy/zaBNnBakNNrgMvDWJoXjD6q7+XVMkzjHDtpePfBQvjygTF0wAjoHhFxnl2exWAoPik
J1yxKN/tkoJ/ZuFLZh5XpOd+oHJ4cYAS7tvu15nGKiu1RkQ1jW78jcRokmFl46qfjW5iT1UvjU/O
BTuMCIBYdGvEOTjNlwNpmBffjRPQI/efefTDny+aAVRvi5WP3IhSfurbr0rnHC3jNadMSseWw6QX
nraLQE0MRQcVPQVDCtb1w1qH9sJ0F7LhDMefaMPb8ycqkyunfl+Z3KtsYf85fqO9t9hZXwtqfKlZ
nIgqb7tOF96AEbEmt4J6D5hfaL2kXWmhxMjGX59NfOPV4JW1jowzFnBHgP9rVE45WX3WAN6GYCaj
5yQ9Xc3lBjd+YUp7dscJyC1wMASLQnmJNm0TB471aaoQi47Eda4EF2BgfZ/NK5ZB6OD6rygloz7c
a1X43/EYHXXvR+/GDmjUlUQfa5nLdbLOBDNJWFJRCZMYJgL/quVELxeDQt9qdoXMmOr5IuPRTE1A
0788G9/Tzg8zoasw5a/5ZRxyW4Fpheqx/C3HgqNL4NATqDmOYvwk1XxHVgxLtZlywO0kX03R/87o
x1oujaxV8Chi/t0VHan3nipLrlBpkuteVT1pVK5ZCpWbThdOSiUBPBisNmXbIQtg9oJU0MizPj1W
wBRFrn2IQPdMYhPu9b8ahSUxSfzZtD8RzPduFk+lQ7j4H3fU/9wdEPC8eRHJopvO2TMytlahFPyM
HFo2ttFl1BRj+MG+wFH9AI/FRQLII43nXJzpEduRgASysV8dnMt7s4ABDnG5+kJoHC46JVaNlvJg
b4qNmF41LIMIAlrPI2BBNfQ70ob+cU6ZaCGpPR5VzTXPVcCt5Qyd7sJRndnzg8O8TAWVz3yHzsjt
EvUgQe/hf/1/6j+IAmcCR8Q63OIyDm1+Or4X0TgY6b1YtXLmhqdaW2IdRAGRowl1buxo66zOYddU
0jkRTJmn3U2EYYecxksKea2rPuec6bpv28Sl+LDu5rktX+8Ilp5P77gSuyDkVeavXcJJQwGofMnk
q6V/4xCHgjBJRMDcEH+kO2DzO9RVPd2UT5LLgtbu4T6/XwHK90QELkKdQbnbEov0yV3gB2/1xz2j
Rrw22TkjBzT/011wAa7rbmL+EngJbBPbm4+r7sMJtaX7tkrXGEp0TviYnStHjU8pHJgfAp2iOukZ
NP8SwiNcNc9ZGNnoafhJ/4PwLzrGplDyDJkDYXO0qkVXum331WOgUweVoDQeFj9zinuPgOJsSPqA
hrDXNb2yXaUngC1AdUUiDi43QFDAAx+TQs99leGOgAiW5GW0cIuMDVr1DwBpNVAYPvfgMMEre1k1
7kLmgpk8pDN2QHbpyJVWFcYGLSAa0ImVx5RYbfloS3q+uCIi4yBE7iteoHtET7D880vuloLO8DJj
BHV+QouFAmN2QOwYplXwUjuAaMejjvsCz29wKQ0dpS5UkaDooWXQO4rAkj39P28MED1mwVcUcILp
EBnZ6YYKS9KYNfEHHZEqM0nwjpDaBeh36cNUl0v0+HXwQVh+gy3lzUCf/Wa8McRyWus1altwnGXO
rThSth1w9x/LE8JSmUyAw86217XifWa2TCf39vgPt8Ds5zQ66godV3YsmJW2zroXuOM6couBtX9R
TSAmCUIlGaMG2cd8y0iKwPYqoVIP2cWFwYlh4ZI4ckk7cjSGILEYe1f7tSZPJIIxdlVESM5s9fhM
dvXn/OMFgJOEjPlEXBdcSjK9jLf+AMZuTx1atkG1tHi5Bwxh1AmIqc6/RhSoQilBihRY9tuchmhJ
7jVv2cf3ufKUDP8Vy6X5z2aj1+QCtZY9qLN74HIQOlZ3tCAzixc3b1xuyPYobWl7O9WM3GWZlVe8
MwxBLOVvTUN/78qSB5QhZp9slslcRMsLt1N4iTjM4eqz002PKhPMEWOFxhOJiLaYKVWprQFcLIki
b3REggIhsRlGToy+b/XjW92/wqTM/7JAh/sIo+A67sat1O7j4LxlWA1KLLwmgWRytWEvQ0rTDzIF
XPOFbGFdjHDTLNdwju8HcDYhpGS8F0Ra66RdzMGVTqFz0wh+Ly9bLZHU/4loWHh2Z9XUePKjtvYO
kVWLC8AbgYJRmIxdbwAtcSexynqLoSWmb+12gKl9/yKZKYqetlafmUEVASyUGN5RclVXZ4CHRrbQ
XB+OBJrZsFLy4HHL9K4x0RyMsbuctvr2tGCCt/NOo7/6nRES2mr5C3enXPNW6rLjBE15HbFHXppZ
PSKRyWIXy45Qbau2uRtbZZnqmgG93gp0sahcpxntE49rh0WwmtV3OwaG4UJdET2JWEvFxVyn2eRY
IhA/RJ+z0YA0rjcsQ3fe5a7J38d07lLPLaJOYhZDRpekz2ZckW3/hjxTLI3AXihj/mXRjrEjKOHN
meRHneGyFzgx6h91zcqJYk2WjO7lvvjxDDIYJPSAx8uS2Cf7v+LXS1RBVc0OfgHXwjG71EJB3FCz
H6uiDw3+kYdkXdaSN6lRbZiYEwVeaRjBjW2222bijQ+oOHkKkpUqE+7rOPPTDW8ibO+LBSFDLqwo
uOrHonTsYlq/JfNYj6cnp8MMwD9XhNupGiPzBvr0DzQOqKuY0ZhTDWVRUA/HMiKWWfsGD1xvA/1f
qFcYS674sXp82z9JxaFYUzquDEhbBMk1Ju8o3vhekN5Gr+lUMGVcfsybUsa7nHfcEksVOeqwL8hM
SPVTJ6inthQ1Kt7xUPOMKQLQCy361zfV2JEREQvTgk0I3nWIk7wIxTkvT8nwskStUfawPfvn8np9
7GiBl3FW3xTfLmkO0u2RPgbl5K6OxzT543NZrTglq1FZk53bY0w9I2Ax8KNZRPdixH9TDvlQxRx4
seXmNkqRcwJQymtQzYKs0BcX8jrXPHXa/88oy5oiU6OtO0U4k6ZP4cukVVwkFDD4F5ERewJdMMKO
OvYnMbVAk45RbOT3g1txJHutFJjZ8Rgcz3DY/TFTZC8EqPm3Z/+7yM1YT+xu8cfNgJTNOCPlv3FG
zbNGp22px8lk7lRmPtxi7K3mIHReaRpGDn1azIP4N3itHiih9C1m2k28K7yDtEurhuEFimV2a4/L
NcrvnX3UxkfJZd0uRqVKCqAk2NTiH2Vr98vfhL+TVqGY4ZO/dcneaa13NcuneMzaYF+93d/zaRxf
a20UmcbWqD4r2txlo9xj9nszx3NtkqpbAzkYud8Q5xkjN9oyX/VpAhpU+Yzp6YgDWyvO1QYWA0TP
WZzL82/kjEyIalSFoNB4G2PxKPuhBUYvDEpiGreH2HHqyKSJ5823/4oCJRmf7EJv7gki7+fb9YYV
oyQThhJtfs9O7Of0DYkVsYtcIPF9tE9CVUbOul5fLS8nswrQhd0/HaveIfPkTHnTQJ8vM4jx+D+n
NwknO9mIl5Uf8q5x2mcCEkExX0WvWHdlqnCJM1fP3/3fBCwoIu7byv8bsm9QQn/v1IprxNeENO1E
uzO1se5Eh/modJnz954NQjB2wSOU3QyK3VEGqnPGLiuvKD9koQFgXMcZb1m1xzx1G/4r+dPBJWDl
AvgWUCCMGW7ZObpGWUosAQZleU6WkkuvQmweZ9frScCq6iLMI8HmRSa5wvWwQWjCGES/598zTphd
xCCMrzvYVjDBVUWY+QIpwGU26PA3g4zX+3uuJXDvPH2h/AqZzj7BHhiutlqFImOO+paRXrD/7UOu
ynd3jwPyBevHIHXglh+hCumQWiRoIl1hLwABzRQH/UH1S0O9Nbie2JhMSf+RRVXHVGmiEZYuFNag
twjRpyghdr5PmWSd14dukFVZrheuqXJr15RV63jw17AGL1GhHBtSTZWUwzqccozwlhCexDpTegdk
LVR9ISlLG1mdOi+NgDZBfcqzIcThHucM4ifb/y/yZ2AMseTkSaQVuWgLNA8p544Be0IaBXWalobS
8nmxkJYTmowPh+2hK7AKnogFcPl9/glgAlDvIjaKPWc1zedrArcdui1SAoQRD9vNPBUD2wxflhJN
6gBfE0G3uCgmQ+0/9OJq9+FTjO5DhhHaUcWNjppJrFq5GhfLmKXpxl75c3wIuPlebfWP/SpA6GRW
EyAHA07tZpO3j636QFTyuNCBKIR8MOQGy97h6AGxclmQDQ5/MObHUQbhBsbb+55/zubYhI/T3zYy
qImGM37cFM34rsIFzezR8UK/gemV6kgolq83kbQ/bnW69CaLu033VKvkEA7aA5uv6JRRFympJaFK
rnKZCz9PcgzxjnP4v6nUtt1QuAY5/aa/wH9/Dt2B/aAZdYdo6UWdKJd8T3kJmHrpawP91PUBcQ/v
MYT7dhqULNXprSf46Pqo7b45B4NyNHS7LaTiwtZXqmRqwCu/WDeIhQCd5On4OnOvqhnfb2UpN143
WApqjzmJdNBzTLihinPG88XsTdQUAMl/V9TZQAwVmJ8LhtXwqG9yABfFY1sMV9bkRLQPRO3v4WT4
RGmUDNgD6rMNrp2AMg8ZY6eT1YqIqGOpgbMtgLm1mXlGItkoFUESM11D++lFOcW9dSk9GNwqtuA5
fbgHvUEBOOUouyxCAimJoMbln6KiILPVMFfvocgwHRMvd/rYkcxwwxPPYPM2huB/1lMyUsgagCf2
S2E9a0qikTwhqv8X3C6JwLHY59dPUPXwq/C4Yx/Nm66Y/VktgAORnPOFKsFGfvnFgNrMB2DeI7yV
HBNUtlSpVY1f0YPo2QAtgI00uTo0SeRS9IApAz2q2wEi7emSGubiq30l1NlbYS/8scbY4NdCN/2z
QnNvdB3r7/vp4L+Oja9GNouTgq0gAClgaNeNdUQ/PF+hjapShH7U3vAK2QhDXMQ5JrxNnGsAN+N7
q2f9Q8M1nwOngU8yFLtNsmpCDWvA0gyBOkC8R9koRoiINzRoawbuVOIrqEL6y3PPXKR+vrlrSzjm
Vr5Lxkp5kwHrK/uqw87IF0EFJsbABa/voosiVC7FtHHcR6nscZBBkmAdCWPUJRGNpINkRn8X9ETk
F9tFUCF3p2pmX0rNC6A8stErQTdqFk30yqLbrtYCKNlDs7te6peQoRAEQLCRXjguoBHG0z2x7B/g
NJye9221+47ACZNqYhic2HQxfCgNq2DLaQL3oAta5ygmftQ/Vkf5kdrQXBvarDsw5pbgVvA/2f83
oNJlRctjybswJe2f0uRsuZtF4Yfk0NiPnuIPO4QmhqHJ8f1rRP9PGg5uYScJue+L37YgCJVP9f3k
bDtuwkTooSt9LaJ5MH6+esOlkfunMNre+rO9PIsdmGD/aQ3Ijl1rdg/gMcWD9+FeJFW4LYtXVJO+
+YlD13p8OZmMCvhnpiW/grrPTIWnS/dMvSutIO87eko+JmfLrfmTuKg5qDQMQ5I1Oc/2Hg2R1jgj
yey9DO2swCNhdjP8Vx0ABkEPjrQR57aT9eodmm0LkHE3ySIzSuh0AoV1pL09eJhWn6DhkSox7pwt
ZdBTrmnQ2+qKJdZa+NyqYdeaJK6tLNOUGDTOBsS7WjUK2gUnpGvLH/s3nTzva7X5HZqqCXTBeuZr
F8nHnhSSElH+/6L/S4O2bzO9+HENRDUHYplpbknMKBifX7VslX/0QZDs32K2GQ7V1eg7XmNMXqLb
kmG5aE6YFp5boSYnSbWZ0qVb2hqw2K4gUcXU/zyoHXliFhzA0gWNSSNJOrLYZBdruLi7mmjlUrn5
GIc0OKDT7qPn5QvA6RaYybSsmASG+KsPe4i2HvnxEDUnLxa0ePsSMCcyAmQnWUI3OiFhi3+rRflO
NEnVOedNIW8ThatrawToA8bLHJ0to9XbO+w1zNvKS0WXTFL/k3sYFMgjd7trBkQg2yxUnQ75LA/S
VZD2rgdZjJZLsFY0MO6QfvUHauMgxPHZzCAkCfj4u3XhBYNE8ZVU9t2r2efgR61zVhA47q4QvNBZ
augy8cY9DLtCHadowRfsMm4qE/jNJEQggbwqZop3gYkAvbLiupMVve07UyzT35fwPr8Gg/FA+eWP
Jy3kUg2Tvp5NymDEi56QmJM4TftXt8BL2EJ1gGvGgr1bsX8xWDulJqEvfRzadH4UDq2WDaTet1u2
xTLBNT2us4c+H7yX71ZMkgL1vKidUV10YLCnbd5RkiSH7ylmTulCJeapNOsljVFEEIokOQUuoBK0
HTIf/b8Q3nt7KanTj+SoJ3ODbQXe5aksH2jT6ztUYB+6zukzu0zaBhKqScBAu4jGkCbiCPtNXwlP
VhTboUr92ZoUpIDxY6AzGs9utt5y2Y6tvHtutws6J3kSsQxYhXdoM1NSahuCEK9QarAP1cdvZ0rr
2MjWQk/8CgFqdutbkH+SRQaDAo2KisLScFf4gckoq1bVhkP9bLvPszaE4evfAFTCq69QdtRuFZ7c
BFhtre5Qn2vnHnKM5V7YsXRATM6rWd3kDPY7iO4k4RNGtEnavbKtfo7+WsTOxxL4/jlqZYcMkOwJ
YBfj9OziA4i12QEg+5OdxtDTRgZ0nTcg2gZCZwbo6unu2NCv0xJyhqIEcnwP4G3G2MC6re8nx2Kh
4G20jD7K6ngW4Q3CLNN2bOdaUPTyfqym8BncB0aMDwzhuGeA7jyoFD/6FaGIUn9WDYiadS/QKH7J
ESGtbHkc3RSU0/Twm8dJGZ2Mx8v7odT5Kt4VlzZPQ7ciT7WsdNPtoDHRnp5NN7xEjQEhTcjsFr1H
6wOAuWvy22CFKkIvYJA5bLpMOGoSBIThPrcsG163JoWXxdX9XL9RrpYP00kjiF0jfQbKVV5Q0Dpm
Kq3ORv3RdWbryHet/8tBaWV+BgyJXkpp51pzpF36iMWEh4TxyqWyzD5BMowXBOexP3Ecaz0PZRvf
lWrqNeRcSHoxSPFG1RkSi/1KL/1bds58WggZnycIinrCo3KyTbSFtCfViDe6GCauwBGfoAJYocsW
+VN3flwywIXrnEfyEMQ6Za3dw4BOfNaiEMwD1S1WzCDKGwnhZvj29TdhGCBZraSlh9p0VdjIrA+M
i/sLrvYWOURl78BYhUt2TNqzOjSUM8d/wrOrhYfhxVynLRgi1J2mc07a8Q9aat3Y98shyzPqlyAM
eABnd9o9X1QeET/go/5pqoiHwQUR4/wPDaotv6+hZDjrrzUKY5mU54iExwZL165LqaPkYkQFetzy
8NYbYBwQOnxClg4vuUnUk15ZTjXoy5ovuRyzi5CWD8mUwHLi0nVYelB6lg97EcooeMxk49cHTXCp
TmXSQg9A3mU5FxfMPBdukkAL99cFkXE+iGV3EuDv+nMrC2DhSylbwbfg7FynszXaIyAHLQhYmJVQ
Wf4B2WeXjieEIc8GjW7lspB91MDngwZhzQBBpkQqOVEnk0LStNI4n/F5JUH84ICGkAiSvXq1oozx
ZACJhgSR11pQ2co4FGLvsBl2DpXuozqJRmJyO+w6oYK0oeCzDzA82yA5F30ZpC5BwaSvouzb2Bll
JWQ77JKLYkTC/XMed17bQrEEHqBZLYNJ06xg3BEhPpT8V7X350VxAX0JrhvharrDOYqp87LJXoKe
Ih/0YVuokwJgt9Nh5IGwf6x+GaAD+YglkX7WjgJXaeBNMOkPhxfRcZ8Bfqvf3Ov3Tbv01ldq+3/K
f+P8fp88DzwdiRBKriRO9l8KDizq51t7U7Yq3TrfUs/zY3NgWzfX6UNcisoF3XbXPtLBy5uTud/h
EL4kpLxJWILG7ZwGxfM4oFOeK3J9+yK1fep6JV6Y2K/bEpjfLHfuIdHTfBBMMICLciybp7CkAqzr
0/e7ZwkWlR+jA5Lu0SIcmBCVjoXVM+HU8ZF/kizdFB8pLFk1H1g2yV1rXsIt0B3jwi1WJ2Por/Em
wtAm8z8cOIubZ0NvJiJlwNDZCDrWxvZK+yknzMEib7Tbkk6TPIWxsYgMDv3zCA4PIbectcxkQhXP
+eNUmE7lhFgXuaLAMP5u2nxiTtn3K8hoByxTv8H8CWUEDnaKGOgV9b7nvXVRFdx+fCb+1cL4H/qq
Y+dQchYUyvSanONYIC+NcazNcSuujfOjzFXV6azrwmuIQKyuTZ42DZXX+XThG0qTnVCToI4+4sOo
rQANrQBNTPP9KKdmqEz1guoSvaIZON8f2vie9LkDeFzK9qIsnYOO8iFY6JBOLAo4fEz+FPwrPS0k
8ccz/76RKTRkkgCtMAp/KxJqLFltf0BXNk6e0ENbEYnJMJwHInw6oOxlZTpMNFDnmdHvM+8WVMXQ
L/RhcbMM1cs43hbQbFx38UFaM2F5KI3H2TpudQzktVrS/VJUef5QDuVkibWbsd6Vh08NsGG1FAcP
IJ8zEpORqabRTMiF7QoQbWpd0f/9oHHGnZkvJJKs0/yfOhfUzRDEaekMm2dzqAVaxXj2OHUXM1X0
ErzcWmworQpr/WMW51vOlKz0hBwZ7vkTQIMsqNxGZ73Y58zguExgBBAY+5218Y89ccqsEav+No2y
Fkm1rWhmLklVy9A4jzQzRjf9D5sBPHYcIVPkCbHnshAFgT/200hDkk8BTbtfxSDFxFSI/V0M4nj+
uBLFc6ra+D0e7Z/NxpxB1Vb569D5pPaj2nCEvFlLSMheY4YeBCfVuARXXnjnxrJPq7kVK7oHkm7H
/BGsymXRZqf8mgVEUZYqTtMo45agi0N5PBp9ejnm7UB1Xp0uXemkVAWRFPsPo0fI8v8VV6XYeCcc
VnxAR6PSAeRiI96givcK0LWTeB2i3tcP9ZenSHufvIYaebNc81FKTUEHsmlKzzhwfgEErLf50JGH
SNGvgQhiqfdau+dQExDf8gzQzGsYTJoXC1hqeeJeC8XA4wIfQvu8F6Je+9tltJvVEd3aBufY1s27
TWNzJJCuUPGjxX+hwiozNl5FL3p6Co8veDsULmJOl0LVvuSFiWEgil0AQ8lIJl365/Q/AG5ISeqm
iYEEz9e7R8OZYUMWyfiL15EKv0hM0JNMkfhAR4lxDLP4xuNXQIDp5hjWOd7uzXBx8ttm5pT1OkxY
3BI2DDG1gz0IXaugWTsD3A/gYZhvTzQoGtYrF9OMx7qEM076Jx4eeK+R1Qf1O/uINd1PiLjYLXeU
xwVRzLBPbHRacTzqaGTi4AREqjHD3+0phoa21yWz9ag+Gl4F3XuBl4c1lEoeLyB85MrJIQEXcwJ1
YDfoYXqh5gs6En7Kj1g487NBgPC6+TeQy5dQFvsgrvwjOQeBPqngiU+jWsp68TbdDZuOK/snWyX7
4x7uQ3TmL3Rq7EsGkQdHAvC9noJbnhbw41JAaiZwaTmoAWl/albWTOhDt1N6wmP59q/RQhn0q5Le
SE1ZIpQ+YyFtmdJY/uOPA4EUrjfhZm1xvgz+GwKU62bZbpj62QR2rr4ou46g2pFN2ZfrMU8nPeVm
2aGByC/+C+BaJST5BY+SMLCPvGpbt9ajOoB7vP6lYiCdMDDo20kTbA8aUbYI1GfZGKnkTfkvev3J
tKQHoJ1KfJVljkrC2+MDTnL70v5b7qvE4q3bcfyA4oldKVy48kJ1mOZGXTB8jwtB8hUDSvILjgDH
hS8e1VD6i9CnlTeAGrQ1Y9nYKWud3RTt5321pL4jfH27ltakOhfYYyVfJbMiI/ZX/O559CHdnBMo
ZUe9zVIlSsns31/AwqdsYF5GTuStZSXkDC9JkrBm6umwPw/EWjnaUyQLuko+L4/b8FPXv32qakOd
Ull881CcUS1xLIo09tOlZ1tIb3e7gR3knHDGAdZWpmxYhGGVPK0YxIgWwzyh87jaUcyQIIipxq/E
jxtplBw6oLvm124Zf9dCr0bdxQDaXW6sxXX4Tqj75WDI0Ze4Gqlltl6P3QN61UACKJYHFjdt8gQI
sv/YoJHQDlBQkPwRt5eJtqeuTwVYzrgw0gz++WLOKnLdSGPTSgZMGwsbtTyo5UXQVT1V+EZlQ+YW
/s5p649POXtVxIrBJGeK6YcGZ+7gU2r7kljQLeLngb5yDfR/oSr1wN6ClXw6OTnL9jDLskzHd+d/
Chniydq+gkLDP8W7M6n/gSQKqsRHSD0fL7p9NIA0elrwLqMxQC2tRdYbbqAuBzXe9v3LrVGSPrxt
zoNYL9CFfkdJh6zPEhiOt9lwjLQZ4zzXhFxsy4YxJz8JxXWvgPB8WOt/jSJi2elVk7dc+AWhNrjk
yiyVcfOKux52endG0DcLPCQLxdiX0oVTQU74vmXcqdqq8lmCulf2+ngux74LoHQDPIg0nq9AmwkQ
yMfnR8yTFseIi4WTy6Hg4gBzFKtLFCIzGu25qHnUni3V/M1B/hX/CAOl4By20gJ+CnWE5uTGRn5z
awJOYdGV/oN7GjUxHQVc4ijGXfQL3IP2AnB1HtxeuEg9NLwqfHj04FttXXeOg+9NXDMRcnRJ8ynt
T2xJjpTn7RFgbaX6xGmO+ckWOWQxywPo2+wcyHtgbAnPT+zzrSKdmDPTl2M0Z/FWKmy7qF1AOmfJ
K2riv52vR0sJdXr/2YwbQnv+1Zet81YLCsFStWT0pYIiPY7mRTZzow3TMbGLRPOIZO1BMvD13dbn
76niPtW6ytgT6teIkzxP7NntU4HuUISFBWtBsHcW+NMrHE/o+AYQ3by5Xqib1JCzz39kyUDy2bLK
o+nnWuj4LwwEcC8JjcuI+GmnQd9XgrCuHlGxVJxHc8OhEZL9tVTjGmIbMlfIGQYyxUnV0UEz7Wcq
0VRpQXOw9neo52a4+ImxulAPxGO4LBLq+R5YiXJYNab5yywW44ApKSB2wo22+pO3Jke7rM3lBey2
mcGAfvsN2Zzn3UeybMBGwzfUUC2SXwIrGHuGpVmdRsyNwthRIxIVWFaBBjQQk4MKGMBfeYu/mh+T
LMEfuBBuX/3xrlQIRzfg3xxJJgRKCuTt0eFY2BE89r2zM1tnUjIksBuJPUAreFH8rS/2Nt2NORkq
D9Nj3CoKQOuEb4AObC4WquoOphmAGJgwBow6Ir7fCMHPXCWd6SR7sCvi0wDxElZACHM/IQtsCgNl
pbI0TkqX0ThjSyrSSgxnqZqrRN+qiLjfDkbd+IiXVQzE3goA0v6r1B+0wsH8h/ZueA3qgGpLmTmq
0jCl3omrHXrhA+ejrESizFcsm9iTihlWzslTdlfJ42J/+KQ/1/nVLuussn/6QdsSOkbmsGPGqZXC
6h550TjgtKT+qxCTNCsuiP6cuLraa42wn0YAy23Jx51WvKpCAUlubGeCL1wncJrSo4weseRKNyLo
Bh5P8UremzFTK7aaJxTUxreFgE9Em09agx48DjhD7Dmxr8nSruH5jSUrPzWtMW/W4xseQALCrjRp
9GE5varXWpGOKiZ5P1O8XU3M2C7ZP8d4hMfFw691FLDY+oz3osArSXUXuX/uQtP3+OFrhjgo9GTl
w6+mppboh7zwvJbaPVxpDoasADhlGFqRR5U7GodDztDqeP/pPT+xXp7zfyeO2hQJOD4oDVuW/7lC
PVvLOeFuGngEnfYEGXoN2N1trpUT84VQlwEpM72sj+rh3hBWH9kW4xCCjJzPpZ7nEagr9IO8lQa8
j3FKnkpENb1mKXAzC9WNjMumiJDyzfCj0iFGHoYvs8wQllkLp8/EiT0rPQVKZNFp+RAAobyw4g2f
a7qDakeEfDgwHceOm5ZNZkmMcU4CY3KlMyXfchasz175W2gSqJpkNG+UV8rb9YgVXNP1f4CmGRX2
D3zJyrThKg+mO29G6WmpVv8aDjCD99dgf1olIFwvQIGhHSjzB9ST5nMVN+eTagjPn0LXPFe2oiio
mi2yTTlAVLV+Q+YcR+k1tu9RHYv1N3fWyQtVUpcNrTaYiruJ+GL7l0tMT//lXOzBS0pwNxwzlGkB
zD3LmTDUdLu1iygPOECOb27aDse1EzjP+MdJLrnDhPOhTQightOxUi+PiOvJR/ozALdRi0OaijtV
J0PGxn3eDjlzh81FkK6QCKCoLbbmgmtzviKgoMVZD/rBZP1s++2S1nXDVneUzEIYjYPgohaU4/CK
jBiC3B1lZN4qBZpY/+0Tg82RXpquoeXJL+KF+rS3fOzoeXUDG4N+zi84OAw+NoXqsYI7ZYL1wUGp
T7DdulgVQljWGCPWMPQEuRCMuWB8g7LOfQKNE3yStTkcoAamGxM8uRE+N2eAvHC/Fqz3f72dGaYX
UM0dNUFf3/MZykUhgvh7yopBbWFV8FGcaP1BzrlTdq6iIU7h3FrlzoI69eNaImBcl9KF7Uyyww37
8vPj/Jby1yfbQUtolFhFrEkSQr5bBOt3QbAcXrPZ1dtyKSWd6wiOoH7wz7E3cgQklJ23jqFeOIgC
tfabTGLr24R8RqVp/Qad78ENE4veJ35h1kkzONZAZDtwvEzOhYYQJS46c5He5AWh6hh+e9ECpooz
lLLxFdGdcpxzOVnSdfmjLa5vmDE4P+F6VISekto1gOI7EpeOsD4d0rRw1HPU19JWLg47BkpQsNGu
N45mOEiBw7vSI6Dz5Rk55wudQs1ZIqK4TUhtu/NEgJfDQ+j+pc+W9YuQUWmEvgD/o7Cbk2jmh6Gt
2GRD20e6mjoVYh/qfycpvolr1JW1rCy7QcWhGqtZJblaNof4c0BdrbADmovggB3a/kyBY+Mg8xmp
xCtwEy/feVLDfdD46s9SHeKMPoIZm3HCPCLmzAGmvzI7vRJp0Lz1NbA9eMKD7UOelo57q7M3maMz
gtJX+aS+jsI5vJPK/HjR2C8bQLR29M0JTgxeMlGYw48WSmxsffKYhTDrNtkiONbCLAdKU0ujysYy
3hdSQB6/YPCgOhxKHBFwEQ5gIvQsV1sWHRqzG4VjKg8V3Nu1PqXmEKpr9H/5aagUm2k5IQ1sRJkZ
L0oHSamDI8+EqBrFOb/gtW8Wgc2vNxZZZ2A1QEuCF78iBU+nhVo3pmrsnaLjhSpKbw3px3xB5cqc
Ek5Gdz1mrewG06QR2PD5/tMwJmDc57EMbac3jYqnEIuaZQtlh3Twm/Q0bE1GrI4I3sYW9+omLslo
pAKmnbfUCnh6644AhzmlVrb7+ZwjW/WgSrfYsddCgQ8lnU8UgwletVfTAQ/hdvRuBF0DFYcqE8mN
4vxT64MOvBrH1/7yuifqVXyeT1BluFg7lteM4i3ma8aAJtmeNyDZytoDD+NK/vja9YCxvH3ISws0
0KOsY3sB9uit/pM9/JbedaJYBaKUaMvU10sYFYTNV1EicdbfWfB+/qvme5zqH54vIwO08Y6x4O5s
bf3peOiETFQ/Du0BUWJWkYJ7aFpC/k00wkjAEpRtlBAz8m/R7SGpcycnb5PwRa7el9xZMmlrkPbc
40+SX5saue+U37/T/SG2VGyo8aYaJXvhfkJhiqphHw+8HhNn6Cyf6/VG20ZoAkibRlCK0Q3rsjLH
cu8GeDNnUe64PP87lpIup8MjR/AW+h4+yqPsfI07Xa4mjnGsopo/mOGUOTp/U2L5hYb8QuZlHEq9
MmUCXKZQq33t1UGP++V6HQC5zrwt1W6OGvjd7BKJePJ2EZFkNFJpZwj1nf9ViaAQogQZm33uINVA
g40YpfRvK+Bpj5UJ3QZJPX6bRWb7gTessRPB3aoYxVm3rFIQZPCdndNCdas2N/9bR0SbUIYBSoE8
sv6Hj80v1qQKbFQ6+6Hl/zKSX4SebJxgnXdtq/1dfN04VFc7y+Ai2AmnrSyv8LQG6TCRHknkj4Uo
6YQSHSmM9+L/5YGS1s6a82I69omuLC2+OCd5+P1nWhsmfjB9f/1h3coB/qSYvMDtxGqN79hveWAv
7Oh+B0aMzA37dOpqKzq4/3HhgSpULygbstzsSmHEFx82GyhSc/UgUb2JSALj1A6JTJDhkSKX4zNg
i/wL/K1nK13TW6h0Nu5k9E4C22dGICTbgAE3TEsRAYmvA7kWeAvUJmfvLeJ7+hVG3vKmb7ZfCBqj
X7gHHOkC10qQDKmMDlK7xDAV1kvL3XFtSN6xN5PA0RxsbiPyiv9/6/2ieuqgGlH1pJga6QV2ZkG1
1Z3p50whVHemJGHv82TNY45/M6r1xaBv6ql+F03sj2MS0X9AiGWltLtNHbFw4g4W8p9FxkYWAsNf
L7fzibbb4tB6AZEEceI5bNuXFjlB363c9b8Z3NsjIjV5LQoEt9e0onNdgGsMntwdh2K2XJ+Jgymv
6i02gv4UUGpZ2t0UYhyeePicfpFhG0r3DeO7WBwK0M21g4MkXvZrAlvhuCoywKwaTeqhXp2L2ODj
66gKGIphS9aXbQxhzX9jw42bJH3f4Un270Z5t8c/JX86W2Pp6wOuwWE4OAPDFsr9RQjpDZg61sg9
HbwCvHKA4OVsS4IxaZgdW8OofpDVoovbeRkA4QkRbcDLpeRUlMU6d/s+x7Gr77uMlW4wXomL6q+Z
ae6zY5NIzJ7mCLfLqRQRqM2FkFtC09MYpR3JqhFG0ajaBQvbI9jfADNsSsZpFdVCR9GmB2N6UN41
7xV9BrITgvJ7JwJvMXtEVVjiMm3ChMyGfb25s0tKyXCtmWtXbTvAruTB0n0u8k9V2AU7mbEV2XGE
+DuF4bOFdaRWZxa2D7xOfPzPrBK5KSHmWeeIHFMiAUMDjonWbb2tFrr2ilpZgNrCR1iXFCropBam
57/mE5OjyhenD4gJyhBKrnMhpaYGEyjnCXBrFeY4nAm9Ni1k8GOJW7fxbLXlVNHOgiWReetgD8tr
3WO2DY5AGaNRbpcE3F/Ga3i9Pam678wjGRMbrj33o53FEcyZpRdJ/GEszEAT1L72VhrpbYV/gpvd
+K+wxTZCYBFNSKE2WHM6PgUSJ3WTobKCUumYc2Eu1187oaz+/SlhUHEWWhCxMLdTdb8jPPuSVzb9
OaeAD9WmPaKDNZQ5BDcEoVjfurMuVh6QoOn2XdtmB+BwA/uFRPo2dCs0vpR8nWj+9m+DLGTLFUbr
Kfoe6CpzfCcRRx6PcQ1aVCT7xcEESK3cj/ROnj2tzIyGNXST8kJHLeaD94e1pP4WJbzEAKVPRzqy
FfEntduA5mwtJIOX4+kGWqvp2i0sfxKHY+ALdXUyZtHfcb7o0nSMTh9klg4lnhPpR3wOwMDFAoFm
8wUOKKJJXS2wU4Q8MWxw0CM54KmntYbBzZ5049iOZIVbumiojgPiezQJXaT97d0H2tSyurvyhNEc
Zf6le8HMhyW01ufji6mHMVK+iYlGbq5PGM7kC4DgG9A604Qy3ZB7CEOk2PY01XmjCdva/ee4aPJ+
zdYPqmZi5nwnn8A/yvk/xaVy512ySzChvvdAhw9yyL46ijg/OqBmGoVkRQr1tbsPAypFGC2IDMhQ
GZy1ee020ilOYG18YIf6t3KJjoYx4CFs3zytRT9nmPwiTE7YpxiR3K72a0iBUE2drMSe761V7WTI
OrMHYu0vb0Yv9tE0+yztc7BEIUrxODtXi4uRkXaypUynnADrHtRY/qW1sGEhX8a1JUtvhItP0+TT
voHMxeWYVp3A02fDpzHKzwk9ixEr9TQ9TUw3XJYo2fi1c6JuTnNs+KP7/AlQj6nGUg2jzAmS1NY8
5680HWt9rZQLGGFwf2PsdplaIy3cnqKqlgClZ2ZPtEPNKjjmXk0lMDPXO3FjQZU0loJZ8mdFojp8
6Cg+gPoMI4rYFnxnPoHPGBiVUE0uY8hz5AtvcO5Nl3tsOoBMeI6a3U9a51fBXDo9sLj0WC1IyK+S
avY/so8zC8wTyXTf7fX+qSGCIpXV45I0NFqVo3tB1DJFSDb5RIqSnPg+wSfMSMYV2r+FA/3ssAqb
9Sj3NvO3PROntIFU6iJDqN7jAZje89rQKwYu3/BzmM5VBk9uxwjw+MoI5W1fGRnkcYHVN22tu7Hp
CA0FGmip8/SB97gp+y1cgd/1HIgX5V58nSD0knOBiRMD6EBWng2VO+pjMInEB3wsvKZwNsvnWLDI
HVvFXlf6NAJcxfySKT63aZlv5DpAcDpLpkP5P2McVyrVYn0BImTezUXbd48cX3a+tb4xiTqrzVzl
NPSHL541971k/bdnTv3sV0X+6B3qi1eUAB5lVVgC+26CYSXiznIkGI1SDNoKMF9S/N3vcxolBQk7
HAbWQW6R+aBNwgxuLdHA7zDTljY81Sk1ponQF6bqpDoY9Fb3vz/6IW2XjdeStHlZiirrCglwXboF
vN29JcKaSoPepbGEfYnBdzaPaEVvVHYvgMfY4Z4clTJSnjqkg2BIDY0zPYrEbzU03/K8OaMdipPz
zMD15A3TiZnP8fqzIVmqa1dNjd2bqryviRiQftsIWglC6ZjTVtUJDLiauS+FSKcbBLE67fdNivw3
v17NI1q6//q64QcWkhNA1GrLyO/f8xoNdPeUOA0CeVufAPla8kOX54L00ofpjqcXobY+ZpSGZbPL
WLVc/DF+YGNGmShc5WoFqO++bIR49bKWq2XIeRpFNdRK5/BFOoGpdTzwLSOJJQTsHXUiC4AMJDU9
AUPY6B2+8ohaonI5JiqA8ISC9XhrY6Ze7rT5DQEbmJPMb4EhmyIspq8F0aKnLvPWT9UkVTzdt/2Y
r8EAk9bdI3vx8egbhPxkojCgq9NfWada975GkVoJzpIeTiNhP4CNxcLnuf0ccTDQG7VRWfAomURc
u+DIWbGA2WxlAsN/tUPD0Walnmhh93CLuwtl9Gg156jCJlz3+eVvB1k3+RfR4tCpg5LaTQOxjjI0
wb5aisxclFw1E07HIA9zcpJUGijc+OBiSy+A5jwGnLpYECimiHk3b+PeqROHmVpCdY5N/EtZafMM
SZVoXeiddxnhA+544hK+SDT7K//64hMkbZI8THsswTw9ExOzuOxwZNcGI0qJiRhtf4tKvA9CfMnK
OiVTBnpzsy0RuoIFLJYTJszQ6OhFO+9auZKdqtusSVF4noknBlbENa8gK6IBGJVJ3JZth1ltXdM8
Bp65/PrX1u5sghdVpIO0KPhbH+rfguaXoRHZLMjJwomKMYLULs6jb5FY3BvKM7C2S6yI6LkSrPRB
Eb+B3Ghu1IQDe7MIKBUT+hveti0AdvpJbzbCDqGvmGHoDCklz1Jg7owtgJEQH0+lzND+KsucBtEQ
w0VJrSXwhJSvN3cymvJN04dFpagEBvO32K3luY+m60bzEiXnyh3c+71Fp5AvwivGFFl6b0mDGdDW
SykqUM2gHLeZOHyzdc+G1GY6dL3nn24aHnxGtiyKRwbwP/58xu4nIjm3LkOtlv0/5H1gEG1l3eRJ
b35TRxkW1YrVg2r12ysSI2pLqeugadxykdnSZQIDOu/Fag+fzo3rKraq29xBWfWRnPfQYivK8wyt
JblSAIjgGfeTt5Qeoqve6a0w5hYAKWira9NYzfBvzOMi/QONofMcwjVyKOLl6YS+fJaQWpExd35U
NEM5pZNzU3y7X458NwVVYPcsZ5T09YbhFnRh12A/CvTTZ0O5la0+m8thj8PY8ajhSLmNXor7WB22
Xx+oM1jTFkQ1sgrKyNIH9s0zQ6XY/k4TsQJOimQmxSOGTp4nvCkQ+YKbGMt4oXoda2FZWnUjmrmQ
o7d8/Vkz0HD248hsLZ6IDnkDjOF33Qihwf9LIwaamqIDN3KwY4FMx8B+BsVSIYkVw/2LoxkgL74Q
6BkuTBWMrwa8/uZEz5KYzWhtDeeUInIQZOlFqgtoo+haw3gVPg3n8mGucHNz1qtcaTLAeYW/MdK+
1eaBa+VEhnqG+3Sf9Obl9VjEhQAptA4rl8qSnClY7ZFsGHGudzgNvYBfouY541aLIlwAKIAzR6xN
lqOX4Taz22eiZ7vxrDVQAMLDZtDWwoJTciHI3O9YjfA0J/Q2RwfRZ1qU9nSsajVVgVnywa+lqA2b
bEu+baERNUuDurqrR6R5+Y+3kRZP8pNQN2sO0zy2l0aV6lAImN05ONUqNrRh6Ua3QOFtsTP+c4B8
0GftR4g9JeRTa0b7V1pkxdrGRpxjGeg1WZojjD6oC0qj89wbaLi/rEgouCiN9HbLOdZyiISjh/Kl
hZ0MDNIPpfBd/ZUc+/vCJ/P7gAzBrJ4UKAjrCInh8zV15LU0W/YOO/fOkgEao2J0DLAkim49g/Jd
Ce/h8Wq+XYMBVgiqcAoBnrOz28hUq6Xl3KfEDrXaKCmbFcAGaMmrPEbgXuxeU2nSqNE+LedJl455
58e7aPMKUFUDMVQxhkHGnGdu+n+GlpYZk5YOHg53U77LVxnEcKeSYdajtIiOhMN2XDSn5mjFAJlZ
bI3AXQebBTQi9sgnh+Q9LyTJAHmhewvCwNAZWCdelxbKw4kCzEUF2fDPKkgOiA07J1k0deQEbT4S
OGKaDr2W7Ip3+UOeHrpZzoTIDfu85euPBa53NH0UySYkY/t7BgXYGldxp7FwQX3NUjHqqjx9w7Dh
siQG+GIVfRxwyO5+AbPOI0NcNhfVfs/c5QS3qLt13JYzEfXFdsej1trJIFyG3OkFiIXwb0QuALjo
M4zdmEf2U4ZyuEmyDuRACx3P13fUs/1SPV54W+FyVCtj+5z21kokcQbEnyAfRpm5M1KcW6iS+wik
Lmdz3+0hCo2EKPACUJjDANkL9wsuWodZx82IACaeC9SyGdidvfFGvHqjB8Cu00jK6ARSkR0zOyQo
AOZfdwt9bBKpB/I8ZRp7yybyS18We3/psABc6rdXrsuyiSAfDa4Gq9yxY11uJIxKIu4tsDtlp21p
aw1/tturGor9C6Mhg7m8i6T1fEO2E2Jujr3EITJ9s4CYnGSS/m/pL7gCW/Tv0F6rGFOzcKne/Y4e
6+u46V/91aHr28HZHxKeOgHsXuiJhA2WYhltzUIg1qKCHzMVnJmd4UtH5zKeBIwL4RTcKV/uPfHd
CJZoviBOs+GHnb24HBqjXI6xN6he/fLi7eyMRB5Pa1e2kiMy+ZR3U/dMSN+s7w7/3Z2B+YrVrDvm
K0Fbqtrc8bdV/3P1OSuvNj6TpKwa/hHBm+1+jmAbCtTMBbS1AvZhK9A0yvKb51mBwvYfL00cqtxf
A28vlJeMVw0dsL9X6dOmeWlGTyS8xAtpxvNMgH/KYF3+5inXbnVd6cb6y+4Bj5sFQNmchqp+BgHw
4M9y07zojp9BDxe97g7zTYMHdj5G+mZhCvT+tKbOeKoANO3mTb3X3l8AAYFQUM46NhC1qTuSWiz4
3tXlwRYuy5poK2M6RmFgqIvWAi3YtjtX7JaHfPNTQ/Tt8UMIwgB01vk9xRaN0beVl0uoqcbi6C8z
IR3NC5M+MfdLJbdef2vNG874rkzfyW5ar8mzuziglgZVVqhS3YTSnJvp8d0pDZ+E3sIvcTmJ49jA
O2JFL1AFtQjOpRiG/QPnLvLIsdFNxO9TJDJSYD72tCpKl/2vgKXa+ekIUskkLcWBFhxakben3fne
RWRZXPv3c8GhepDP+YhygW+kFB935j/oEV+oOy5qKjul6lJR/2DELOFizVi0BZk8GvSDPK5OsHqe
6rsiFNodEW2Eb0R1Nvd9wCdyw4LiQ57hHtQLLwEvxKeNhyIy+eBXVCnPdOSxM3qoTo1fhR1m9R/a
n/MoMNkPcB8AbuHBQ7WaSBc757btoFMBWPlvnRJ/4YAzP3TAO7sZqrvmMs3JK+5bu8eUYv/L0DmW
1HGGVrZoSbK14QYusVUB5GMASzTrl8ertwI5NqejEgtOS1halUCzQW34cWnvCJRrUDn1qJYL8MOq
IKz4WWbyOhtNQshskRfo8zAxglMpoFJiVXwnetDuYG1DlOT5CN39yHQhsbm+uCdcq6scCNdYLHRX
J9pL+bowjJ9tk3D33czJjCx9OlG8qxhbJJDdjOCFIgPnGhI4v9OuEU9whbIFNaHPaPxMhnJnk25J
0zCYozr24zaCNBdueI0KpNv/jhvEhp4j5Tp7cKp/Sp0fWDDmRxV6elML31iXh3+ZkIBdCJYbkW1i
ic+cZH0aHWZWB7LUdOV8Dm5ymcyKH98aTHyPNEHGvcd7p85sONSBDsy3JoOahRUNefCm8HXYOSGW
IqDRpB9cEBjzJ0Az1lBXYMKhDzdxJoXAWfoY8Wo5ykQ0LcM1Gt3Ya9WlD/BGSo0GXKzsB2QnRxTc
bbqkjXuvL1i/F3V5pssBCQk4j7snGNs+vqTTqcO24XbP2ww+b/Tp+H2ze+9GjwuKq6nDU/euf/z0
ibpY6arK+99CVeCY++t96SQpWq7np1EEgyzpAML6NyftAMElSRRhFwiBoJSJUrfzS9ZdMj/8Kp3/
RBJGK23yDxjmyHZNoD/blSvrsT3l7qAqgzB0Z2HPKT9+dcXKSQKaq87erzZ+C0I75Rku/OWDJhhw
goRtHINYAQWXRJoINOjRQ+JJzo9r2poBcfHCPS1rVDFJAheOmGtiSRrLZdLgQfqcM+GnWv2UDTny
5jVdQ1ufqgPvusfvQlgL7JntW3X04sv0YrUG8mQniRvMS8VzoueqLFeejwRWR3CXxisUsUoUnzTV
O5xCiylxEmOwzuknYMSnaxSUF3LjrLdmywiznR/KqCB5vM8uXXiuNeNyTtFo8ee9TzmjOIG5ixfX
0vjGKZr4sGVNFt6Y8ka/8u+91VOe2QpmZZR7XK0k5peM827TzA66Aioli4YNgjBo3SIjsS4ClxET
WhEZdJDxg4WrET73eDXVt7bd0WKVyTSZwjGLD6m5dQdWZYU9FYrZRYr0HajKfloxHLElh/pfql9e
ysBk1bFScaf/vBswr9ExuOF1k2jpgE+o6r3zSt0cLXWD/tDeN39n7KpgtN6qZp5eNsHGZp4bDDem
9vWbb/KCKrtCdc7PdESVxXOcNMX5ZlvSEZztuFH/R52H6E1AR+VntjDO25YAEftj576k1i3aVI71
+h9Ujw54nw+Lo0UYBpMHt2WFdX8ThEOb3RZ61Y5uJjqkD9ncpjbZG29BbA52LVB8MdDfP3LTtHxW
DxqIu4UfPnXpQcPxcEIBK3j/wPXctps0jB5trAbx++3lPXi/e2KXWKZawNMPVjmTwGNLJNWtfszl
oXWKGOWriy89LSzP98oDN/E7U8ix0Vx44AXZzGZREn+jmjbyA8aSV1UlEMPmtCHz8bbU808FjrUU
VlTzBv696Mq25emCfkUOtSJ4wlLCYF+PsSqtaovWtK/LsoVOU5XAny0Wiot+tI8CF9noPRhBXL00
SSB38eVF9qnQYD7OnMFG2T8vD4nU6Sj+HlmPfj2jUa9bYR/r+tC2yUhDoxSd+Wl47VI9jC7KnkM4
X6FMrCIQ3RcFzda04ZW2wD51YbiyG8B2d0spwUB6qoxfVo10aluG7OExevGtNaZ5awrIRm53Yw5U
2QeuOHJPHFvAhU0uFg8XI4fIlexLrMCAxkAf/bo2vGSXGFU+zPKXBm2QWvujveCwd4rREL643aVV
FaylaDeiOLQOrIe8pzM2nMX2dYuWrpNmcugwRc1CzPiMm6erBORSKyKFfYLiYxGEBTbRsZMbigVe
7lSGqylty8m+rg93a55IJPFMMVqVIteTsFBr2TkpVfpO/F+swk0IJ0ImiXyGvGWvuztpP5XE5C+R
zO9mg9l9JbK81lRXSpREaSPegNqtYkIOmvF4H/rYesjzLcZ5FHEw2a2yIZxtNe54qZCa+AHzwuVF
+fy0jcLzQvhOFgj/RIXA7/WObetbaUCKqUOAP/ThbweVai+Inbve8igOTuEW001e/k5xzo54AWHa
m/Q9x4Lm2oeIoxeABXkXxRBqDTBpKAUdDU+k0Dtld+J0V+OjHjI0puCL5KFFrWBG1DIQNREGx5Gb
FMS80XoFw1WK9l+0o2NKW8jm9Smyp0iug9byj830MHTmbeCepfmpHwNfvNR+Njo3JrxI6ydqlVaL
LYZvlBzT1OIW19tjZxjJAq0z6l9gNUWFP/zgSRaJ6Cb/N/Qv12OgdqLiDb2SVUYmLTK1iFYinYfk
tleOb5LcUHoqsFbsakimoG3hbcakgHtpYWYl+smNH3on2zlu6ZFJqyAvbJ+X0dOn8+lwElaHTXxc
6i+SL5hrQjCZ1D3TAps+L3qbPvo4fnE6ccOI0BExAAgcVHZ8+RH9mon8fjeNi6wzD3vj4MQoVp32
Y+nxv0M2p5Jx9RCFveeGh85NN9Zk5O9uBV+K+LUtceusaFRWgfppgKxACfDCIOHSxrqg2PP7lyS+
TDRlDg/PgkBIPgf78A0NmUSpEtbg4mI5UNbuVv8gtY90TLwxdbcmlUt4n/CCgvmjTh6PjGK9k6kp
hNt2y093wAegt9G7SGSwzrWGt5SDlFvthO830XD11BatP2GiIHHQtNuNcyHUjmJDvEdj+XINhr/h
YmzXZPsN10U7ygpWDdSkasdjxy8uNrOfprvScsctqamFXyBrU2Ybd+hlxTfnTZdH0hSBVinJkuG0
T0Hz/MR6+Ch9/Yuq2U6SmbZHvMlpeIbZ1se3YCz5E8044+6r2TfqWuYck5ngIW+0gCkm4xKAisTu
o7sJkJrETa+RWWuthFqUGmpKlRGZDsmEvqSxflyPFsKUJ5wz7mCN0hSiUs51hoQMCoTWzxr5xDSz
ra7q/viCF3EU4BZfp3ctJ+TJe+E4iVMnapY7U8zEKy3gwrh8dP8ykq4Yw35A1kzKQa67CWMbcUDw
5U0zg/pPcHcLyNLLNcf9bzzVDMCOU7qMhT02t4cAyLO1rs69tbpwfwsT4Iiydr6KwIdV/jodz3sa
MNgq3LbmYmNC8cJQYhEdwdQhce4r8AB3sTCrhDQDqS6ToZCYlEqoIBXZhej8ndsEezz3qffM8ujJ
ik0tKzlBsQ3GLEjqIPqdaBN992LOzjvCj95+5f66XMOUwQuW9aye9ymQrXq5AYbWQcQfq7IMgx8V
9AtLZAHmRS85kHHWMwFMuFpwzhvnEuIiai7LQMlTo94PNBWIiBX6x+mCzlURZjCCEFUP9uRjJVB/
AU3Rg4dcpAyE0y7T/O2g66uqcObnTEJ9p4C5lHMZAJPx12Nmi0kd/Vht5WWhohynPhevPITrjRA8
PsVlEbiYv0J8p6HUiDW4uBuVQSisTo1j1MLcY3rB0FC3p6uwRXViC3Slgj27tUA1zX3RnGbEj5BY
eP6tqv/Ftp3NSm11sPdoi5M/05q50YOj1FoqSmdGAswXC1FcrHoesFSOd8YIpk2Olh8cvMwSdPFZ
I7uuOYBzfvAojbCD9ad9NNQtM6AV5ODH0Fx/SFppvYlhWXaybrjp4uaXo7G8LEo9WhhyOzrI4qN/
gngTTmouYJSnT2Au6CPu54unlpvTykgSlydOZBcfPezqD52CcruYXYMwXYkpc2nN3sy4D6EWSTho
iAw9fKVN3yIC2IWFYYC2LNUHGOItm9y8T3lG9PxBBE/knLvgmlkWB8MsgTa8T1AX6iZvzHlHbJhd
kBKSEMMWfE8EBOav16O5kkY7uFIZlxsgNpn7yzS8lZFeOTKahQ47NLnO9izDs+1W54xoijQT3vfe
aencqQx+QIe50fHS5AZbrj0aUr2iatWP3ujfI43l7MuppwmWOWSDPaU+/B01ROkWj6JG3J0a7lFK
wRF31ho4pUAKuBvQ4YpZxuvx1fDL22HCCRqCYG+Y4pCojw9Er34GI3MsOniHyiF2w7hf4pjTpfqP
xoAcqlmeYRG0NaAGuIgyeBUIngbOjYXzWKvgshrD3KFQlaFj0OQ4iyDQVDchIheJGEIPP26XPLrR
yOlXcVpyuWmkWvZEYFlu1Xeq73l4T8nrE0Ihuo6C3g1Ywh7i42fpF0MVCRKAbXtDHcU0rUwdniOj
5nIM720xi9/XTiHvnx+yPbStHY4eazjNrLAFSAJFgy85mlPKBBeXGrLxdHkQfLfCtQMcV8FxwCz5
Jug12toaEIAVVj2Ra5LnTro/SWolEAJmzAOLc8YEzxdSPUZ4CPRiLqYvMpWoW0LRuyQVcRS8XTAz
OaRcOxDE8vn9cmPXjy0Ivo1P4N5LI1NdC09B7jCf+hQXFHzLcTXzJxsojLoKDZvv6DPkm49XwMWe
kaow8WrkJPMPQSj9lYEYbPx/gHbQxIi7I+Xs2nYx31lYGomHsWx7JlRk+aPej/FXFp2DN74Y7muc
s3H1qw524qMu+LlO4+NzAL2pvnguo7IO/lV/LvUl2yPcSeQCqmSGKA+jbGdZhiEVGL0yn8hbpUGv
K6fqhIDFCKAUOod35mPjfZp3Ouo9GSJTdLN35qS+xPOJtQ1coBRertbqJCztdT/fHgklP7Npz+fo
MgbJ/LJSkTilD2DWoAWbulYNJbH/AOIDT+jV/vo/VCCh2rzVTeQRfXX/+87N+D9kZO9Ytb7b1Vjh
KkoOKfNTCLk80UxVwASi961juUp0faEIH299jWJQtPXL5rqlxyUPG6YcmJqYidxRoC8SBD+jwOvX
Rmhqu7ZoWU5QSAgSwTCV9VAaK1BCjFA7b8pySADWpQTL1cRfzbWcrXq+hX5HADaBkIx+zOtFP9IB
8DN7tH/q0t2ct4xpREI47ejca2K4V8NyAIYZOrMnCs6mLw0kzW4gmsocm/lQmrIMeq3t2j/Njfva
kCBAyP0aRStVCliXAA/b3Wceq+KfGzEjwJWV68tgEOQFtg64a0R6xSXuXQk8cvhmvakfHg3gt8cp
zC1bC8jkAoATMiLcip8HftFJyHwPC3tXGLngJRKBpXkpg2FQnw2VBIpb1Jg+Zsg9wISDjdyAScMw
vcF7xVkPmI0JQiFImS/KhmZNWEqUwi4FNJmqqIvvDS+cidJeW67L5qlTIAEC6z0pJeTZcqhtvr5k
MbYgmXoOd4l5YzEKZZkusk8gS8A7RHsXee9PAaFiygmM29+EuN+XbLrvGvzztpdXzMve0Y7rhI7i
CCxHAiR3QNCGIFcYy6U3263TosZX8TS+nBD6lIUp5hu9PXgU0hVHUJ5aaXXumh/4wK3V5fzE7WKY
1D/hOlZn9c2ZnXuCQfjJbv7NBeZUpa6lK+fmW6kazNR6LcDy3tEGILqJHpMf4h5+o03Re1oz5PgA
k/yIPzBSyD34w+1wX4gAVshXZbEv3bTS+wh48WWmrwYuVavj11oV3FUueuqBZ/KOz5PDZavYgoS6
tf/+DT+IPirSVuu9t1yQ5FUC8Sy1faxNtgxKDDgKo0xNSnA/IaWEp06LoOpDtfdtfi3URctiqFjz
cQ8Rc0S2o7/4tXK3IknzcmM8sF/TxVFytyxCKjE3UfA/Xj+NN1E8SPwKAvrdLnht8WpKBav9K89u
NpQTGei4fVSnYUliNIV5Cys+jWw5xBf8Ezdk1qAtE697xlxgVa6yHbdjchU8XNlGZNirjvb3JUtf
vlxR2c0x3ZscBHO/6cKClhFNGBmLHOb8GgAPPGkgguD8ElaQzRegpeXR8LgqimM3BdD9gcdxRS7a
+c0+JvbKApeH1o/nXgt055baAY2vxRVO89g+OiKyAWHwbVVYITbPF/aorOgMjDDa2bf1dFN2PQ2M
m/TI3sFQ+c9NT8HeRhTHn8xBTAthpMg+iFTgcNkmeXrFlJ3d+ALea3u2fxPusRuz4RtVxOylmF97
AU1KgdU/1Pi0eDhLVz8ys0q5bUSeJp0TLYbbk+xmQ5GlgPAfzVKe3rFjIV90A+HCiJCTIdb9V4+q
FBBDmffJ3Hn5ziDTE2tsiX1XkBHTcv0/DVnOiuxogigAh7GwnYlZQ4k/NVLh2CQu2ruOYXwnQJA+
AmKif90pQQzguRpaErhq1ecNE9JFfWKUUTcNLDX8CbP7uvdcEzCqzwjUg3FJhU5NK25j2RG1TEpX
PTOA+Nnexe5ws+WCIF80RXl5U0Th3vpUxB5W9EAQYJ+5nYq/yLzjFodEume/yduM9ykadZTk8Tey
ruXsNoz104U2OqmblPbvgpjfGctUZvai5rpz5qXukZmfVmMUkOrRYus51PecRReNh4NCA1dclKKF
Z+OhovBN6FhkHOuhY2KCe1UODRC3Ro0dFEvpe2KCWtlTeRedUZ2x2sr9z9jbh6xoclKPo+DzyuuT
JEoIw5xk1kKt796RcjzHMmV9s3mWDRlpgDj/sm8vAliLri049Yy5dLPWCHVGsyexM8cw15hlP4g7
B3Rkkb+qV80rDyjhu7w2r3PsUMhuN0ZM1pjt6hVrOy/Cy4IHqAFJR9HGWfmV/ULgRRP5RAWPUB8E
c8pM5Qr/hBPwFK1Pg0i5VFCaemBrwOApqvlaJQQRDqvfdW+j/wIIjgorBqDI20Kzvq+Jf3KmDNQX
2fALe2vyGzBXsHLCM2760/Zlqg+jHqIQb630FHmjwU+uWr+gkXbABGjwFE1OtzrlapjUOgdNp//9
bM4/BICZ7PWaJfLMFYsFWVGnIuhxmdkg3n5/nhao4FJmSyVYbv7ZXCaFOYiSCs6Vl/bZGhnTz3QN
Jk6LjepPMuTOb2A+AxBQphefY+d1hnivKnsvt1lBcvxZyIlwalZmXqeb/WWlZMDqvS+J3ZyHJKe9
Pofld1o9a937bjz/tIycwt1ttsqIjH9Sd2dqcnfAsKYeXQ2IZ683iwMymaDVWOzfo1xhOAlnqebR
qJAIxmZYK06fTExOpVdv3n6V3QAGT89Ni4sIkRVi/BlTKyjDpPP+nBCFyTOdq2poltgurSfuoUmM
pcR2As4PSYyZb5i7v0L2oJtAyxy5JTFJpXicK1uTVcCHDVmEOF7x9P7fhHWGllVu6krhswLbwTo7
NL1Maqd/EXGflwElstnnDSu7e368yeqVMugOeeG7FTe7ahJx0Bq1BNO/XfH+I9Agj8UApKQppWxi
0wMfgbPq1tl85gWDxFbB8HcHW9WHijZ2OlojACIDnOLEnMivltIbHf6W8TkBgXxZ/STZepjUOvIW
1QfBsKY2kQ3kNCJbPMHztF9chxJvYIBZUT7s/m0r72GumyyXNLJxuwHBz5Dw8ES/PncUBB0POGAA
vxsWuKgf87tREBXPkGJ+77NJaNG0b3P2uifrRIqxZ49cVOyNhHawE6xjjrjHVmsQ+5SjrTkiKkq7
ndw1C4jrBsFXY2oIbmQxAzD6vklTKdblPYYA1Ux/EnumqfzrAB6ws/0V3hbzVSJJwq79doqYoVaT
+JvtypgEBdeP1xGj/7xLwDb9wds9TsMqtMVj91gjSwkEDGK8JRsAGWVsAiJX4M22RWFUshVlglRB
L3YVvxbxSWMpue+BbZGM7njEJ5tJzG/5FPtlSf6B/okZYLRIaPEf49szjkB3T2PWC/HGz9MXHFjN
fph44p0+c7i1S2xxoPmHGKrRTzKKanSAO06OdHo+jPPK7Pol05uvC7E6QgOvwR3eSVH2shLM9c0q
UaQCwWZ5CD0/dz7q+qY0J1wYvKKdoPAfp+gnx/tWzsjWLAm7jmcA+mHKYYkiYbxPcqWGkNk7CM+I
CCMgboK3CXTBcJz8XVASicxf7KuYIPndHI9Yw610D0V+1Q6Jn390aVKBvBQ1p8GGurNFcHCslMuV
RO9qSolRPy5kSsVRxe7OsCiPnVVl2jVndRE+iHDLwHLjaGoM68MPs4fqq/1dsEjnXws8WWhENEQN
JqM6AjB24lzklXt9AS+uirRMpAcOXMbD13Te7zF5N5zXCGlbaJ9T3V2hO9WszRkybhlvimX5/geJ
d6CoMnkI3j+MpAXPLcrxPt3D9Y9xMr6shJJDscKI5XgC9R3vwzYIaFbrAwNDPmaYBiXasw02s0S6
uW8b3b3E0z1XXAe/tkmoWVSW6P1GpKGwDwYVbEgVCvN70Y+XODql+H6+yaHw1cXtCeqjDjHsWAhL
zndXIlX3WfIRxmRwZDrM9OfLlHyEEY7ohqY/tSuR5Lonj9qyHVJBYo2m1SAVZehDG+idR9VEZ2M8
ugj807QgCmQcZ/z5LwtEwlr8SLgvIsx8AlB0+6my5QHEv3Ub+SU869bHLtNp78Rx5QfDPDIEF8QL
PQSVw9CIFEHDjiaVMs7W5Q+vvbDDoNdcko8xf9nkSSoGz9ufhqLPkz5zImHuX1jWO+wRk5ecE0yh
nkoa0zJLEAsvz+Zexfk57a4G8suW6a+8bhId3hWg8MKdOCqrj5wq2XyUQKhxog2cqOv0w4mLWFz+
iBp9PaM9mFvHsbu8ocJzcx9LdRa6mHPqPPkHJ9C7H4n6YhInFpQiFGsOF+IpqXtftntKBoGfXV9N
vFvsC/hJmgzmARM0VVAHyjUFApTvLIHBV6iMUjGUF4+jdpgi+uPiryJZB8WHSWaoAtugz8mwxScz
lH6B33LFcxqsmVJiJ9TD0jdR+rbo+rtf/hwt2wuJXIVOR5XM+NdbkbTiXllu9X1Kas7oYuyWeMNq
HT1+0EQHaw9HV6jwFFVgT2R1iqS+nGSq/grgj6v8Mw8E82yMkQIHVGDFh+FxO2KVWBiP+KieEd4m
8Z/FhYRWjUzGbmYUyySBkkFd2XUQ572aHLprJpzzbvZdlh5yfnN+sGgitsKNdRlAnvP4mH8Wbx/9
AmQSEitsTD35ZPV/krMtH2q7uzYTA4VQc6N/Ge9rhtqCFQgnoNm73q72Rm8FHIXGl5HbvVO9Hann
igfzLR9RGc67wON9CwKGx04qO8bEkn9njriFgNcEN84pswN45zstoauY/ZdFAAjCbE4MeihWo1nY
o/XvYozFcJ8tf40zvGnG4YwLWCixk0UOD2mTP9ivrmuH3z6iXZyeVFL2PCznvhJRTAPMFsc9qpF/
5+8Fq2Qetl2HxdqTr+d4DAxu4sO2yiuBc0arTaSIg7Ah66FooZ0wQgOGduj+FC8PgWInk164M4Pg
5ItxQOl2+Toqojh5JaTLu4V/jq/oAOhdsYO3EU58sNFf+JDBP6rEaoq3o56iya+VaYeZW029p1J4
+VcTZeBpASbkdU/or5RKQEVPslfJHBOgCAq65PVCSsUzMlcadlQ75yWdTY62pJGGXIU322OOX43a
IgR1XYJQ90L7CsNAI1L4znzbWlCdbXGqXpmKqJbv7qc8V/SrGlgg17WOhLxYqJpJgYW1Ph1Ro9sA
5ogkacnKSa0Di7TGXCFEFmpa1RB4R2W/WFcjXF5AlD2+7dgvDnez8WEgEX26e68niBeZd26Ne53t
CaId/c0akLsGIW4Lx35IwzV9KWOqO2sBdNWGyQ0KdbLixyKd6Sb8lyrFfyXFpVAl3PB8/YL2ZFGN
TGE31DUR8QRHvDcmRAmeUtqgdenaac+nGXQ7yM5nVYDvHUlYyNDSYKQYXZXu54pELFYXlztn/se8
F06HVIJzBIQyaGTft6sfUZJUSqfp50NZdr1TV5/beVJGhLZWjDWQppw+Ea+uI9krGUqgMTCS3yT2
Le/UH+oMykz44UP8nQim1rQvEPBWdWG1m1IxcAz0qVpgPTgJLbCPLCWTdsH4YEL8VdRwy1uw1GUY
+sfTyBiO2MclND1oFLdk7pv+U6wpXP+MjNb+g3p/Fm9WcbiHiMn6m62Y4lMZ/CW9UpM8DoYeu/An
7M1ZB+VEBEodcXlMe+/DE8yOxw8KGAO8SfDrM2VwZtDQ+g7W/bllg6Zj8LJ29nvj3PJJQGUv9ji/
jTSHXKy3QPdYt/lx6belxIcvke+O35Q2E3EBQVJPTv2LQHFF5XhyqdW3lvpQSUUXBtg0DjWS0kwA
0xLS8ROS6nH6NE0YiW/a/aS4Dnm/1FSgZaqLwBvcqORntJMeob7aRVBcFsLUbjlDyunNd2oMo8hH
nJo3RPV7RBDIFPOIPTiD0MiUQwpeYacJFpcP/jFPQOFt73mPi+Ly4iv9sADMwIz6pVNmc/pMqr3i
kFDYfyIDrVZHueJtFpl0oC8cMNcd8uCumb4Z/89IQANHD3mY0wb2n+aKjI4u2RiE4CyNE54fIX5z
GoGoLY7Lied6x3MpRJmh92meFQqsJ35WCAuApSpyHlSDDc67T69pLPH+STkC9busx9ufbTCQlHjP
c0Eq51C3GPT6LtHMk9rBS8ztEZM0uerzEzZ9/DjrhmqzChGv9THoB4025TGOJRwgHm1T3fnhQK35
YZJK/if7bpYrWmEqO6/qFL3ke8RZUSY21ZIFOuIO5BxobqynyFg6YtTBgCPWzN3zF/bYlgZ6WvPQ
xheogYdxtIdQNTHqR12WTsrN8Dl4dgNTRvzzE8/VmCnB7soh8te0th2RLC9ubL5ve//ac54Ggy11
u5IBEfyZk0hOiM6TBAl7YSM3tLXQ11QaZVgpG+JOdhQgrzMD1rle2Hlx/P49zR21W+aVGR5uK5Zn
92sAjMCTN/R06POPkCTCbuDfW1Fhp84V59k9XJnSu5eRDY0YeiuJv9uVk22/gZVxT0hXGcyrq5yf
D/KmWYtqcfPiQm6jqw8SLW6B4lLHRy1ssshGWlUzOEFXf5gvy94f2Lvj/2RZybBsL7wwXL3Gykwo
Ilpo1IS4HjcH2s0d3DJA9wGKukN3BXvvpMN+sxhGWzUoGZoY5b/EcZTQ0NBFzfmi+4uwEDej83qH
9XSiJfLPxlpOlg6q5fy1S0FJl1tkcsA3HBF6b86qtYNTmKCB3M0ZBlRyZUGm6I+vGslitSTq8lbW
lY/PtdGSBPUpCQ+4ioaVSHk35WKr7LK5+KgTghUvXUBu8dHvCxyvnLQhFTmIDLbfXImwHdl9V65r
Segno5+JWh71CUzyD/s9hX069wjouapo4YjZQRo11klPL29NtGkfOSKcHfZz1EYUOkhQuR5h4jbo
D493Lp/FQfdEZkiN/iWgNxGpY3KidDncytzY0MjsUknIDK+BqPiwA7/sxazVcnoKuDHGH1kDBySf
9NH29JkREs5jxYUzh6OsNN2rtrBt61iPgFVMI/yb3QVRZYri1+FiKCBfx30tE7OAXQa9p1lun7lS
qG1EHD+DspgZ8sXzJIzbTwYSXGDk8kyJ9yFcK4KmTZ5XRk01vlg+Mu6iLXO9rVLx+39XOB8z75gI
WXRQl9uUbIljdFK4/ygmg1Ylg08LE7vVSv1+5tZSV5tak0FSz3ZO+gPzCX0oBdlhvl7prILUJNUm
W+1Ak6Ue/g0rSiq50zXcZKFddiPrc6wuFARejlJY5rAg4svF6KXOqTv2N9Sb02Y5sElDgTSH1lBN
/+eDFLaT9lwZkyZWNu0e3stNv+z70eaDgcD8DTFVsAu12lxSEjV5BnZNXVHVbmKE4UQ2StyYmOR7
9d9YNwHZ70daj3Vz1UZqNRhcZgGilRxtBcDOU9cAiZjsL9bJbD5BUdXBP0/0/5WmTXv9p3YhhKDQ
9FBTpDDp7LQUANEAnCv/5yMuBonmIm2DNUg18IHIEZw/CImH7wXbr4i8JdgiWseaJ6TzG6ubcKP/
N7ik63Kld8B82qO1aBIszNE4CivVYB/0HS0+gGPou2Fkpklnjr7iQaQdNgq/kI0L26QmN2WakLVf
NEV/1pxIXdQztKyKX+RN5wo3f8r09vHQF7zKfX8O5/bkUY9wO6Xft02ThTLsydocEy5Ly+LUf+eh
w1IUYzgzpIbsIsz9MLjjNbfFbNxC9kXflg6gqRe+FSqGeLUKo3uGg4hzq3C1FbKe6vzkyR4miB6l
8I914SO5MERakLXjp41K0Lm57DK0J6c+3sruAb8GbHqMgAMOVOPkIAzltr+k6Y8acmjbGhbyFRfB
ox15pPR0CwW1MlJLS6HD4n3CcQEcgqyWXnFyg09GQZAQoWxhvQDy8U5TzsV9c/kg2+HjpJkK18a3
9/rtuvAv7eminVqsIecEOS4kV1h36bnvKoSFokZHHxKPZJzKOerlVSt5Qf3queDTX+XZ7AMNMI+N
CP0rROkbbQL0YxtRvm8o6mGewYuXg5AGbesHT9X4ysW0r3H5pkKOvzObscHnRJ89GwYXMHzEfS/a
RWDSkJxYggTK3GK95ybz/dbWL5UQMpL97ZcaHTnXQvOXCrI0Gv8Ho8igjvnP/aobCCcgJInJUEaG
ZxP9C42vSooPaSlCg10VpieNCWzVG2edf4lXvTvaUkeAxEWrbhzmNxjAndxi4K7jy6XgVxge5mCy
czE7kmEzKXjbTwfLB1K/D4K72fOTeI4s7oSZQNADHtiIdHhXJg9+az3v8Ctgf7K4pHt955e6MUL6
YrgApGfmuBKWpaj53QKyAP/kiHbBsF8WIq1GaYHVwUK54TxmyprJyxp9sTaA1SnCfJJhISdIAI3/
eZiQyHUL2IEQhqybnS7fA+Xeo6vbrqAZzrYXN8i4EE5DJhiXkQdqN67nY6wN19yHmG5fwbKQI6Ru
O+qekhzhjDajVHFQmAnAC/X4kMtQ8uqAueQ1TMdF8kejLWuZbXEis8ADHt31PKRSMCc1xNGqPWS5
NqWApQwF1zlVtWV1ZTxISB8jX44mrX64XKJjpe5i2Xs6VOehkiSmXOtkhBFBDi+dIEQXFd6wgQtp
JEpz2Q3Mx1kA3umYmhaZQOlTKZm5G4e6z1OTtut1/Ji3lZvY5VcFVeO6J2n/CwxRQY/Nb3qNk2Ml
1tHdVUwNMq9c+qSywL1osSAkm+U62i5YXbxvN7+wQ4gZAavloAh+1I0eVxU6ST0vi1byVU/uPkPf
iwT3+dKcyZZq6KEM6N6SGMrbkUFF8NhWWASc43DlKOH+ZaIymtKa6ceswYO0eDKe7BjJrXdHX59x
ykEJrhnJSXIuMxWVRreRrWLmlv/deYHXw4YZ3h1U+PTSfZxeRKYJdL+DCJri6labC8K6Y+CfIZe2
4mzhfTFIY0WMLreGESdvKsTNz4Nj83bE19eYGJaAVQ3nwsLBhkgv9mcyvrDFvqcqBJfpUxtEN7QE
pbKkFN2fhg4x8F5tYdtSveryDn1Xn0F60JMyMFNclTtEJKQTGPStRuO7Cs5MO/gLIBrXcQMcHTs3
x2UocpoDUIp2KNQzoq6vgnzVW6ZevJ+Oe+v9O5hBhlqOlZU+Z/0dlhFbH0Uq47H2xxfV7tAFK8Zh
VHBp/5axk4mWv+lzl9xZXTCI9IMJ8jtL/e4Lgl7Q++dC7T4eqT96pcoAwBe/OAzNI0kk7ZnypR22
+8qw62j0icuDYysMYBeM3tZjR7jWj7BtLBOsaGQHKOgJMLle+4euq/Fq5Y8ZdQKDawyI2GtuJIUK
DrC/ZYzNqX+4bJoNd2RLMHX5FhXRMvEKVLoUDUzSW3cZe8IDYb7UUkwzcHH1Ec4BgMfHWPbh/UKK
tJZNgW7sdK//C08hFpLS+3Fq21BcpgQN5MaOOq5Xz6Te6pRW0kEyjRz5ZJjieNvBcq4Y5VrzY4kl
aA+yHlYsQ+C3dmtROPh59CkAZwfydKzQIXBh3cJ8xoYoFy9K9mBe7TYX6o2cUXbsFnZIn3QAWHy5
HQDGmdwbbCAwOlBIoCdMsGtRwT1H5236m6flZoIBQMV2DIAYH9FbBM+rcpG5wuRyIg3Hn/7tXji6
rsWDrN2rVx+mOymhGgJeyCtMxoC/Q8sDCJcwh4k9b9Aa+uZ7xKZ/yvZheVzu39/FfIIU1U8PCJyX
myg8tPZhpfVupFPjfsYqhQTSaYAICvAwJ1L46cpNYX4X2P+Jln7DDXgTVgqJBvb6io2VoluALzyy
+ZgURT8/vbpJmrJkLCDeM8wVLUrN0J1oq9rEmA3w6+P6bojdz2W2T64jWYniVDcUZDa3+kf+QwvX
414+rQ+yF24USB26c8OnpNBdKqZpRiWYGREXeYrejX0yAK/2AfeD09hRdk9CJUoFxfedQ7wI5whQ
UtX2/IE2x3jEQrdh8PRm+fv8YKATAoO6tS+MZlYqulHoSswrH0wvn1Ei0spU1RRZ4oYXW+nDRkAh
VQnk8xuUO7dSlkHqFPzBXe+l8XkuHr0+TgLO5jOr/5HiXgmGWdJehL8EYvEb1BTi5BkufsGtK0Ep
mmvMVWlqeE1+L4rW7X0Ywb6Qjj4gIvahzIFvJfBVN9diNfhi0bq4lGfbIWu0Zs4HXdW/I5Z803pB
9YOrytprjgjdj0D3US8sdqRGGZ/idKWpWuLybcPvhnh/TQUK23TyDD89eiuRzDm3JKjfUs4YqUUH
/O2V8KOJ5BxGN6lNUAPk1Lk2oh1gFeNWc9oIeqkPSvdM6thdHr4ErTXCiKTUyBC41Qx/DV1USmsM
iIIe2jxyoHiUaoyz7iHEWpzknCysJ/smC4eV9i5fiyFuhGJH5dPOfEb5BKx9DY3ZJrEMwZSxdHxH
3AXL3i7TEbwM+2mP7u/wrqMkfF72kuqpPxdagLEVNCBZ3KnUKfpSuOpuXlqNDLI5/q0v7U3Cy9XZ
vRA/YZ7Sh+5uFMgR9vDZH0mJ7FGm6vinuwUnKnKRApEHaVW1HOTnvoTyIkn+uYqDmg+diVHgZJU5
vnfniSrZ4JvkznbWDCiyjsXNfkAxDTMKqx3vDwsYInhdAm3Pm0m76oao64zdDFPAuNk77FokVOiS
Hl2njoiQrFkm3j/709mY0egEI+WPXS2JqVG2EC5LSGAVeViyO6Ly3K8v9NhMcnjW4JE5mHlgcq7J
SZX0k2k40iiWaTfcMhLd1l/2XwMlqXg7XQ9XrQTZ66Mw3fWpJyvH426YBf8l/vqlkI7KKCoEb2XH
1Thz/xU03BCLGHnr7a1LdGdyNzphYmrNLUkvOS5ztQrtbpep6wkRECuJZJ/UPjedfRDb+DFkMpqd
vZ6rFBFUjK5qcSFO32VbhRl5CG7LNh1bhOjLevtoCdL3dq/cO708L9cNl859ABOvZU8REoWVB3ms
F5tSXyDR1rU8wLpLdkht0bXmP8HU2O7Tj0UgTEPAb3/FLGtyBinkuy9TWcl6caLXdARJkh7jK/GB
FYCIYM68TKwBZlYwbSLutbOuAPBcg6jVwgtZnUh2NvsU3BE+9+FIhGp7R9A6+yXZRt1m8hrVFkkY
j5bBIsPGL+OQETBIQvj6YAmGk6LTdgRbnJNkoAKC/hInU8gMppFqSSR4oucED2lw9dC7NxfjmZJ4
yx9yUIHMgJl9p+AjpiFk+Edc08DzUzl9z3B5X4dqYy1IjGuan9MLFRX5ylArlDOOHM1VfJ2wZ2ij
9MOxPnl0PAXSa4TNTyo2TrpL4CUbPDJRxbYQavLIetG+wR6H2RlGBHEp7qCqMIHm6eRdXg1J3VRE
i6iLXNhNDp0vvhPOAkyup+585eOs3SlFLD8k/ncF0zqOJbslyKN0N8n28aFJliUpMLcDrcksyXT3
r2hlNa+3HLd/9Vm6ei4wIVVjRPgNRch/pwtWZAFOCVF97UvpUIISYS9DFo9rr309Irz6ooWZA+ef
/rG03lhlhkolqm81v5L/jTXlkVz6RB0+wyk9jaVGOSJTvXdCZkl7+kpAb14OWTFdbbMzT7XB00Hk
7da0Rrdaz9iW7s+Y7I7x3BI6Bk3L/1CfZAsr0/JPqoPpf0mk/kdPAZsOFUyXp0PI63nY/ewoX/y+
dvmzi3GY3dmNopilFylo2/+iV6Ir43D6IP2FxgAIT3to6DOo3VO/EpGPqu8f4056uOWEltws55nt
kfTLrvWUX55Z91uGCaPtpGoCPac6VsE0TSJf9YI384MkKtW1wsp+aig/ID58fWvpS+6nQnxB6u7b
8tid5S0Gud3lRnmpwRIvT9otVjc5pmv1X3+a9t+vcvdOJ2eOS1wpApotMl0jmXsvZy7txRZS4B8T
38lYGsmykKuqMJgJTcAQnPZhQ1ZFB26n8wtD8yC3rkAZkYjmDJnhD69K5PnEq3u2p0zLY/QoTCy3
z/EoIuIpJEiGfKjUltEyXpMjSDjVdXsZfMijhgrhnEyTEAPLHaBr4znCg+S6s2m52FRBcgMSibmT
bNg6lTUa80iPpEDfXbHSrZ39QoyyqaFfELpIL871iHdTx2ievwnnoR/KD89qsLIp/eZQLghssXpt
dnWsuE4Hl+Yo0RXQ/5AliZ22Q6sJQTSAV1AvQFUZ/DcQeukeM4QZLvKozzhNwHJU7iiS9iWDBYz0
L4AFF/oId+1rYEQlMpUlrHuwW1ymiOpLbhYiCcpN7eP7bMvp53/fIGVovCXsmozH+YIGv9iuOEyN
T6d6t3uQQf866htySEb5hdcgVS3nslUPU+ApiLZIQjq58fHrR7mBJYScWDTEGyRM4STQN7OGGPoa
nJcCdNhIZ6YkfBVjbsv/DarnsjCkL2J5oehrmzGlAXqUH+HH215WzDCJIf3WBepw7CEQjru5bz8E
ovJgAOH5M6DZlews2tQYJpbhYuRXB7kdwYuP8BUkyMTE8jGNz7tacjeLqBwI/7fBXu0L9xG9doyH
BQjS9/Nf8FZQ+ULvNSpYPNdztGklQz1rVniuZh999WkdKuQsXtnI6kaeKFwArXNKIKY/Vvy4nsSw
g1Fd5+lnaVq6UQoZcTzT9lvEh7jb9qjhKVrUX8rCPX6fUlV4+TMjqESeiE56TD12kjnslAk00/Qv
q2oyXJj4NZPO4dNc6lm+9uptzlG9j+M30dHDoMnPmzDtHvn2Y9uRUGUVryrUX6cO79jFcbYeMlHu
eEjazxxiQEg/PuiswVLIr3XJYFPSux/8Xw4sj0N8eih5c+zsITtcledxfOBntytJ5rwjmYKurQvA
1C3MBZDGLzJiao9TOuRr60s6s0+0EMcLhNbmzIGpThcNXazhO3ZjDY8NzNTSU1ThIhUfBcE/CG3D
ceSR7ER+b3z8LtxLjRqqzvDAlYcKJaw6fI/TOy0/CmQyC3AmCOvtkrRezKpQErsAdMpSf6YK3UAL
qLw2OhbussgBOSdGbHx9MyjaHj5m++r3pHWUEAj8TnLUI0WjyEBiCLohLKj5msaLAGW+fmnZnHNp
2FruFOhzhkcgHYYUxk6uuPg9TL2xWTJBXi8UnzG9t8T9IiFkECGMyrufmiMQpyyqoOCNPTj6HaUJ
9CKRKZ7fX2Cw/G6wai35siQl2wdQJLl3JNVPm9tezlycXhoBhCyn6wPcLUvoHvXHpfg5KDlkQCSJ
Mz5I8C41jy9uO/1KE/SiN5VwcEr96+PrU0i0fdSaOVVyXykD9CyoGCIwjZn1f68ojjsfFOBc36Dr
o5tjbO4N38yY/WFX0XJIpgJxqpNBzWy/3EJVYv94Gmrp8zJjA/sLvDCMNhZkT4dDtS33yVSKdsxN
RPekp5YcmSwIUf4yhw1YLKV9b9NygpaROJNwhl8mMFeRhoKkMb4YQ+i2I5Hto0yYwEmZMD5aw4M9
mhTkpW52FTsH0FfIK83BMURbNNY9MrjmPa7gFXn4SQ66ZzH4uEILNAV8yX3qcgqom05FRhirhCYf
jgmBEGOaUMlXx1J5c2zjYI1r0fVnJZXGYLzNiF1BRw7yEJLImX9PeqFJXhpv6BTqSAT2gNG+foag
ldxFpcwALBXvFOj7TLWZlAIOaet4BI/X6mE9LNhIZdu82ufngPfSsecNEgjwBsYSrcg+e+KfDg9o
802aUGxQDKwxvESbQcmmeKXOTnaA3riE9NXszxx9ggBcHl1+8Uia/580Ae1vUjLkaAPAV25rQNtr
R/aRBIdnbfwOStPjJBXfhzyQwIIE8/bOmziaC2KAIATQdDdgmrJEshFBJLDs+Ht8KSdebPPqeyTY
sxrlJM1Y4aPp6zIKMvpDvV5r2JFe2Ujy+CJ3sYeUo4JUAPNoqGI7AiqliFRRZXj69twL29MJgFUE
f5rnruEVqB9zgNpFOlPzendqJiKiBprmWdADb80U5YRtSFCH6JCqdVEDQM3ugzPAk1MwQlZapHt8
W91rASFPItEXAr8qIFiCcqoQ96VmLJClm2Th+o/R2ul33xxeYI4HnJZEvq0PdJThh2TMJ9Mpvfwn
M4ckV4PzYZvfs4+fk3sX4EICXqVQG3nmAJiEzVLmKuDb0L0w6Z9mY4BHyBEaQXi9Hor2QGl/cNaj
US5S1ZxAM/tU5j6rN7YBsRA/JBZo9vIfMBK/Q6DZiBpaRBFo0mnbSmqAqwjjecsef9xXvIANwDeT
gIiArIfO9HC6xSt5LyidQAX8/fQC+E5P+TsAvVKTeRaqnZl/RZ9TRESsaaegzAKxbFDGjVM0Yj+s
F7FTOAbwDQqMKX1rOdyj7Ohc/ukZ4wNUe/0VR2EtsmWqlA55iaYLdhAaZxg+2+Jm865iUz0d+k+G
uLGsZ6XsVaPlxdcI+jCycn0bDPZNHyumgBIhmX2L45DuDyZF+YJSuq3fYxeC9vw5N5Rwor7jRxOA
S/Z+HXeCfp4bUHYNWhrX44BU/6onpg5GuxW0KzFNV9gElwwz4HplBfe+UcX4IW7AvAGrZNtt9rAr
U1v9fJUa6mujM8FlMuwPWFx2/gIwyevulq3ZiKUoqm4J3o8JGl9kMAeaBHSgT8vDQzHtK8OJ9bXi
O4vRUvSM2IAxdW5EUiW15cPpPle6mqbSlteYYr/9uOuTeG/DDjLEp9z/YHppOAxPw84ynE67Fjvb
TO6Iwa2FbsKfe/zTZYYUFon3ucD0QnsNBk5Lb1zsaQ8xWuAs9pN6LEnvOgO8wtOWtKHcpKou57KX
pPAUUezuotgsBUdMr5Hw9qfWhej3BBxOvfltsFnKv1Y82Lcpf7FX7wNR4m70jXVxfWCNlomCH4/W
WKJzcD+IHLaS4vN/KNm3SYsohuWDH4iGpuKdP1AlzLmEjVj7tvs4IZwyij1W+oSyz4z/hUBju00o
NwOeFx3M6tDi3/ztqbVw0dATJWKFs4Zsc4sL9VXE5UgfNfbctJeD9XhMVgU8r12Wz/nn15VOUPi/
5uOYTTYd+qyVh3hzzv3iVt5xwAE7+J8Cpr0mMtyr5I2BZS7xXOOoV/6oYoNX5fCEzaSsZM8xxDp5
tbYVS3SeAcdpRHgJu0RODklfAexGquOM9GgjuhcQiwl9ae41LKu+WtAuQmRO6Cp6aKFWJJsJt1Zl
08kM7Kg3XfVlKgO8W216Jrdg19KNUeuoGqa9O91dEx9S1AJyvWWyFTz/91JoLf8jqdGDF1lQ7P2w
C/fOoJrd4FUxXefqmQ2mxzm9GCbok/XUtVsAEcP95N8EXwBBOVuj53mTdDDSH88yKt1yvvuhZZK2
L1Y6K+qpJKX4gchOsdvaLPjxvwSJn1TNJIO76rjWb5i8jHyPJiNyVNY+ASupfy2qNFC3ZWPkDOho
CEShZOGi04kuDjO0WkzN+TP8DU83uOoH4z8tdW3mJImEbquPyzxYjRQTAT1tv9FWxcFqpmhzI78i
94SViUqhdqBZCTkWqhmibhdXtXEUPcWFLWsFXpM3oWto3cci4Nr5Jtq2NQRcz2nOFa8u1pCaW8/H
mvqU9t8ypPBbiPLITvXyCNncl2gxVOOQ9VOFqipHmvWLEEYF0MbD8BFl+6Ckq/0Z04HzeE5XmeQo
EMfwgwLsx8LY57v9QejkkGkAhYlXggyYFpeh3M0CiHwBH9KbZMmaawu94Ns0dYi3c+LCTSaRCFzF
ON/b0JocRDB+78Sq9pAeD0ZkR0xxyKVVz8pp/HE8uYgJszXIyKMfZhqP5gGPGxHs542v2Ydj2n72
605Q4TUbE1TDsFeWLhVqvf+YV22zMgd1IWqpZo2sQAmDhvmcyexE7YbQBUf3ckvdkX2erE9SgySh
Q/DsGKwdyfWsM8kgVYjBTrbkSatQdvV0Nr+MxS/qMCKQjHgjkB/2lv4MLyfyzzbJgkpnyW7pH/gP
FQS8Bq3f24hXZ84gXzLaulE6qidNYsSxlx5oJzO+H6ofMT0xUfnlxn05wwYwe0/YVm3jQSPAMDoy
F60rLccny/aaLPWbtc74tbnGXm9RMrYquMXYuMV4ZsJ0r5cnD3y0ub+JNmDkh2BaM40GMajZorL9
n8K6SlYcLbH45f0MbScPx6am2hiP2wtulyzcLO7gvfsopWEU+0h/IX3hGPeUH0iIqnSZJEF+JBTm
IKZsforX76Ae1IwsAKZaNnncyyQYZfEjhf8Ggj+miFka6woQa+BuRfg5nfGkTWCLKVHJh9b9BLmS
/MUXjzvKQhmdfqCnaFANNtGfxHCQCEZFfPR4dUNo60wXXl70jMjdcNNFjJdHXt8jX4fLHCY89iNV
Ts6vkcvVv+du0dJOGwszMCpsFPQ2FEaGZ5O7RrDrvSRrVmzjiuA57HcLwkIJLx8iFVhqRP3dUq5u
YPe9CuwwG7lQ69Wayl94X/RCJPfq8aOHvK3aaDPqRYXXpWZ3Rtnu/RZGzG3MXVbXRVNqclsi6JLu
OuB+k/SoVO1ZvIeJbW3XxKBp1DoLnfKcUGAOMv2Su6aHbnZfAdW2Gu+yiOKhgnWGe354V90AUPXo
v1t63HrCb6ej7zm5lJ2U04oKuidylJ2fkJImwN9tDaEzVTJ8VNslADOUa9fLa4qmtIBXTjyA7TCc
ywSkYenVg6Hht059i2aBp9YbE72ACMtYQ70gdV+cIPXaEXYl41WpH9OSLIfNg3fmh+xr9MVR0elf
gsOV8lbTzhDXE2YihFzpKmzsyflUObEttYlYYdoFFx4++O5v/fNBRIIQRPANRE2OilDxgakhEfEa
RIsUpviwZPMKYhi4xwO20nAhGk6QPzYnzOpRS4g/rvwgOGVcPDHBYW76nBsKUoUonqKB30O4HYi4
jQd2yLwNcBAuNyA58wsSvkeXulcFu9NEVpE5VtBaKVuQn/JbVXXqgvCrx2l4f27lYrERzIaWaRKO
89WVPf4Cd60/Q0pZtkDzzl0WdSTx8cYXkOZW9wlaeOU3Yy7fgn6yc+RNQ1ik2XXuHosaza/uZW/Y
LlbHYUuapXvdYHQKxex6Enq1YjZbnbJGfcPSWdIpT9SPODA6KCWcx3hTMbqtbKGw6yH0wEPDcGu9
nD4dUgqEL5K3+fUSBF5WchRZkmC7syFcBaYxdMUppTZ7IPDOSS30u2nhcy/NsiQ+H3KSBV03laxm
bl8b1BzAsJ1fh6LDI3YegKeva1Wela2p8rsCB+kpeZAXytnOXJ1Eh1Qg77ZZMT8SfYwMPbXdBGNq
QBkmowSMicn+0U9t1eA0abFOQcLKZNTvDPBORoA1mKVfM8jhm//wns5szW8Dk11VZy/OcazaWvwi
SM+PO+P21HYoKXjDwVcnqU9nJtbadwrbEFdFuRHOm3iqfAF7z32/FzAOGEofnbnHJdaJwpjLAfli
CO7oluI70dB8ohoPtzX59dzhNVCtpFc7/CaFkdKlcitlAnYOyBAJJzgp2gUV6T/EPJE87SYv1ijA
5uvWwZDhfvRJzOn5pBt/WrWb9u1WjaEeaUrzsB1kn7r7WRjGr/YL7rrIH+6C/oeb4nkHqKrqEc6J
534ucl7NYr7n1crr7HQsxOQe0WMtbcvne4jKxngfpcS0hwNcWCyXUWk/a3Dz8CoR6SRLN3yk/ct6
fMmbV6YlqmC/A1tjcDi7jWi4YZHB20dhqSWMw/JJi8O0/G1Ub2hEtZc5/Vj4Ap7g5vZmUrOyx9Fn
BZW95LcR/dIMegHcHVMHZOVvng/GrDWeTGd5ChdyDFPKr4QhzAD4zGLti1ju0Tmk243/bY/NOumi
DwnWRv03ZjndfWeyxsklhL/Wh+NpPWL0wEtUrIR/d70kH7/mgKXhpfjMeHdk0b7/U3UnTFjyvH8i
Q9Vh+MCyLOhUqieYfxSOgii28Mb0SpfJziDlY4OPn9LI/hWSnb3elidkE6RY70HlKUdYW4f5HVf6
4EKHBdGgzKvL2f5EbJlG8ae0M3syug5o91XUp60v6z/hB16fSTMOnthvewd6M72tPhwhBPF+eekV
PHvD5cmAsKTRcFZt534Av6G3C48VBB3XUcASLBnJFnRDMcxwicTBOpbpUIzP/+iyBpEw074agDqr
9Plr/cfjWFZXkO7/fRdbYtXvaY9LPx3xG9BU/YRylxXY1iZdXJj/42YHOBuMt3K23WEehPkBzTBc
HBZOMo9ERvW7Je7jfZuHOmxEup4n0NoZHwfZLEPQag52kPeWjoSJhE1VUa2l8wOaq5Pqerz2M8Kd
5uxdWTQboTAfH2U6NDCDC4NypAt3sZ+c26JwBNQxWPrswqq6xKZYQHLADaSZptmAdLxuA0he7E2N
FTYCERhjS6doRLc1s5r8a6y/DbRV9HmKQhmYTm6yuHXXW1wBuzmY0jK7Gl5qy0C0/uZXFczkUEYI
toGnFY0MTIhfJ/XMKd12V8OcEM2Hihy23EprNHudbpihsEdXCT3DfjgnOlWApfb7oOpVFCATKxeZ
gtbMq9ee5gUbIOUhM5q0yUKTsmIX6LuQZzzaz9PzW1jdJavqeUabPwd+JlB61F+NFSHb6HlOQsm4
8vyGZOKGUsp3HPL2I91SuUUYUzpqzn/nJkPACN0jDqJT//Q1RoOKHd+j7M4vXmUyNYnFQgQ/jhUm
NKEPeDUKVEXwPcj6MIS//iF26EjEfA5aGERnBXmfVwMu02q81zRHPZCKwtHWiF9Bp+1cc+ZmNjr8
bcEOS+e1SOy/SKFQXal6DpeUbNk1dDQ6U7xLDLxPBcYt0lreFakojoBKFB9ENeBs2KAgkgoABW+3
huPBDQSeJZRdxtz/SNUuZdFI56pqNVNF9vLvX2XUvvKt9mwX0PW7sWHM4dYUW1ZV+pQA64gi6sEa
MdtII7CtD+v/oVduCM6DY4gARYzDvYtjTfcfdKByGZmZ+iE57wcZQ00AV0qAzFCnzyao/XQUHb/j
/BF28rN74wDhRnbWaxKp/M/IlyNh3pGOlNYaCzypGzquUgPQ3VyF9Mjrc09/loSBNeZ6hqkNLTm4
NOMKEz6IPGCCH77tJ514eRNZ8P2VhAJiEPHfj3l0fby8pgs2DAv7FiQiKAmJu5TWqJI9eqbO5phL
lF4KM26+n1bnWpIEZfU4OdmkWUwgG1LjoOy4lRmXcPYRNy7NH4imEeF3dCfbkyltYM7VtIj2938J
DaMpoNeoqia/7CzaVket1WRP4bA06lFbjZH4FOaCpxMM4gO3g9zm8cxQG3myas7vRw/ejnnt3anr
idWA7+nI9r7uIyDXxA3VeZATuYQjf3WKhqtYobVi9dW7hml7KPJ6viiUi2H7HR47Tf5reNvEqJw4
E9Zbb35GRJLQMgMMa9Px8Coa83Ca0Os1Kc9VlLmvbK8I3OyBKoGoOMM8Y+DxleBa6dhtFybX0EPu
B14kphk2sphjiLYL/8M6MAZyqeJ6nByTmI9VaJuhoel7XY2wRGy/YJYjzM30BE5KRMBFNT6KN07J
9Z4dqVUS0EVWgPI6lwfSmd8z42dXwrxumctoeZxcJXRiAe0d0FB56YcDcXKSbkz6nEx+ZuVKhh/Y
sDEx2qA5zJwQeiFcF0WiRFY8n/NlDpqni0bAWQiEM2vl7axbIkDD6iZpYjtEk1oJKMDiwxBu9CGu
WW/VziDdXnyb+Di4CIUn0mzjIGrqpIhwW+nnTXMpAVCrx9VQi7mAxyiP34ZxhXVXtlhMkIDIrKai
uKRWF/lOhlgMrJP3pvTM5nRAMqT0GiF/CIv7QLzGVc/i9YxdzvthbvyJDjMc0Cs7GwRsKqdFUiFJ
D4lJ6l1u0c3Mn/ky3c7XLYttbszbZLk41FtGkIdMbNp91Yfw/61QrP/fi2jGqOpCtck95VZ11r3F
QuQG+XASWWYCxctAN9q7d9Yl4rPyiy+WT3UovTezsrjTKfaBTX0HwepxvpzL3VedarQx5ilJiy7s
hDT/2fuyDptJuHP5886/UI5BTJVz+2qA8WDa+kVWGDZoQ3PJDJCvFFkcBxKzm/4t+PJ7ckFeTg2z
N6DmIIAEWXFsw4FqRy++nUaUgCnwrGzNoVpD4il3M3JDcu3ZfDkVJuwIYpdgf6YdFBonxBDR1LNw
lwxb06H0jubkNFied1mABpXumkN86MLYlXYv1cBzfd1rSV0KGAHxANukzvS3Gt4TLx2kZsLCeKmr
GTQ/750kS/d8MfWKoyxvy0Ti0cxnmzhUtgYg2pNidIwJRDu/qRzHUyjPXWzQn2elZboOAGjcq6FC
lC27NxRqE5lfnk0pjSwP8QcXTs2z4CwDazrXzMNO/f8pHSOB3XfzCITLCnGXgvFQk3srlB9DDwrv
Zf+Tb/h86rrJZZvjlua1ZMsGbqWkKwrr563KbtSeKg0W+jENJksMNBUaeG3wCrznv+ZymS2ivqXo
sBOrjlL5LC6mCtmNgHuixOAD849rohRHgszAEAg2RDuUyx4iMqIFNqxjoYNi7gX/KoL3N2gKHY2K
FUl2GfxSX2JSCV+zycUlhJffk2JB1bn0YyOpP1/9sPvSOz0h9aZDJ8Kd+ZfPWRMRE/WW7rUNcDxv
x7OmqNLXk1duZlMyPW+yE1kAwVvt+ZHbUhbatOo0JKvWc44C9G+yWUVnUBZKwSUKhyPHBDr71ozU
yYMaVdNXD4xSN/cOrev2pr++wWIxrLs09ykTQl4KHPk62KWSXZSHzejoIjtS8qgqTQvNtcNkLDBX
PxnO5nw5CJRANZLOYksy5pXsBunZ0e45eDSS3LmtfgbwNlukvERpqf2LNv0qZaIGTn+ujDesBEPu
esXji7fKl7E7hhFmTl5GpiK4fMCgLIPLbVS3Pwx8YWpCLw3Xd2hbLUr8N8+Zrxr5+IFSbGSq3DWz
ICEIYQzPh/Hn4d2q+Y2F+lEt+mhGt5JGE3r8LBT6oTnKWihuG2lrCWZiv7FkvQ1aSfcPNC9o3rz+
S8mrly9Md9dZlV/vW3CU/SKj8v8ThG6Ys3kbkf8Mp+23xupjXut+C+Rieb50OtGn/dJXupfwBF/m
GC+PqggCkgLqJgsm6pBdYtE51TDa4kuAcq/MTS6wDKhrvnLpxAExINZuw4eT/4qRqxK98aM6G2Ub
nMV2fHF8u0VH2g7So2LQCDw4H/C7qsCQ0ZYdPEWGUCEuetOVNFXHHl1IdFH9pg2isqKTf50XApjY
/eJDtjX3HtdyJb28m2CUBDpEk2HtVkE66CT2sTe8Tmj2z8H7V7W69xTADgSBNC3yL/2PyNiH/THO
X3mabpDRVwC82khd5/6Az2wyA9MWQHU+svWU2aA+C/YM9y14p2bKeKj5yHUdZAbYfGO+5pDSrq64
9zHURpJsTLXn1rQ28muW6oAqCHabkru0b44KynCuoXGK/7GJvHOLRzGlUOKBtV6LFDjGplqfwV2L
cbUd2ittbJIH/c9stxVxE/8V/IvsbJykUNKOPr4d9fShN3DLIGL3kXlo8WUVaXDJ8lGdgkYRj9pV
2ch0CykRUrUmiQckV3e+LP4WUlU9vHUURbQtDM1fG2oeQ0iZ5RRf+dBfBRNLK5Z4c5P/L0dBVKMC
WhI7qFI7+Fwqp3E+I6tOMpmHtEhjqpSkibvihUn7M1NXV5Txbz2nTkqrOt19+yxFYHHzW6fJg0GX
kS3ztMbsW6LiE8dqL2xEjPYIeFXdBwoX3QbkdzVrYi53krno97CCWjcLPt8/tKCzNtHiuetNogAP
WXsgdHIg3RL5fEFCUR9DVMQQ+/kkDs8o203rDc03P5JCnZpiv1bJfayKxvujWZAiLTXSFU2k7MD7
kaYoSm4VL8yITfSNBGi0+7ClzvpkUMTNMMp4nJIL0WgYnngfKJubB46JdoYGt13EA8MB0hN1Ja5+
faOnmkgBOuzyL9pPA6vA5C98yYkhCfLPm1lB/kxgKlq9od5u3d1HQlKXlbDYJ30W7Axj7afyo9hT
lNDJMVnExuS5D7fJ0gAcozH92B5wGhffOjLrcw1UnzfhFH9WjbV0enHbAoeWBYLQfHUwWgZIZVXX
zeABP+f7MtBgPGCCnZCbeXSKGaZOjbKsNWen0pIxmCL39fO39h0H+sFjeuxwju/2NM2324LxcYpK
DM+WcCpeSRk9sXwgCHIIL/nwuWkZvd5LK1hdplgnLDaVCbt7Ll/WCPfVVUBTEz72J3C9oK0SvEdU
GtysE6AMIlznCHih7qWsLU4A4lm4zNCNJMBEn1jj/N4XObGU9UeYXRI543x+/9cRYx7tseDCrjVd
HCGI9tjiQiSN5A2I8ubP1sutdoiDwt0IDOcOetcfbQoC1IAKPNXkigSfoT2b37fNHq+uSDr0LVO7
LRYhEOhQu6jhGq93d1cL48Drl1AM7uEh5nxQYcxA7E93HG5dWLEPcGxkHSLMzAZ6NU5yoHdEsNhB
fWS3D7cntVGXB3zHDWwjsfFdYd+pE2kLkz1rhCkVz7NCcG3AiFLAqSN7N2hIT2Gi0VyHfTR2BFMX
kcvbCBqZkld/hrGw+UHzFS7jb/f6LV2HvZiWnwkpEkGiCkQMhTGzKwluepPYrJ/Y+Xizx8vYWCb6
uQKtJC3V2yg4EUn8VWpg5TLK10UtsYBiNJ2GXFQuOuyatbpZyRNlGlNWqnytv+WxWqweX4fiF1ud
/LigSag1gbg0WVpI85uqqy/TywhimU6NEZPkDXyKuyGm4h2kllqjMTCK1SB7pW2lfx7++5vf75zY
0oXE3q6hYRGh7vmil6JFx0VuAhtZsWXUzOiHJc4yFMrditPH7IDgKqZYbhN547+6N9sHt1b2GfGj
FL2U34fsSh1ICki940Kdogp8xiUfcldbU31CTYtxQaceRxNn13RLbUJpa55srO712/FUmA4sU1T1
f+HkcJ/zwvNQPcim6vq6m72sM/3Bust9Tr7tCogBJSH/jE7hzwl2UKwLPk/x7XXpTnytV2U2C4kF
B/e7d9SaaKVGDLLk6pjNngZGMo77DbnNuYZaXuEpnk85RaGHE6kxDR5fAA3LfuMWDHDPTKPdd03t
wunAzNXCsToYbD8VhRe6uGicGMk6Nv+4KNUVmInYk/8b6uDBFyFDoTGcuKksdDZGamk2+X9n4MRq
Z4huaa5+z59Ev+pOLCaxaV4QvJuB6lmOlyzk8qcxSqLzTjcwDXmo/3aiD4RLP1g7LP5qe2CEB127
djuopnN82St8UtyrGQY+JYr8bJLaTnEE1tJ0oILwTFNj7Yp+mwDh1pUwfirz36P3pfJ08RYbf+Fa
IxBZpigFB7zD9LQDtXOn0fSLxnARCMhiuvT+HYldjYszvu0xspITiAHdWLDRlgy1JXgrxMfABY1L
EaK9WlrbNLOSRPZFZHq0vG3DZNAWaj0emATzaZQiSu2LCK+UUR6RLtaeZiIliBcm+t0FrxL09g38
oTBjp3lUq8CKlzAMHuI7Uu2z9SwSKGzjfMRpHUZnuuDZ03oMyqmA4AWduzwA33V/v6IjWVWVCGkf
hDMG7LVBf9IWStYnUnf9Q8fCy6PsA36XSjGWj6Z8fqBzVKcbG8skIkFLJcVmoNXcLHpncPC4t18u
OwRSltMDcMwMRzmsEEz+MsJ/1+zCdjcWctdzaccBGHq/Z8blMDSAvFBVWFssw109GGKpFuHdA7n3
LI4DInl5x+aoawaem8HtP+oKOgpWskaFvCYsxdvYl4PBoGP0PLXmCu5970yTQhh3r9er/mcT+g10
Jumlt30o0QMB9J1D7AnMK/03KMYQJVZJaTGQIy93yG5aLhpxxi2rC1oJwgWBB3Bnx9fO6L9Z0YM4
NJxBVcv4+6YRFDYuvv9l8eXkf//cy6NfczCMJlH+Y0Q4qCmxy29tl+VQzOLwm9lYSREE9AibUKG6
7wZbVtIXbdmuZ8Nh18qAN3djnVEzlcweAT+igRCGqOgkakKbhVckj9W0m5/Clai7tiMLRNoUY3mW
PSfbhx7SzIg/IZu8taC4FMwK4B42QCiWYrt2mSdhisA6c8I7rDUL2P3g3+xXODE9Tf/F6PNRaaJH
T0rsCSl6CE+Qc3KIlX3wcG58Y4dQ9V7kxdNTRF1oCzOntZW5TLtwpcMy+4sD4oVocV86/ZQT898U
Vb1zZnNEGJJMQtLkbtQn4BInunkEu7DWsQaVcUzzMZUBDDZGNR9lBQ4iyeYDyGaA2uRdx67wVZPI
JKTGDcv5Pa42e8N3+A9LqYLZEbLmShvF0242TRmq1zSd+RpmnmvqaLdcR+XjmX2gqHe+beTVkyuN
5SC+D3v8QJxjQ7I0B6ECpUSmKsbnamod1pNzrwEitVUyzRiB5HcvPixwjBkXQbtF17tHllKaPBfN
5vFBRh1F/kqdK4aJEPcQfmRpfUEzMrFOXs+r/XLI8tKyEch6RBTFZoYOtTHfM+KpDKHeKyIVHYs3
N3NuDGG3lVbsflm8K9W7pUsLboCrtxKqhX1oBKTTHoQEWolSLWrmlELBOv4l0UmQCLQhYaTwu3QL
0XGeeXqhMWn8LauNLVY9eM1zujVSx1yDmBjRMhb406BVpx3ZhgBiGtYq+V/IxFDJSOCOC9nfS/wR
CiWsZc7e0KMGy2ODy5rm0kU5l4SyBJA1abyckhCtbk3G12C0rfiXJKYIn05R1RGxrDl8eB+6TOUU
tNQbhrvnQRKicxGM/DXUWu1PNIlL2sEKYt/BSe5W7NCsTEzhsZCBMw2p+qbQivbmk28M+bR20L2R
3kYqif5AlQ/KvRZw2gRKGIXbcLDIwoVZ53kQKAVOqD046zuLwBMqxVt2Vw/k5W8t+iHTna9ccMus
xfwaM+Z3mwirwnVf+zl1R7XH0muLh4eCnPtK05Q4BX5+EzwYxW1ddd3IwtVinw+m16xp9m/sFNuc
2YV+jI8wCOMTbElFyYZfxXtTGlIkXb0TADGzvEuTewkFhY76AYLt/KOsxRJZBVlOOzO60Kn/noas
o/t0EUAh/VGqfNLqVszbCBpyjh6td6YLrH9huynRU7IWsrLRrgWAwUk2ijeMhZp0VkFYqzY8brmJ
Rw3Z3JMhuvLwU1nx8cJGdhcDlfMMz6sdvInlcXtiS9gRX0gwVlftBggrUNhtl9YvjObFk2wnlF/l
cBW+KMXbAWwvXeGaeUU3XthQipmAZbrTyZOysRqxmCi5/fX+/chm6Aw0AyuQvz26qXAGLOfcIu01
gJrQbNuHM1+rEQQI8c+14/MqZGndMDt2WITgeRGNPdGEWDuB4xNRpHMqGwFM3ZrNcfgf6mDfAcmN
Yrac8i+ciecbKM+8vJCzZOgdaO+Tr53x1kjageuTkIDuQFoi/FTLii3S1vD3FgYBdP9EOD80tNwL
hT4qAewMuDXdRMkd6JCUyH/44hoNSPh+PdknqrTpeeJ8Jin2sWJ3mhtVVy4fWr1fBTOA8CxEIXyf
3RafS4LO7wScs5B9q5/CxLVpW0y1sSuAyhAQ+Ed+vwFzUyAvxfOzHi1l2Cbzsg/yX0twDk1JNe6F
JJeddk2XRXgA9JkBkfghJmFk5j8yS0ma31Mh99An0vZP7jb6PRtzzpqBYfVgD2KmuYkSeKgyFhNJ
QMNxy8vhiVIIHQunYjFoibhbx6gc+YZG3cy4yywgZco/A/p/76QSOvmimsEok/AtkN399nGf53Jk
febCo/GuuutlxCGUrwZnvZYNn9fXM4xoxDy0IB3YXLkQ+nNVI7huLEoXYHCva49u1nRGJFTAHRCr
3W4aw0ZDlq2WHWRhRSVZePCvpVNaggHTIfhlyuCcOheW4jS8NJOWA94dKPDaPkSssqAgG2cp6U/a
KEglN+Bl+VbVHxzsuiO6Cih2cP/TWl3iNXlZ9fU7cgROqxsLtAygpqCTnRyz//Nne8HMD5ThmVwJ
bXTEeOrKflECxlsZii5IqmYBm/2cerwfgw7NC3Ln6SRlM0d/RAOgxOutfircI1tTfOXE9fE2zv7T
Vcy48QxZ5f1LoSwhihrUcT9YcOhleSIoRvuoPLbkuqWOqiGKbfSPFsRWyXnZClKl3MEPVu0DXiiG
rDcDPFlTr4DxUP6S/9wwynHXFJrqYuG/X/7bUVKhD9W0b3nXEhhpRRTie2oH09TZbpPD2SPnjQUE
S1XGPkwBrKpvNgJ5eJPpy9LoT/NMCBQk44OH+G5QGg5BaJzOhEhPa/F6IwIoRjPaDMKwK0ezbC4i
JF+CHQpoM01dObVjLSqK/f6F1XK2gMzCaj9WnFoupMhWdHZlfKgJ8pvNHGHCf07K4FawpYxDE31j
zrzgfGcXmf6wawy2zoC37AnanHyiLY8Td5R19/5Vl86QtGg7YCkzN/okXbkZ4jUD+ljEHJQXAUWS
gmrbLOYeVSKX9D20qDETDd5tnx2OEbn811skEaLu6fe0EGWGe5xkShtiJyDEw41z5ixTrgqrw7O1
lJbwu/PUR0NA7R7n0YurMMQYYVNCx4+9IOSxHYMYlmmEU4t3S74e5heuH+1Xpr+rtomIE63afVlU
ihBGUk4HlXYF1jAWSWAj35z495nxSOG23fMJBy7UjS+6ZeciW4xcjiIXDamyUX28q3NyQNiS2oR/
qk2JyePzR7PJ/xth5cyoG/gbuDjRBP25jptg6yIBB7hrgcKrjBlzFXbIiSxNMC6F8oNCKbAEL1Hl
GK/rlsowpNBplPNc8ovNqx1FtvkPmG4RJEdMtb+u0d6AU+rER/q551W+lq+kYOC7efa+NUAT8x0l
NfUal6MZK+KgvxBVpz8wYKEj2q6q+Y0sTPSn0uFXMY6KCnOTpgdKdFyggIdGn68RdxeZc2iloBXd
zCF6SrMjIzhaT9vq9idwbIPfvrzxWVdiekiqBruwNNgYBDWk2WXuhY3QQmHOR7fx7nio/AhHcq3P
XKR1U1z44B3xWZUEglqxR33MC38vjU8YtZUOOfeVmTFeITD5FSEjBUduvfbFcgdO+zWsNt8lS7BG
ZIrJs9PUytugYCr5r0dOpYwZSXkFGOUujKiOy7QFegvwmCwwntEBTqPbvQkvMWNpDt5nz7g4wTQ+
4UJwUSEWHLMmCIC3hbgfb11jJZ0x5H2CCC4HwGF/lHIs7c7NwS07K35KIL6AfYSt1+E7i5jRIjti
jRewCYkG2VQL2ULSrS3tJJuf1Jy/2cxnuMV2XvhhCCwhzMeWa7521SIBp5E4n3Wp/WbaaS7d91qF
E1Pyb4aCYI1EJ4P20UXCA7ChSFrZx8kWoEIdW9vjiE/XYXqbPtmyTu42VxLTxrXNWbuqN1z4FCSy
wILl3EiCvLjVYnxQ2AQiJFAi+4TmEPmnacgrTXoknctREhcIFyzsKMhlYKBiDafiOPRrTxQLREdB
s0Nk3S2D2jrz2GhsAQXGPd/Wp8Ij6IpuDIWDsHYP8pDOASpnBAQixqhGu9T+AmuYIkssBQGT+83E
VhYDEU7turW7cLyrypiUkoPuUCADGUnPIqFB8DVvW40M0xlLR56n2Sf0x2HCkf5NZ4zMN/hxH89O
/wzhyHcD+Ul5HorM1zdUOFyDGmtp1eYR93oywmEIKpLMm0F4pXGHIHQtvCD0m68JQ8ImTft1YOTG
/291nuxxnOwhkN71UWygTpHwY9hhLhMhPWJccyF+wDxMKhFR0SmTirpbRUQOs1PnWD6DjJqtLczW
lY/d6eEcPy4Lm4NXWywn25BRps+75PbMSF2mxiqBVTp3Z3+zxxROSt2MbNBqe+Adb2tfa+YNaUFY
MXwPJZUQJRohywaPQ95PaEH3FT5jzcgubViXLA1u2ZKZLvjX1kAgABDe+BgE5hPw7PEXgURAwnW4
RUCsruS4d8RBMcOki5P9RD56wL2tk8rbI+LSDw3n4q24KxgJsuU4MqLpNKw5Ysf/50sW51igRB5e
QKkWpybJmhHhpWnoJ8Y+0ZQ3zdF3QdFTmNds2frUZe1VVdxW3P48vkjQyyA0w+Y4rClUh7mYN4/Z
CQwaUOlKYzFKSiXBQu9OzC9fQffPUjDu8MrWKKJADRAjNV+E7Ot8P0VUknUql1BwbE84IDUMdzC4
W+V46hSa6DHCkMm/aYucGCAdWGu5LF/6EPhdVW/71bPz5o24zhjjO8noAhS2q70i5teXhSxl55Dd
a6fjSEQtp4yeWAOm7Tf6YnTDF8qXByNNZBqc+dSricMmQ6lCPg/TAgXnIUvXWWMURBt2pWkx0oJz
LwoigO2Xip1MK9z1tND5TibxLGViXh9SgO/UJ+ybkZrTavmEQOKxJvWr5WGakpV7gZTk7hdvhe6c
C/feF8Zllpfm0TXPrO/ulfqvOTdfY5dHP6JiM1aV0tyvDI3vsqzWEikrW398EPHOiwctLKT6HHRa
wjmiGRJabMHy10snC7w0bUW+sXitndNejDN+dyQT3WTidUFvlkad9lDd/75GFkMk09Ki/sXZBl6G
gTonBi8qI9Y96q+6FD2HfCLwPYbOi9C6xXCfKFQ9MfMy+MQbWQf+UHWvnhk/VSzgue6S8Zum9n9d
qfyTfdq5XoZcroAUGn/ABgfvb4NxScmB3zFZGoTyDNiCG1Wzmc4riF8/pMk0UPHI3KQquYE5owZt
tLcrJO5Q0N14jzzWO7vwPYkbGaljyQt7cvchSqJ6ZyrmbZYXjULHg/3YIV+tb226WQDbJuH8vCyJ
KPzvETVvzptnyb5zdOo/J7NOgAcllNpmjnXr20z4EXpOaffNin1LuxaCMPAn61lVtbWrd7MwLHP9
pVEWGRaaAMQpxs6kj0jTvO7bbNeribN9aY4vrYE2pw/F+hFINvoQkNCjSTNM+e9hshosW88YqfaG
9ArdiuAOqr8auZPSaH3pYNZpen1V0p/iX+a1xA4CxybuKDY+vcvc+H4ryUTPx5u3Fcr0UVi46N8c
97ksy0sDRr3rb0ax/fk3x0I5o8sYNxlOxftzc45VFNCRjhH3oFKI2EaIEGbqayRjg6IlEFQrs+ar
RfyF6DoYJuphzUJoGO/AVgdVppEcXxaOfF0p/6z5anubQwIgiBC5O4ox6fAOzh8fc/F3pVtEeDDh
V1gPtvYQ0C16IXoQXOO6wh8D28DW44QpgLvIBRkvCDKNLu8zffj3CE22RDIE6YzDklSMBLPuMl42
sxxsxd9iPsN3nRtQFJPQwjXhgRtJZGmhIYKHU4W3PzS6JeZiQWBSZzBEDTWqOkpq0uLMC+D+SkrO
D5tjJ7AnprPC+qvYrcfHl13OWPMtf0Aj+q4fe+qwyKESDpkd2lIL62GSrfMDb/JXKGQnruSw+lFS
EMdzV6YuKJjSDBKiSv//L+YYJ2bREZTXSd8BmdHJY5yA4Tbg25n+CxCV1ANrBxSbNpxlyLe3HYLx
6ohVuE+7oir45LFgowcg79ZVaMLnJwOxR6bPZqIKGwvg6uj9JnKaiblDkB4k7NkU5FYLFOP2nTWc
sHAd51ioWxyMA/hSQ8qZFImJj21x+rSOYWT1B7qSvg5ceMy3UY8teqiCW/dsdQQPI9of7i3GqJ6K
+ovne7qc/6aR1FeI+zfCmo/UIRkwtZsQlynTZIDf5qq9pIoQAkDW1+Ji9CoKpBzg/1BHexXzKya+
e/vwksvP0ynitMTZkOvLiVyzpOSNYOAAXeWgMfX8szHu/Bc+/YvZ7QV2O1XpKX74acsjMtx+Q+J9
jSgiz5RMdtWiBuVaIC346+q5CQ/1ySzfoV0ZWKPwJWFno7WWlknU42HR39DmMH6o96kgxn2cwRWG
tXi1X8sDsRdNdNsr1xD/rkwTFv/B9R1Ks5n1TaFRA3G7+lnCp4zGVVzGa/smuCv2T5n2XtU4SIYj
TZMItoSrVoQuoBXiRNG89pgRhWLbwtYCgHBkj6ReI8eHrKNFuLo1v1KdDZyu2EE/gs8kouUkhqGK
gJjC3PtRcqzKdLrIpCamBf4eX7J0meR5zWo+yXbtu5CovcobmZSheiC8b4qyPg9h/aFh3z99omj0
48glhDKKtH5RRxJdJ5tmyG/VRqRNeNGFsKm9Av8R5bBovKNanlW9cvzg9QuNqZ/eY3pnYbxqBSw7
nCbMGBIinRmebXcgAr29dPV489CAOO92ppeSwuPxpHgt8Cz1uTfoUdtFkZfDunSMejYvCGTzaaGA
dMbkhPstF5b9sepJvu0r33rcYKCn6KQxyiR29/FmqDElLJudq4ok+khCnE0IigMYPWXdWWW9rETj
22m/Ggs1FgnVYh0zM2PePONFyokcOnp1hJKaqWdEIX4RSwPKujnpr/SWPESjek2tbmWPoW4DWCz3
Qw5UlgBwSusZnKV3NssrLlGLdZvw8hsiu6tdxoO0o1KwvZGiuXVS2ngss7oSiglt7ifaAbiRKBob
jVvEROwB8dJLnSN3dVmwk1OZ2toMl+ZargAfScg7gxwwSFhc0Zpv53qfP5BdkFHp/RR0Zda+H/Gx
P61ocZCyyzWYX2kjxx2Q5Rc1RGlWA2J/ZZJJ90N/TdbO8C+xrnVtPECpc9wWUUEYbzWwmA3ZvPtC
rYprlj2uOv4pFxFkAgI+pjctiRt3dNuvfFfYMlSiMpzhB0qLkA3Ttm4kZCEC+zemvT4ITcAif9ex
nNWYd7gmRXosDZr8WcA0HIn2IsXzJk/hB3ufSEVY+xmqnLXKnIH//iR4/S/slXyGgP7t1ZzqvTFj
tf+ZWtrckhskNlkBxv7puxKCNQQiBehQ4yTTCU2LLW2IN47fZ60QJF2CYOXhnXAJFtRPM4ZXpQpM
dTBt9mzqG8BUy2lE/Quc3AhDs1sJZOQwQQJjTjtrpQNdol4oKpzrhOJMwLMMHYchYmE9dGn8GsMQ
mu7ui1hx9g+Ij7E+tXNnxg25SHPcLXKjMzFclk6vT7ZlgMhEHpS5JnWnlE8WGoEVanrJspKyXwtf
59nYS2qkZ7aRojgQirAuNFw29BcmdxQOx6MIfjG5oXhE/acfwAQnjE7B0wqmk9HGUEY3L22lm2bq
UEL9PVqb7Yfh+4B/kiD0P3B7rWAvu3LLmpZiFB8o3EuA7CkQo6v+nOU82mppo3Yd+P/AvYihO/4u
AlptE9pAbxQPvCbbRaUJ+VjGm7X359w2xbyBYsig5rLiNhC3mRhhJ33kTUvqVeukgxq+M8tbires
YrrNw0FiJyoI9H98rbxRPAR+feZ13y+8PA0WAvj7v50FfLZGNwaR34sLGqlSAWUjm0cYYlSzPCL6
nLiL2KCtUqj9n104xuFFTrWTNOrveq5pAbw50kh8hcdfXjX919xDvU3bqtMoewy3V6LIq2leDxZQ
Kl+J2NI8gdP/Gsg8r4m/xjA3ObMbPfh9xZis61WNNVTBOEIHq3Z1eSZkYcIXUsxw8P2+uvsRFUHM
XdGdfdAiLlHKP007gXUr1wjuF+HFCCxrlz9EzmoR1n/uc3kTcy1uha5vjF0tbivTwPgFb3pbQzpH
tIm81UvsYOJlocGjM6J8zZk8y6uMa1NDxkxD6Ok4eqF7y+tASp1Vd5demdlbpzR3HEHatRLAf5tQ
7qytEUDKTqcGjg+ZnyCDbx6nOWySvVk4m2fAkuh/hxK7M/kvvU9sA3bshRuD4PYDb5cMwEHLA7ML
wzyRnjIhLo29LRnwbjIk1L9mh0mIKf5xkO1x3bvO4gPHQpm4h4O3rvSTQap6sYnA9Wz4H1OSwkV0
29+DrU0Xxnc8NYyvbK6hBMW2Z+kTNdDshlzSxYkGT7BbkC6/MBXa7L8Ckri8pUuJjCA0cmv9AqB2
ve2n5BtMSKESSLSnDjF5tJY/pX8HZT1o+9yJE47xqERXEeQbbsppVLS5wASY15nNj6diMv+lG+re
o2bxtJ6URMU9faSxrY0tmsINW1WDCaXBSMnRSn1Ux4igUrlh2872XI2Cfjd5LJFs4dWmmfi41+1a
kEHAJ9KCu9l0EESKimamL7vi+ZiHeJUUGaOQDg8MUgia0i2rYErNqNjS4nIwueigtBAJGkQJpI3h
qfHGNERUZEJu/mIYOo3ff7TOzfmlSOn2RXWIHvvUYmzsO+usKNe9f+k2iRbF295R6zsiHZSSZV6g
hs/j6muKsdHFHVC0AfM/wqpURGcg7haJ19bIjhtPJSXHS8Z8lWR7Om8UCIhFozhIwbzI9JimFbU7
A69BqNMkWWD18tWG+8icYHvJDMTUr3TmCiPAjdMZ9pd/FY2lHl1SrnGLXraqFsx9AuULqoUb1wzd
eBrt4vJA7VwhO8iAS6X5xisfiYtBmXxxVAQDat1dndi9JD7lzlNkvNBYCyfRS0qUOsMVssnN5Nlw
O2B20AKuPEg9L4ISX51dRvW6HY/l/puUXzuzLHoxz75pgP/QoeXEuiwKkhFZuabckEvzsYXC5L8h
gMphyaQK92Bijs9Fp1hH0oQ1PyTvdN/pOoNJtVOs7vXYtEHurSPzfZWwOyI9wXsoHTtp//rXYH+a
ovEDQIeuzjJWvSIa0J1tF6RKFkZMMvSpxrRkvhpGVPDOFH0KAuxGeSzdfW8P56iBhi8zTa7VFT9c
mBcMT1MmQ64uqkzsUS4/vYHRWE9Bzc5lFbFYa3Sv7RkAnR9GUbeCxpiWMPoI26kK8KmwdgvdyZH9
oORCSWBJW0DRl17fRM95aMXAuWvQrpXrq/RjjCTlzsdwbd7ahdlg/qDmurL+pnfA9QPUGCtv46SZ
z2dF8TELax4nXbDTlp+sdQC9B+uqNPN0r0YrpwfY9415gpQVsjrBPshmEoynwdf5xef3eYHUw6qK
XGVT5vttTfUDo8+x+UeLGvgiKtfhBtrWqzET5nxitNdjXsf/oX7O/m0wUeMKUKEPnE39SXPPoOrc
FYuQc0QgBN68mEhpJYl76ZI5lp2Skiv7kCSyWBWEjnsH+nxL/jC0cvHXFZNclSzhzxSTh575+WU/
3M0GUJat/rGOpKIaejxLrLurSzgkp/7xYYZ5Jyp9ySERfRZLL9Db8XNfCr5kuCKqH2LIhVnMa47l
/jEmU8Nh4UZutUx3XGjqQU8rzcXxhH4Iyqqpmp4Btfg4xu3c9MII6+s8GXYFSHzurJr5CqBlYQcV
qrxGRgbeKqis1L37UZ0eofeEz/j0QdUKRK3iUIZPrw6mJM7vu5Wt7D3KK4yKos0Ww1K3ssoz30MH
mlu1wZdJBioPYr3a5LsLTjp2iMLR4U+bGC3s9QLojeKO37rnm3KA6BCA/mVE6GPpxO445SLUh25p
PZXJS2Svg65/K5KJrHOLe44BxSZlMgVpW+w2mQUx9KApTFmbXuagdSqyUs7+tYXh9rEa1y8IDoXW
4qGnW5dU6jcC5hXX17wDgugFmbX0fhPoKygfjHGfjzZPze6hJgcsAVpKyCVtcW5t9HCw7VWNaWyA
Nw2w+/8TLMdrWactvcsUeWT9Xb2f6hkGUz0ie+Oownj1dEPizBHZGM56DnwUFPOVpfDhUq4hu6f9
I4VsNT9WPVXqGwISeNVquYaY2rfiFWPOk6xaAKFHfj3Xt5rDw7LsQCu7cK5SNvVkcI9mrFzbTsQr
8XvqQg1D647+SPV6XBjNNs1/1tfLyFNW4hQ+ivW+ohAGDcbI85a+ovLlZ92+HhYQ1UhN6nzdu7jF
oio6UchpV7y5nnRobky2WAOdQ3ThL4SgiOaRxfZWz7V8ZzBEhuJa5mgXIcsZrh23AUTsTRI36aJm
XnGCkuKkkQs15SRxRHbzqQCEZmS7RvrQ2tAFwW+022kEgZlRaWKSuAcBxgsEmuF0wO2c3qPVumRf
tgZ3/WylyewXipQ2N5Pb/MfIAVEorviI20uIYfrtGq7KzqsLd/mO5+Maj7cFWRFTZBtOyB0VtW5P
9yhasj6soDp6Tx5AjFadpr3b1d0OKbW06uVRfENKhB7/DjtrKwqIZ6k+i0tYcNuK5X0w59R3EgQj
ZLpR73en0mctQn5MIGpnue5VQB6lqj26wxXuliCxI/Y3gXdsSF/HApm3kfvyrS3G4pijPk8izwL6
V2GnVRyYvLa9c84GmmgtwzHgdsgOpEibZpQBuMcjf3Y+lP0c0SMTQWC7l0OiKFEIQon6kn50XBBQ
QmAHSbDdFoFvesr3rdBTUyegMAiSwo2ltbwGwnLjqyjHCivvvnod1VvxsFDSWfH9k8dpv07g3FOD
oQYpkN3SYusEldqzhNM7lB6Sz+nNp37UDXgQuedKzzB4/qEBlF3SuWQEQ2AFbIVKPfxA+pj7LQXd
6PyRe/vLcSriwrqbdYB4cb/nP84xvOvHkYRYehexbdQ1HHbGw2BSM8faB5Js3KrB2lfoNrk5e7l4
fVRfowetv/LsnSsC7KksGXd6lruJzi8XPmSoJGFHDNr0jrP7A3pxRzSmSLLkh1qXySJirFMAQhtd
lBSuQdFxcwBchmULh3y5wYWB9S3E54TQycXWONo8PubKs52p2tk8rKdmvsTRo/lMd+vGYwinaM9A
uknkFVkJel0grweH09shBxYm1JD6f7OvQtsj1CabaJY37HQGMWvDI5XFM4ZqppZRZK2lzblf7mnr
snDSq5sgdMzhda18Eb0uilXuWvwG1xcQkOUClGL30ST0NzCQ4MjLzrInqmkTeZ+HHOKPQIMhODoh
fl2Y7KinJBclQZ/O/vdtZqqWcCOxsW/8heM6wdz20P4/CbTRYKuQV7HU08N9aVVSBG8Ao6/APHXt
y8HDsub2/AOqSZ2h7zxxTcbd+WdeVQOdOCw8isWSHu4PsbXb+V0j+kk7S4qdmNQM5qsbzyXWmoin
74PnYc1fdJnV/Y7QZZqj26KuS9LfEtI9pwQDm9T0+m5azduQFXWmeKNyvFCRCZhLTzwczLdLO6BM
fOpnmfwwpOhU9b97U9TrKq+P5olxhzMoAJfNutl4w8letI4r4BG5kDkYP+yOf1Vc7a3EsbiWYKfU
Hrgu7l+4yzY5wDnJISpufEMU2yPpd275s3VYOHpQYFN6zOXuleudF4Buu9obf2mjwAT1ddn99XWE
JKv7V9exlfY7LBCl1C0iE9UtJLzC4+syhicPp1JSnsg3iSyw4nk48NPpNkwj6h4wCrtjYcEmTggL
tbhH+hgX8iX9UbETBpar4FwYPQy8GG/l2FciRApr6ZPq9u2tgYs7SOFEF5kbr5WJZObA+QGsGTIZ
v030VHVZKUdwp0ngzZLcbecUmXoraPdwh7V2kUclUZpo4rPl4EBo1wtJw7KB36YeTJQ6hR1JUl+5
HGyqMVevBtUTA3u77b+1k8SIiYxagE4+2u1kvax0HJOj4PSAuaJHjyVXNsFXreXsp7OZFMwfS8NX
BvNxWor976kOWUqLA+DSewJjfZvjMOIscz9R+KAo1t7HV+i+gKYU0ZU0Rh8jvgHpDF5qiIIEZhkc
aB9/hFsX2GNeDGC48D/2CnrTqMbgz0kjhndG8uOyB9BqqQIpbiqUWMoOvLFlKVfHXOTic9diLFB1
1hBbLAeS9eWyleNCZvS/EgEgvPO3iomx1Abz9oAYWQVmR2IFtN3RX6WUR5VSGKDF076vEE7U/hCo
eQ6M2HM69pSBaWKwxUa81BkIC2e4gP6tvFzZ3UdrcISu4G/mB+j+hJWpZRBQbWfTqABJbqLGavuU
fSNpSAK8TQK/0heoKpjGib23q5F6Y8Ss4f73Zo0pUNLb1c6vMWiXDTuOuisL/mMERRVkXS80eCBB
chDDCa8aq0Cgspe0sE0iFBQQ4XonP1Kf6E7Ue9Xomx3DWzIM905OoI3XTmJaK4SlyNHDmoTYTUwF
tfBoslydXaVloLxbSRDUzvj9+SozLKBIWxThxrnPLDB5ShXH6t5bU8X1d08KYRmRNuwR3DyrUtm4
fBkEuwjyAA8kCL6eBrZ/GuNPeQdPY09d+mNNW86MAzbIbVKwgajfMMu81z9qXDLxfLGXDmbKKuLx
ENmkDj0ydS1ppa6b6M+/xpu7Cs6pN5+7lJ8Y5SPI290tfzL8uT2p1Q4mKpbK2nFKrkCVNkK+F+1v
oy2+LCHhQPZzv/ettqD67YfZpfsnD2o7te6Xt2CQdWeG2rwdY3M+UgQkARtUHRgO/eqSNLB2gVM3
qIr+La1isW9pqw8EjMKtMc1/6E19Bm/ZomK2EYs7hzjeuISlaJMWZdHVlZQCgMpOKP9MPs4BHwei
DopMxVAWs+XKaPBAvZTyqWe9egF++9bfN/OuTxqi5drwVp/t83jIu4hRGwUPLT4+NafE/Nm3UQ9X
Kn9iO7REhwPZO5cxVSUF4Mj90UAZEAp9lckVLVV17Fp5cr1Ii8yRYQGZHrd1r9VLwvM41kSY0Hwl
/upyR4zKRDjo8ls28ciL66daa471KvotOGXCqZE8hBukdhaquWrsa/5RBxLGS7GAFZPkghopOLQL
CcYUuBaM3tgf7a+HcGqKOD3My66EjQTjW3JhA3GPOoY4KJsFRABF9Ud9FhkT5YywIAqYqRsI/qz5
Kaj619RKMJzOW8WpokCUOYM2L045TmWOiQY4UH+jLiJG363pAysjIe9+R1g2DRjSDCJy4cSCLrSF
FXk4VOWdC9h85ua17QL+A+xtz8XuQgj4G/nznOaIy1D4aeSWT11MsmVEHR8HBKawcd4gCGkoVIEz
1r7bLcHq2I/3bPAmeoOaYI4zNZEWRDpbFBsXa+Gmkfb6YLT9ub4DbCUgpF6fyu/exNUqJeJHa2zC
j/Ecof+uwfttsbReAsBkIyAqpXv6RJXKXmNXUbIiQq8PMfq1ex1YQR1qBthIAJM4fvxNJeWzONYr
3yiSmhj+mC5+IsbQvFvQO5Lxgs9+/qfaZ7eHQBSmT1IiL6h3ptJXgSDbSw3UX9EIvPsOflgzN19C
7FqhGCmAjwp40UnGYeJSgb27TUTUoexZpWE0yJKZXIgegJCZmwtBlspLlBDgTSeM06PZQJDp3UpB
d5CaZJhuHPTMJ5cOlfwWVw8HbiHqo7OsbH+9n+IcFTIXO3q3fcIay5H6yG1ToKH2LEyXQt+NVY/5
ZAWSSMkwmPGZzNbTczw1mEySlssHE0r0zMDQhEERgDJ8H7NUr6M1QLsZLZ046YAocWRwieQpwsNF
eet+k9Sj5OxUdtjYEdWuaJA8GuQGvuKyAGHiIAyNymuBkRf71ue28FLKQXAOstok9bGH2quLnjXc
6DAUi6FsqIRbq4cUZg++kM4iqrOmB7bLdWVz5Gby/t93+Iyn/KTdnGOb/6lUTqtEnEu6y+E2A5sN
IJyFSJljTyu1dCDugMrTrAXksywgVC18HA7qPkr1+v99OBuAygpQkJs1tPKNKeO7ar7iJTgKSAYZ
SKBAd/Uv0bO+EuDgDIuQNLuDagYXSVthtFQ/1rWJKZ2HQotUImd750QZD3rj1SAl9KeVWQ6Yq5sZ
JECTprJSeW4wrwAdUV+2zJd12rdlcfUfa2gLfg8nLa3V7LTIdPJjiQqOD2AvY2YKSVa31CXG0pb2
1yLrOdEML3M5/NSi5Yf7MweHoyKERnwhHoRuj8Q2leSz/jsz2VKb085M2tHKTPw+/97s8ax1fDIg
wT3hao4QMfWIaFCst/ihh6l+pad6ThfwGic0AURz/iRlzbWC5BvIIqxX/w1wqW7M+fArumfvNOE4
9sDcHaLsYTA5zHdGX/692sQLUFK/HPO9TL18ZH0wxUat04gIG1tn3KnLNXBPWmZxGc7wcdu7Lv+z
lp3JZWDciRQt/budy+V4t8FG98k/OmueDGFFmNFzLQvYOCvI4Z0JIYvP4lQpHmtFAVUTT9WSg50h
G48LDaEGucYQFMS7uq0N0scrcKYELglKKjxTt2N2hbS61i1suVmFLfKS8X/HUL1X1MOXqfCL6p7I
9lfh6EZda6sEpmyf4c6MKbYtju8lGWfE8HrYNuJW9hrsCUdmd5/iyU9GbWy0bUdSpVzazJbiJOTD
A3T/C7DD9nsUJSsfG78p5k08mBJTCmVSK5touYMD2V0Mc9IPtEOeeGCG/ccUI3uopg1IVPhmsDDk
7RiniQ7tSwIJ/EYXKvk8O/7Z3QgtPqzxCHtCO2K/n3kOS8mEGmtOZMB5VYEXrGgrO62vvUG+7dJu
TCGkpEnSR8PcJ5GLF6qKdk1+U+nelp2A/8Q94dsMAxAPJ/i3MgZ0jlNHODUIHrzC1P2/lSEnlM4I
CD/9Z3h1qknwHXENS8E1jUYiIxgp1e2ggFzxBJoUM+zbIlMj10qVVWRI5wzF8Znsvgtgd9tS+Tdb
Dzr9Ya+0K0JR4Azc+8Q/Rd+2EkiK+r7IPGdULRYP9bdJfbwe/8wqhrcRoKQcm6plPYllf78ntlVa
qMtz5wmxHGZgfvzHR2IsxfyhCd2jugb0rGOuW8UFLozHNtNrv48UvcrcvObBCEvNG44w9cBVNb8E
TXUnY3CTQlinsEVfMLuPn3g338UP96AXHuVI7uYKZJmMd7cHMQDWECOOKk/Lcu/DdWcJn61QTtiC
QPN8ukiS/fIL9QEB4NvJx2EopJR7WB1azwDHqUU3PdftNoDq7RJ0vM3mcoDVCAIZwZWbm2swSZlm
Bd/fUle4oWM945mADRvezmriy1qqfgqcsJsv8cCVj4Moa36AyIvoPLPALVP3trCJhSVuo5T8jFB2
el/bAIov+0aXd4SlWWCY9Ol/Z6x2FhRleyCV0y+9l7wiVezd6a5uaWKmvmlfatdppqKd6FoTGoCo
FeZflNnBAaz7PxbNMg4WZCdtFw5gDtIC6npqvmRGa8JgXWHNG9LOPCqd5otsoJPoGD8Ay0mvnwOH
3MDnY/q+qVVUPjqJMPTLaz2FrPUrgVVS+nm4nIjrjgdNbY3YLirzVIZVZNvPVcSbgu3t3ka4iaIt
GBNBTmWrFWWNw1Lw5iUGcHHgNgCvnIPWPoJX/pQSDiNAbKkIJYPhTGihteVO0RHyyDbr6drDJzBg
4cQKD20tbEmmTpwUkHxfMlyQFZwcqkexwEZnPFKqtXr8CuC0eGZU899KHe7zWhwQAGZzaphpYmQ+
1xsf4GF3UHSgmrkK2UJMnqD3BsdcaX5MBjF2lSal6X6liCqwziA1zenNPpIGMX+1iHAnN+LrHAFV
ec/kr+dkF0UoXH8sZgzM8nHAufcNJrdmaFvoOY6nfo5vbiDuQvCfaCZ5yjDl5aJMx0+A4xiIobHR
I8Ox25TaCsTqTF5Au8mXK5WrLWrzfLjybJxOqpHsx/O0LRsrp2gwoJuJ16wuSPcylgGwc85FKAVT
KE7cddoFj7Op+3ccjF/GmwGdS4lgDnrrlzKweOia1gt9cQah7GLfoAVSuV06ynW5VlfHZ4t/BZTG
rY4t+rUcgFUSXLbWFvknSLTJTP3I/zQfwUjPRwGdHmWH4ZTaJWwF0GlnQpREjoMYfjDhssEqBQgq
LQUcGsXHLnC8C0nI5bqh6djXRi+U2E3NKCkkKHobVm7nq0yf94gA8MIDv5BQlHJnv6DU/hI/RJn7
GNTGOVuJPe8m7qnLULVcpBgEbcMV6gXTAd1J/YUqpTKlxX1+rF6NeLFh1wUyh5qZd0F7Jnk5W9dx
ziDAV7q33wKYw1sg2eV+y28epn3lueEEymz6QTBCuUAKAJNvZ+u9KdGjC6RrupDP+MLgbPgl8aWc
u5fKg7R8yrcfj9eKwZXPZ0jMMMb2XGi8Ph8bECzIRZ6sn+CI4AvVbt70CkKkvRkriOgqxlQ8XHb6
yzvKtZvvSkxULfHi7JqcD3QkhaMI9U8HLo0cqqHPWMzvc3IJrnthczUHQ6zRroCkiIStgbl4AW38
A1v+Rm0aVf1aV98tk3MoCX6jZhBdXke4kSW5M6z15yGWwhQsewfIeunJuO7ql6dI1X+Cn3DU5o8q
d1j1pqvoENQjzgETMxPKcR14zaY/lPBf4NlsyfkeRNdrf9WU65MkDEGmedL1ZIMhuDWpxWjyjXcE
7+NTNTbyaZ2PfHzYbshSDVumvKSL+Xp3rs2C16WBpiGtVmJQ9lbn4Dx18Y2XOn1hDgMq4UszQqWx
rQikAiqob4UyQiSQ10CgrEsH1t0bHuDn3VXFLSzDU08pL7abuSmzYUxcOdqd9SuZsf8Xw/zZHmp5
n+0xTL233OBd3txBm3MnA7NV1yPT1iS7xGrFNnX53rBq3ImFRvmFGsUvLfPR6IA78n2UW27UBpn/
nww+z3ZLysxyLktdMyD6takO4X/WS8aAih65Qg5LwMFvPPeCbIHWXumay/uqE0mp0a2KcEqm7eLR
3IriApJ/qY04cUfcABWaaecIF8ChSg+1qgmJ09NuXPgasoFEk2KOECfyU0vs9wdRjCZ8njhp3fSW
iItf5scFljWEoGyE4Yxm7yul8veNSqCpN9Q538paTd0WvtQWUODQM6Sdh8sxqt6W1bX2Tk16NopE
kJs83/UJUbIBeFabskcfciTWTEGHIs4Htyl4r7fLdLvDRMcLFJ9QJT058tu4zJj3GlWlidZWHMKb
8l2JSKEi++Bth8bKM565v+te/zKAU0CbTHWjpcowBKg3pkCCxZD/+3NCYaT3nrYgXdXTlARGN7p9
MaW3j7a04tFJc6EnKBsY/QyhopdLXH+9/6XLq8PfQW7Qqb71CuWMb5OLtPO7VgOczWrDZrHlu3aX
RmnQdizDyaBpqjJmFJ/8wZDruwVqjE3ZhbNktzhVsgat/QptFwTZFPfaJE84bxTXXisZbmAMwHUU
bjrjir3RErNWamNjubR/6Er4BSYTSNqtBr/OmbabjrarafgGN6WAvtn9cUNFQvz3M2+sMhJmsuap
Fy6rTB75ypkyGXCyG0lK1e4sAUIxyG9GCO8QR8SKVuFhuYo55LNgClZPwjui1dRfvOs2eO3AqsWc
iT3u0Ys1hFgQpSuDbjHojujGjU+lUFmdi4LDK4s+gYpTBvQfAKgJIREALO/1kcMaC0TjlVvwvxJk
zFNXXmvgyWy6oSiImDphqjTeSwZ9kyVFr+gtdNVxS+0CHtml+R8H3BBoVIxHuCGHHDIHehBlNi0j
5ugYw6IbHUujDwbBBNWkdq24We/qJYrIobgSEGt2Jjjiaa0naj08JBE6TwyCSGziwTBVUbNdSlyf
tfjEcSCt7I8GggbSEyoK0CTJD8yUYG8o0Qoor4vsD8kkRLYf0eCINgcHS/k0q+nDSn+2C6rw0TIz
HMMWXpwB9PO5LI5rNVxD1UxwFRKsJsuik8TvEMPsr0HNB9rmL5xEyl/LZT9C3Fj7unuQSleHMjhy
JYsfkHApCyqruplhkD1dS2PGdDe9+tfN9ipyxeJf6PAjo0Y62DshHs4fgdb7ZU/kfdRCU5iUsHWm
PpX8EHsvQ65Nc500HYKljvQOJXCpuVtdzVSq4FJ3Cp/ysz/wjHno1xU3ZbjXkodf8MYxEfkYdkc9
9wfNBpwg3SAmXoGAHKeR49qkrKhIsa4Q1ahM5Kn/QxUr7QLQcSz+9jewsLqI4GpvXjdLLGp16FMX
29ATQ5TZeAiuwvyB57jGDFCn8A2zkx6sQBpNeUyLNxjDf31O5+N9ru4SpZVjF8EUjuZFO6tGWI4x
IcTavl+N+yixgtfZ5AjJkHupFIuSCD6x2bxUGDj6QqC1NxMTxEkMYzwgfgzGYq9LJILZZnXr89gS
+Wddx8wIVnzOHnvg9buJr7pPbq9suWPwzZnruDR0U6K8NrTyNwCD1u2pDJU5toG7XFW9ONgOvCcC
hAVmD05RBnOJnt+UE++7PNXRw2Uxqx7VofMMxndtlJLibaPA1FKP9HDfaKX8IF+WXOgB8PUESABU
6BrqdyynITk+qB1vKhoEyjW/NMtIv2eWeIudJi9tEFdsflrBu0HdUiGqsF+mUC3TgRJVpnxivy1e
IyIdBwJlzNoz0hae69vlhUPJRwQawA+qz52wpOP9IB2CCezSsLdrdkaAoPCRELT3/WIsQCEot6Px
ELMDQw1dt/d7HlWJJa4fLQQoMZR9SZ51EGeLxxWL6aO+hIghKnBC1gmxzw6D8ChxP2wZ0KJmOJkM
iFHaUKKrFTCOrbwjOymYaiWXN4KOEHLtuRIEGhMUWfBDRsbRnEw/WBxnAGc6PHEMBMuyw241w4kC
eaoOkUwAAk7NRyE/7QRkcOuHNk7GwC+FbUTvEcFiUNpCgFCrZ2clVF6KfDZG5u1xl6jwWy06WdIk
F9CPdkKmmDa2FX5fuzT7ZDsyNFs3eFOygYwdChtfD9c5YhxbmMbwbQP8Am6L9V5oqOSdtvX1MhAJ
OuRQfJkQLzueJY/98HUSd1/tB5zFbCu1DorqA0ewYnUrHPWvAP6SFozNAGQJwe2mBGtpLgRBffpu
DFWNzUTzC/wFBDuwDbbdUzUq+merDwHqKbUk+QcS/fOUPYbzV6BUG1NpsXq5sFJIo6g4yE4buYI9
Z3SCAYwifzJ6r/cL2FkqZq96VBEC+HIUBBGU+NHgXXI4QdjqKEmtOQNTPSt1gglF/Q6iW/Ey0u7j
ExOUTkEc2TQdDIhhNpGKHGvD7p7vHiJ3Jqs+CffOVrHV9dwxtl91U9TB7NPWaNNLx7jDDUUjOWZx
OLyAYbEw0A9s5KVWY5msfE5Oue5FUR1ykbeeKTybgBXMttre7HUC7VngVXrG9lw08M/Gbld851OF
JUJMq8tKQwRPaw1OPQUr6ivklCZrGf5rBQWgitMSjGueIfH+32ZTW4IOGY0U0k9o/YH0QhYtTd+P
XiTIdthjspvUyhGBPBrNT6z/y2HC7m/nMOhhq2fU6JZsVe573ik4Q8lw3gAWQ0Wa0kwV1JodslPC
qnXwDr6D5KjlR/ciPNJ7M6l1r65GOf4JXHe2iR7F0TifNr+t41AUyAyKKqa7h5Yf/P2zO2k7Nosj
Lv55A9QKIO0kzXUb0Us8s6sGmLlTXMQO/MWrD7dKE6bxVPmSOHs2bmAleNu+3gJN3vIhKnrK5Lz3
3U8S5rsYdo++xad95g9hUw9oVCc/j5tL+iidP7EwncEkyGuU+PaUdnI8QoGnOm/NnCS3TkH0DemX
8uVJ0QbdNFqs1hksSE8wXts5yEFcXRR3WjIoLOUCYstK8i2K38HVF5zlUYh15ZW5b1JJv1u00PeT
HDl8k3GKvIyeCm9YoTey1JZ4ekAa907yUS50UqBhPtOs+pFTNzcZ/LtkpsYEvx8SmDIofGZHX3YE
UeIuGogYyzAF2AsKcdXo8l+8VPGZWvbPhuxE1gUNHXXEpEYZoYndL1Dvp9FIKEVo5gRwaf8TYIap
dKEY7z+NubCu2EkghHj0h1YEft4kT4s1XWRbuqZKt6iwD1K4unCvTD2YuhUYh922vaIoKvRjjwTq
9oPkxf1mesjMlEsnitUW0XVu39ttrg/YqYLXfpTvpaNDiXdzbi2AChPGxcEdUKa6xaVg/L09HsMm
0WpD+sLwn8MnitBmY939/WPojjHVuLQdvxxHm3isKJtaSfzU4MDDNJjvcG7oA3q5QznvMMZZpJW7
B4RKUBQWb1QegHdc4wz0MuJEd3h4Ku7J7i9Z7n5th8QXvuKVkxaHyYSkj/4QDFsqzoBj+KaKu9cL
Ou5nTzEhIGxSGCFsbOjw5342iAe0MI+4Dpa8MTuWwF9W+S4ubh34XYEEyEg02EF4Iv5XUoyQt5fw
FmqBn1Tnzox1mfkXbyKLTA0jhm9dyxObgItYq14U49Nl5XqMlbbREWpaqntpCaHNZVZNm3LDFm/X
+vJ1iHmUIS2YEhgCRQdmSulFZbWLTM7gC7jrFAi0w12/CPvci0qk2qhLqan6wcjcIK2MXSBPTsS3
QAaY3ipvVaMYdRDqLoyeiG17euunqjUn65YcYza+L/SQpuHOIQmxzfBOqBTpkiU8+y1TW/5VSIqD
0WdQJG1w+cZZfsVwMEVRxKKmvSV8zjuU91sjQqIL1J1qPyj6gEAwGGYP8bAzvoQD+lbM+6fJs8fH
HrH8MeVuX1HDExyWjWlOPxS6doUttQ39CfrufHAzx81rol4nzeYp7/YMKJPDc/7HNjCPrPgbi81M
QWtArbDz7Yd9GQBsBlKcwK8a1MJIteDz1yKn/gdLATf6Z9AeXBFjh4c3rNNB1Jkd0Schk9BevDG4
0IJb4nz4+DaWdqvZ5oi2kvqtYniK7NrrFbraQfnzWVUloxYK5WTIX0G8fDxTyb22hATEy1aSHd3c
YdXkQqy1nCIqRzsUv6zPAg6qnbXbugOMvtysudghe4UX5V4annkVp1i5ax/adMFHYNSzgNqttlli
QF/Vd6rbpj3Y16DN+mUmjRlft7JnXbyNz6JTbO8lrXq7HURLIZXspK04F7Lg/vY6VLCiD0Ay8ZGq
230JpdmFdumYV7k1V1Cq0BahcjZaXezAuDFiWyV54Nv9Wz+wZ6XPMaTvoOES0zOMK9lzDsDrYg7W
V9QvkIDkQH4mARHHcJduB5PyZL/lEA96YcZ/s5EJ8Ngf9Tx+ItnL7qJXUS8BgjRcflGDd+2/Gc11
cozN0EpjEhhyUlzdLNgdo8eR0805qzDnJuXMudD34dH0kEquHASxTPGzOnhKPUa8jfuFAbsf2FtF
5a1ngUZTMoNySzXWPt4otO0+LKiyOTd2TGYMkCIswDvjuLg/h0gLr9ijpp8qMx/IRSHbqj6kDMBZ
vj2RnjGeUVOqKjmiYC8NmUSSLGgidQttqbYKE9+qMD+akjurBsZxq0CS1snwJqvFkYxvL+K/ziWR
I25npUbKUHfmaLYUGdVqKhUaraq4mSKQpoW1HHU1UbHF5M1rSnDnDk2VoO9ECcvdDQiwEt7Y6x77
2TvKealuGj7nZg3leGpAmKOlgUwqIrwmYMOmnNZQUjXDmS9Ui4FkyD1z6f/+U4wj/om7UUNJHy6/
v+EIw9/GqQVfU6/yDUPchYZOUZBB8WeuyQ+fQHQmgFptOTIqQHINtO3IvPKfmAQolvqYUKHDP7z3
xg6CTcnpoual49xXD3kEv/IqqX2U6oAaYVJ/jjYzuxS44CbhFf7Oe24+rcgpKXD7ohtOSiGsMnwv
hZRlxjLB6HRJeUDlIqtRQ63r3kHB/SORPSHarqDoxkbqSapWIl0evmn0eAw4AwEdfXEmS9tyY5q+
s0+trX69icn4P4cf2ZwHNtkOyAdHcpmGTZb3Wco8kfRdsXeSc/ybxlTbQGfwoY/b7zxTltRgJ5ly
APqkABL3eequwCtkguoRUCguyVpmTlRW5rj4k6E4a+zhYOVN7xUWLjDsOP5xuSSgglw5fPqsQ+6R
VXXIT2A2TiY4N7fJrDgtnK8cNICvZEHIgZJwatd4BV+mwFY3H7RtwwVW/a3vorFgFHLQSvC784M4
p8pECfBFe+vFkK8cpRRQRlk4quTPO2qBvD3l5c2VZrJtFZivbpKVLCNbQQh7yr/BAKJ6xJf+HQH7
Xu/mzgxKZaeV8dgEKHGD6CkAq0j3XMTkW1bja8+aMVqdwOrKCI3P8dD122jRXkXh8LlBuk6Bwny/
mAWrT2dsk5eIioMGcRNd7ZgTvgMmkLvPXpBj4SaA36fEFWm/EhA2jiPkhlNhRUsLY3I7mq91yeP9
4R6tVbK4BHL2jg/LJVldJG3jdRe7UPNqzWk3nJfc87y0E4LokI70V9szO7doAbbR8ba5HB4oqEtt
od0Yfu6rt1Lz1Jv/DizAVtT8wpDaxO2VfX2s6SAYqs7QlliMHlB4YUG5oIozN4AyapitYye+rWxC
OCcpN0Yca2ZZZDn8TSyVDaez8PNd7gJ4hZ+BabMqYDay/mF1g8dwdVK7oH3M3EbkWyXsTUttivNi
TORJ1xDt47w3SJRLhk2xf0NxAlbudRs+P7NSSYDptnd0uizc4Fyi8j/565s/byBvvMqLWumXBs+S
/yeSdr9hw7xWXYa14w0M09wgB6MdYQWx6nwXaQb1KLh7NkWP8a6Vg2ZDzMfaNPJCNj3T4rSI/RW4
PZwbZph+dwE/2VOdni54ZHFQppexizH4gg+PUpPYvxyThSpMkLMYtiUAd7Ew11Nf/LdUmSqs03rr
dgAYhinUWIeJAbVn5jv+jSXl9XBT5K+ksUQkT9qYf0+1GTiI9oppjWlomZl/FUJK6Y22w8Gk79xC
dsud4aqrnS/lVGS+G5/5bqmQ2dOB0SZxYOwl+CYGDlDDLUev8ohZkwxxV/5tls6EMuo7em2ZuEdK
uezW+8RlqRAyz5MkFcCPw1uTXtXwhzl8i7O5m054UzU0IowSUlzlJotcVpPPH/TVYbQf7bVhG71b
I6B2viVZ9kv87l+aKjLi1r/eBdbUXw5abQmdpQtx/mUio1TugDPONKNAaD4/S0lO3CxgOnjTcmYk
km2ffpiGjvVtcWjEJKs1zWCeLgju2M1JF6KR/hqWTTwUaQfDPROVRa7ycn5nJ6uG+GE8XGwFQ/eB
jpK7R9/z8X73dNJq7SPBOGX5OzRvFqQCggCVggOx37H2cg9Ys0Xs41NFPaVpY7OyP2vliCaNHZAL
WSfa9zTtM5iPmDTiyAErq5ddU+0FJz0FkQMObBwbr5kIbeaSW5v2rhJWd7EIiDZwH4NMsrelYeKs
BjlNQ/vKUh2wzqykMHRwt+C9TyF07cWu3jft0qOp3K0OOKEzY5OWZHnYpoorQcPZDzYFUh/dbOx5
ZuCLvpa7lwoVYS+pv37x8Uaf8TULxEf84xfkXReOFp0E9DTLHxByTB18lJfyn2AfVnW0D1nMxcPc
xQYSeY0wL/URTmEXsB7wTgRhDx0y3bSczvxN3i+T9KlWHrU+6zx1OfDc6HOW2c2dUg0NBfwnjqiu
mcceFmtMvsWvftO42W9lvFdEjU8DnEnUiycCT+cLvjJSEdPg8XhC/mMvGx/3DtD5rLP/7YfU9ag1
jm7BsV8DT8MRbw0uyuMR1RrsLJLmb8eUJFyOKfZCJsVQNlNLWZNewkeqUJsuUvyFuZUfM3emRfxc
DScrzkyvzuVe9KgM6nAig/fvUMFsmxDLj28TCWyTxJ+rhCnkv15kYyRRFdi7/r4WbTkLzE+1BhoR
NBLDlHV/0Xw4KYFZyskMezeYwSlopl4umADyxiIeRJ1F5JFef02lQWFLVg9PsV96ujgZTcDusrOX
Vx+qExPo1bzD1KXdxnud2JzT1KvEeL9JgLah/u+TgJQ9VqQFCX5aU917R239L+L6RE22bsKM12ww
MAWHnWtPmagYMUJRx4siHVhOh3N9ob5WzKo0QsCt3doCjoWrEJ2Jhe2utIYjOsl85IeQjRcF0y/L
YyF4Z8pfrUYArOph6Ck2uJf55eS7h1d5IiszoJdrO7E1Ol94Yz+WXAQRQmpEr9EwYXeyX8Z1TRTD
iceSYKbNz4dkKpYL/yiIuBlWPHrUGFweh+MTBjtq5vICuarn5zPIMYaZs0vBQ8T5nShXvP+NGJul
rCcbWE9LR9sI8Czqz4h2+sg2XEClFjbiVlt5++Dn7iLR8ql+PtJvNhcEgRGDV6nnyjq7cgqhlN6T
c5VwuuwGBL7DwzlFalHD8xhmYSslVgo3XnSTX+jBrA8DhyByVYYA4WK/3QJhMscTQ1BjRYzvDX2Q
5H4HMXeKeTNYeY2BkKEJttXOFTNtyoMWC0WzvdbfpxEriC1mgnfWW9nFNXikZbk8cmMhKCjehv/f
cDQeBYA/kGUUen3j7clUsq1YgDQyHT//vuHbJS6YrhDDm+V0KSRsDcKVG/5scq3WPWH5lUXohwt7
edLdyFVVJG37MmJQrVaw/a+TDfCMrg6xT2mhyI/TVpHpne3slePGQk84QJsRy0D3XnkfZd1yckQb
MU9xahP5POEvzD9B3Mq3HcToruPiGpnpGwqm/Lukd7aKbarJht3qBEqvtmtIjwE50hkgXty20usJ
DuV5sZRgSobEm230Cdes6XypjFN0wkfuTZ9Bs0HtURfs7ekzY064I+LqzY5gepV48j0p+Ed4JBld
YmJKyPa3t3WFHSZnmgxHpg8/DkohrBsNMlQWyQfDCX3/g1D7sYYuCKwBseMit9tKrZig93afbo7c
2NPK7sk/E2D17mFDkDjEgdYWJgUup3RW4v+fa6HtEPN/utyFV271GhZG7j7sQOtJo1CCgkIGzJaK
DELlJ5y6C4AEeWSsH/77dE3/j34Q4TXS3iQLhVSeKuPXVvs69L4jX+/noML6xnuYvCXn4F/CFDPx
LIv9EUPhF0V4dEwX7Qq+Px14weQwvMIozzcguSlncLSxkjchxaD4N2QbCX1KyRNdK1yCC7FQMZce
v+NgpF7PpyZtzM3lKgWBrlEACEsrFkFjg8AdZnXiEUZEJow7to7IfDBCh3+Smwtkaa+rgeOpwnfz
bzM28/96HiD+BJfBnm64flk1g96iTCxs+V7+Qof2B+GJHtXNKLh6u2xRTIEGsRRv3klaHkMfitfD
lFWNayvsLjBbj7vQisSUuWhSQb7HwFpeBRG7Z4tSZ2U7dWHKC/xZYNsX7454XEZ9YiU3y5wH4Wll
fQhRx4BD00Ac6XFvDyBuzEfo2oRv4L8xvI/ku4x2i3jAGMStBvqWNxmEtwgMFEgO29LvW7aCgHiG
d0C1+iIO3ZAdtA1l3hM7VFrGnEcHyL+hpgRUvVBc/isy4b5aesa9+IXGYFLuU4he93+tjgvG2K3K
zQu7GCoX3xsliL1cWQPrz1rZVPPlGPhzum/zoHPiyuzotiHQt6Trp2CSPnPUSuO9g+D4ucCW8+5j
q89gM7QzGHPEFIaONKJSJBSdxsSqbgYBcn5PbV9JoLM0j9Y/DMKpMXCc1Ohydwn+oNBMgisML1c1
8X+0JCUFq5FYieUY+8WrPycmIGvsJOuHPKtqJp7bntk0QDOt29sGFLhY/a4F3cfu8ixMa+S5U7AI
eQuGNRoMg+cnRgdSAcGjO4xQbSUQ2zqTqFtC5mXBz0FBxGU6CmhhMMDyJ4Yra4rj9+TCFqcBX+LC
yL12otkWm02goESUUrP6PYRPMYhMfMFnxirkxYc7bDncG1kTGSQgdwpCN7zp4Xu2BjKxgA6YfWMC
21oSdBTheAGTjFpFDQG6z+i5RN1rsHt3xIo5qepowvUO6XKxpaIR4T0mRHiJptajCqRlkYY1Vfag
g/iWEN4agQbPbST0GZkMCSEf3ZOK1CaaF5HNHIhFg5rifUQFJnmo4qX5Tns/Uja9SDRr2Ea+adhO
oeUTzNzq/FykLX+U1dE44ml+3bCNZsOlbu41mQk109Whu5EUleRARBq8HzoRKXrKWSOgm8RxlrPD
/PksFxR0REmSKINN3P/fSmFD1jN30N41kUxuoqEy23rMf6cjjRcYEU6kzkie1PQ6I20HiEoD34xe
JgK4dhsKGk7vEA2M7F3zI6Z6pgQYlXofO/Lnv8UUvXvrx8g0YLe4iWaa8h+K8slgU1g2/Lk/pQTo
PSPfYD+GJUW1uVw4aUF/yUbCN16m8jKIV8IXrZu1llfYQGmuQuEqiGBErRC/T8lTNgXn9AZNtJcC
BDo3lpe6keI2XbKuppUWl9zoWmE5TXW773325aTyP6jRBMHu5JZGE2lcEPPMd9EH+pvTpVtTl0Oj
sg1NYcWj5IjDRHvv+bVJwhpOmVqbvCEEYXRu2S9ACtovCL1xQH798NLcg+h8DKAmvW9CgU10rT+C
dQ3LNV+AaprMM9gbjOTR1zCNlftz5BAlkzocrLFDMppasOo/C2+nX5wpqb3wdHP4hWlJ8hA/8sXW
0TL04YtqcpgAThu12cNw5YmPR9Zbya9Y1PM5DrDGFLdfdSGgvkqV7bTpFRWB3IuPUmJmhNSDBfOV
cXhRkpgOK8s21l1nI5+Vz548FCUelk1+tJ5dBb/C79x+a2fcAKukGqICQXB1dukhDPlAfqY89AEa
5By7t/DXEOwx5ldDwos1urXKQlNECUgqLIatqY47/auoB8+X2GjRFDiRMqVlxgCZbOTj1WaAvt5M
G5WOe+r27xXpR/M8/mIv8GrsV0J1dVGnk+Sl4P+1kYcqKEZu6/0k5KIBb4cjjko+Mho/rqvBKzLT
rLcLJAikD3B3m+7CjumtnGZqxYZkSz5eznlH/Mt+UchuxGrjgirDLrBUcp2h/pKfzqvJljwevSE5
wvv//9d1610EI4AhB/L8eRtubdCwzDAz+1BRxkNBZXRcfQFK9WwU2lg02nPIcF7afNo3N+Z0Jz55
uL4LaEvGRIfhTjY5CpElWjFRFCCZb3m9Xn0w42z0UbapvtfaEQa1mgLp8tLnVDSyKnJKVDFq3Sa0
7yrTi2akZyZeY5N8ziJfIDzxpdQN9vH+igoFzUo0RAwGGRrt9EQfezxIG5cDP9MBOHfOFPyltw1M
zFHewwmJrEWTIqaDBeXSInnlHmsIVQPpiMNmvrtUZB1AwhX6SPAjOUOf2v0DTs+RRMPLkan4CnLv
jXB5bqlI5gg4fvuk/RhqFyxF98tbro9VwoRzACcajlYsF/zl46ceiEwGAJQWH4w8eK1YlP0J4i99
6NvBTUNhragTL04AjgMqQJ2OFCTyt7mewVj1R1jpYZ2nU6bCmZ1d4aEnq025bAey90ldhJj4XINE
usV6LPK2ciCKUnRJOtPEIQUHb9kry/D2RcDhTX2m3MZ5iia0+zwsMorX90kLFT5b27VsoXVExz4T
glmbZiKyjsZaAEoRoFjY5GVG4dKTSHfdf3nLQtHKoL2fCL0osJ2WJWIjHwkReoynIB2cEXDbxlTu
ibTQEi97SymociNKQp/oYotq4u1fhKtrc8XhAmg4JZAxbW0SKPLohfXxTuf5AHtjyOaA7Ix6XJjZ
vImIketM9uAIOTvkADi5DKqKxvNRIpeCIw/2SmN7VSH6TGdpNCVSR63qxnWcT9Xi+46Z4pb4XYTa
CytqT0xhQgsHt4khD2pFnBYUoF26J2vaIs1tdt7cDxgjvu53mUZ61eEXIVTBDL5AZRcpJQmOs+PI
Y25xGY5ATTK7lr0dTvM4tl8VDNUhbDp5nV69kTsjUWAshwzOynbWowC/KDQuGjipO0SC+b7doYpi
V89YOchMxK9mvfVdzKT+jUJABA95Eg3w4vfLQ7Ch4qBdn6cD2K4tkaUObQS8Egn5z36uOhuOTUU2
uzk0dYJZq9fWMz+XUSA5/PLzD2hTSVRLZJCJ78n3Gzz61LLSJv+LdO1bqTWZ5s0f51yRdrVi9pMN
vmunxtG5FUDbWypjT/yNgA8VHgwJ/UpVlLqvDwpJzAKKfCZZRLSTC+8bK1DCHKIdda2Qmn5C9ntw
mfrLpfAhaf8SSIRQOLbuHoJgCQNZzsSnuZHGvtEDLQ3yrwvhTLhia4erm/NPmYLzAiHRdD0xvGUX
VRZXgHI9v9iGoxC68nY778vx1Pz5wBkomxXzf6QrBbDycgTAhjCQytUTHkOud/7BamNKes88IkR8
iCQRXDVG1zHeGRmL2TfUnnLx++2TufrhLAyu1SRozmcRltrlp5q4/mVpPxRi7v5FSAYyZo8IRNds
uyZiAAG4ODpSV01lF0jRsn+0cfPgVZw3FKirrVqS0h3GCZ+54qDeMGYjJNIUH9Hn6TXIAoPDPx0T
iEJi8wYL86eDZ/yb7F4khoeclGq7xzw4OxWj+zPK4qkRBhVi85ekpNUs0XXuLuadWCdIDOFLq9Zj
C3zA4QljruQ+pT8CUktu+RJOAng3xaGRSFg1kLJ68ZRkhLTSjHTr5JnkSlVx84+zrwSgFtt/KIFQ
4bA7w2bMtySVxpiZx6ukd6X4O/ZtM/lbGcKoxGljW/7zql5eO0zVvbNXjMWb3D3N1AUIqaW5HZ6h
gMU6L8Sk1IaicZauFtB3RBk3Vr+YxysTb5fiZBHDEVfoRL+rDx0iFMqHsykMFhcYaeIxn+QS78JU
At1LrZK4YTdDc17OD+fIQDQJ2xkZ8cKqqm9j/XOSg+75nzucpNnwW7cOIMLwUs00EC95zkbEdKTl
ASXB3fnrt1MJrjgZZZo0lBH+NNqahvx5N2ZK6kuMvcpraGH63cqqGtOmRC0XLZy5eWugOLic62Ms
B+KntfeZu8O9Tg5sbBBanwF3aLjtAdj73gXyhBA82MBcLRIxO8k9I959xHpjvFnurC54NKsKnBz+
4LNpkd6pE1cqprpzJaMXLz4V3IQlTtIqjl5x80RY2FtQ4wNicd14w+H7KvAtxl9IuwNXN9NfjWjS
bnQxVJ3HOhQ3lnx2q4ej9hDLTUSWzawNvybleP7ZUEbMVgWk8P8KLSnNxdYFl5TO2ZYkM/U65gHp
PQpAmOVnreqwj4mt3josKvw1Wj0nhx3GV/Q2+gUvLHCe+WhWvPvMl6Vzp+7yhwJONKYoG5p3Iusg
2KOgDeKVGL3tfcryza/bkwR4XmfTi0eTpIgBXMEOBJQ4LExr/da8nEe0LwCvUyFUQ7D0npdBiRRy
u+4DKIQlr0xJYVlZE+QzjR9P8JPqallf7Xb8pDCWMwdbytTvucqIZlXo4CL2dLTsQCOJdmRrkEYg
SrGysMaxYp/Bdmk0m2fdLDapfzgqfOoQ+eb3sxuDEobEZav9UEIHFPePDl48Jw9wBJN0toOS68ZU
mSzdI2wBVFBX+go4Syw6is/79fuL95S4KNN6rMGY5VFlE/PJygC3aYOx9axil/AMVZyQJsmqDlFW
cILRbFcjBfUB/srmNCmHVR5laEOmIeSh5tcegiT1m/2OOlwKYUVA0+/o49uE4QXuNv6CBU2fMCCh
4uSO+iSzm5a85kIXuxtzv1yBMUutytjFSfnO8XLa5JikLtG7DBMpa6lgGcHTk9/sXzkIBInx4vjB
QlJpx6q3SOPqWKbgI9rP8z0h/L8nnDEhxhsHefNPJQaMcdM7ORQ1jLmBXb2tNnyZd3riKgvZ4PgF
m10Yr4pOoocGqmAwKItHjlNCZib+lmoiwerSWWPiXUJki+rQQ6AcH88OLwz406T0IV6949xZG055
zvmwl87lqkuoLkss5QesilCmtX9oBgfUcSRVi3lr7aI/RMRmWRQowW+L8jDLjQtw9Se8b29PTAWp
rEI8y1w23rRigDdFNIzYq3mLqxaAa0+nUXddJDqfe7vKveKHRyTIDwwsM89nvuOQQ33bJvUGa4n4
+H13iibPGJZtrn1xPw2ZIcfRfkSbXCidMOSHmNxVSxZbWMRPyJ5WfKnKgArB7Tw2/wZGMVcDMab6
BqQ3SAblK8szqVMAe6TOJOwpaL1sg5I6ap4a04mlQkxc4JK1d0jwydhcSPHdL4zwp/+6QNpLYTx4
jh6CBNFoPKH1h3xGrcfca+JXVwEIdDkS/4rggG6Yl6wGMM2ZvgrzCRoD+3djVtH3x9/twmuXrTKK
X66KqV9W7yeZERMQmzm2XWlkwuLkjq93PDMcdGWwJeOPQOe5dLdxty7w3Nna0eBidHQIpYPrG7+G
+5aGL7tYiEIpgKDbUGYhejZFFpNTo3vxnT4LkTRTBUrcbTbZFT7+d7jsrxBs2SRP9vi6ZqIv+kBO
Jxr4gAvvLoI9AaXM/ehN9Grxx7eDD755ID+Cel04iIUt9WcKbd7tS0JTrAFuV2l8NCFnIi567cN2
msIwAXVhaQ9xvQLdIIvA5Z19sBb8Q4JwNGMbmMX2/V+26j5WQQKE5087Sv5J1Qas8VIsrXbC/XLD
Hdzx6lMg7fRndQ0I5WDDVj4j3TSLfZbbzaDJd9+vDS325O7B9RcEi84NXTVbzozl3t/1S83Dasy8
3flW78p+T3hX555kyvBgW9Q6Zu+Owzus6oUl+ZAohsV+LTOblsLeX+QGjHMFxd2rYGedUcUI0PID
gpFOHOpQWYKpwsW2X0uyjDBe4rk2bujKCD+GxDT3DEKUAeZ8gDIUcHRmsbqxV92oJOIfsAgo6AGe
lcQ2RPFt76PGFi2plzm78+8eMRFhp5/k8sG+KfmQ2dEWcIxr40cjaoc5iDjKe66CElmyWbmxs1RL
l3lpOJxtciviYmGc653WReO2l1nAq2XLx2M5gqXTrjGWc1DZb80OratJj0dl02Sj0Nq0JxIjimeb
gBxyL+8gtcYxcuS88DzAIeu1coE0wihM55OSJ6KzSMXVRWEXeiUnydT81dmyLkDt/eAezru1zZAP
j0d2bn256sR4jV/+IQs7pg9oyjoYJPSO3PjU9HBLGS4sjP2HLeFjn5YArWU7YxjRkTCuSWeaKDNc
Lm/lTNK4k1CfROlW0t5tOEF3YOWKGv9Y1+g4mKgU/FT4EwWpxA+LYbgFlTc8cxPVq1TSbUHsMU0/
vGCb5EzXnLWoeU9fxW0rFQLDmiKQ0eureXQDilvcIqrthUs1VALH7M+igJihLTZVW8exv1n3hRVU
Wq38qn5BNwSldmkGuhj9tPcyPHhI08/3xBVoeE7XztF4RiLRzgAHUDqra7TWSxSu89QvqAvyBwYh
T0e/iaTELHaXRGv4B/QXoYzoujgFNZJmans1A13V4LFQCBYYTsRo0NJy6RuorpBOdeYcaapdKvnb
A3VmureSxUnEb9SzR34+7GpWkSD4y7D/CiPXn3W8q4ewspd/3DJ2axBVRobLzoVFwW58YIJKXOFd
WBtxK6WNPHAcu+rkR8Z6ACx0I7GS5uywGu5DpNZ9JXAbUlPJoGnY7eo+NL4rx/TKuaa4nokFcpGy
j/mLfw6uM2Wx0uwNwHV2Pv0g5SnDTDwa81jlXnCx8vGir/nruupwIhgDuX4ZOBVWWSzJH8bs9xJT
bJ1m8Yahd2mqTtvgYoDNdk9aqT5uGh4gkdHzNW3JH27LiIoRNMS4hITLmc3BZLkuISgX3drHPbT7
S68cudw7awTbWGnB3ezBtHcgdla257LRNTcM1IqkBISmdzO1OOiccwA+IeT4OlkyoJgztgHSId2m
ydTTr8O9K/bjUc5LgeCOfMaWeYNxUvhzHa0kBLJZ+3SjoXIWj0TpXdkCVrZxQ5dC41Hzz2BCYhs4
97NYAnbkiBF6ACxESbnj3OiXdIht7+eCMAelvvtfIxNJpq7RIxiwfGRnIokpus3bwQNBEMfBxVTE
tdgSYyl7EMTnzV4uox/cmASffA0+PK9L1AI9FgQYxB1KWI1JcLg38VGEzjYDi6FocsK+nbA4qqbF
2BVmiWBhobbxipbzlVkPVVzFoaAJGvw4jbOH5je4DPV1H80qFhYaUH51eH57gp24jXj02IuwtCXE
XfAA1yMzz2496kYI0Ui3S6JudOIF0d3BD9s8T7pYcSCkHNXOBlv0DwbKQCf4IJ3n8UEttMPQz7He
UepfN/29CjjR/2VjCOuxKiLWmDz334gaJluqRtB+tIrIGS8rglpnwwV+3nRHHX5M3i+ql2Kx9gRF
MUR9MVllVAoiyyaWRSxlc7ClvSB7Pa6RmyPHHqD4KKefV4ZMNB4iNCV3wd+yj2Az4Czi24ZJhD++
69KJLMxjqhrOUzEcNoXFbbRWBk+qwY0gobcwWqwruL0n1BXxD8ue5kWFykH35SJet1gWgD+zVLEM
fRbYkYiqQZPYQs8wUPp0wPLzUPPIRR1A6Mn+FbwEz3fZk+86DTlmP5XL2yLB9QvON4MJOfvZcwgP
3n/89msfpG1qQ6sIREIxyOX/enXSSgWKINABFfOIsVLXKniXer+4WUD8mUdFbXX/kL9xr0tnt1CM
3YzCRT26xbIFpGs4qTJAWshdxNhnvb5PuYvy9b8UVJe+do+nY+u9M/XylBpoeKJrZdwh9t8+zhAc
fhPTUBHCSluaiSEEs9HOnAfe7T7FlcUxauY5r1Wki3pnAGWr7epY0Ppa47I4n0ysCkM8CT1KUn2n
8J81y8WU8NLNa+xGmAgXO4JaJLAjsxZLZNAYQ4M4BKt7QlCvJV9M7RV9/7y9Vwj3V/JAN7iHuViF
LYFK6wXh5lzoxxWfPz2hOX+drNfJzWBFTszLThOHIhSTgNU6Knb0SPKJcosNEKcMUztL6EghM8rq
w77/omuyPGX15L6nGvsc+5ZPB2xAOmHptfWxf/joeDtMQtnwwgqHHrqlbIFz9E+YDOFfIBkF0RI1
MPESzgUAkYN0dJfrhIjslk3oPn2PeFByrtnuyu3ZZHODrxoG+IY4ouee9kmzyZtSDSb43gS7gx1Q
zfgIHlKqGMylRdI1R7eGd6r8BlFkj2V2HrzH3cBnMQSa5ZXhJnbCaTgpFuaNeubjOZnVsGFuHz1O
ie66ZtEWkqXUdbDHYkWU9VhyBQeCdcVX4T63qPlJLOKTO006dKXT3gPo32hWUfcD/hR0sAqejU/f
ZahR6Ad9qXo9NTSWExqDKM0uh+nPT5Wypr65/NaMz4A4n2lbf1tJ9HYSesQnhzR/gvdUyi2BVkiC
eei2Q3+z+69lVkbV2QH+Lwwc7HW9bWUvirfjwWdIBm5nHK0MTLSoKmRqBLrrs8EI5bYnUG2UduJ9
4ql49S9SIhT0jhQ78FzSoTphZ1ynQxwHst1LsmwLlpj8gSgaN0NhN1Na+qwbmf3P2Dj5Cp8JfIaI
U4fROXk+fWmAQSWqj68Un0dwjJ823MzmXeOiOaT0bHFEwpOAAZa0bE+soyuZG81dtDSIv+ubikAa
OtBrIZ/cxqR7SV/MaziCLP1qawhXtiGe5XEO3cveke+fk5EAACQ9tr7z4eWUTlBK0N8TB+0ktmSe
Pyg2Kk+VNwpMy8X3Aa/Kbpgu46paLdVU0oa85GeXHGREIvg5eAi/1K1jys1tVP066nNYjs+95bmd
5QTGjvPnH8ZiTOXwF2p/tiI5Kw2wDhdTNdGdlFNU86Nx7cdSXc6iBjUD208XDpev/EQ6YBkpudeE
STXn485jnXF3cYGqacShcjqZ4Uqe8Cji/DaL5zuLsv+ajJXjzK76Wf/X9G795yzhw7vOSqEVYCfl
BuxPNyrUwNEOQYq+otDgsP0D9KySXEQQCqe0ECPRzzDq07PenBSH5wSHY4eREpINqpYGdW8DwEcL
brnu+30rYrQdGyzuDXJTEHvf/Cr2vUlEBG/N1fCzTUQcJlhceihBkq811pCc8oV+PHuGNDHrElmb
heiDtFh5XwunEDJddsoqHC4l2st6koF1xKL5IdllQ0M3cp0TQ/ttYjd0GiNKAGgKPFxsSATwVqkT
sQlyGOlzuI4VPCPr99NYN1vKYo33eYU7ykobDl/RbpbKR8hZkdxYQBuavWNT+c8Fx5VucYY3AHj5
JHfJzl9c772lj+6KNMIsQRbAtbWNGlH/ql3/Bqz+B0tEYSbdW5WwXukgxsVCMEYxSW8jUmtCzyMI
oxjErEYgi8Honz8rOY0BCWd0TuwM07YYQRqH3qsSeAYuHV0rx7Ny13Qtyb7aQdEf1lku/kKimCLA
G3AplEYzl9fEP2zszj4A72BDe6MFjoy+r9L5OL/JVTTuEADLey2Icvps5o+UF7mrflCMpFXwJfeK
3rWmYz+IKMXAjESdtfwR7QYovewnwshQAZRnzCSyZjlehk8TfD83zc5kRyn7gtloJVSQbqQvYIw6
P0V11E6waH+V3+SSPV3krZb0Cq+PrpQBaiSypdYD2SgeaLRZ9EyehO+7J3ZukpR+6kHMUnDdqa+L
38pOq4zVOYxKybmXwa+TZjd0ck2NoK5E69lOwf6lKjVbn6ac8j9RoN98VUA/60JwSGCI3b+5AVzn
ej4O43BFqj+0zYT48r6kM9945olld4VREwNnze4hNYmXyU+Md0ybI9JCFTNyTS62df1YXPJPj4mH
M6f0ueSH0ZBf4qj5+osd0i0dP61RlSkjcZ64ugE5LPVugt92FSC8suDz3sf74PS9aAbnxsSdgNNo
OXqKEFr0wRg8Gh6a4P3QBTZLBdaPIKJK+QEqxJGlWwMw4Y/l/6s9L20ee3B8glYBTE42cltccSiJ
qNxx9eAh9ORci0Bj//6jfHiqrEuVCeyZ08Hkq7K2bM+9XNfFP8YTtpzIpU2h2zJV5DKUYdMW919N
biwTzlSbhk7Xv7eXpg4iAFy1sIFqRhrHQ1SFl5MLqAZxpoQgCebsgdK8v7o9+qgkSeQpInKzi3rw
4QQ/v8T2AHFOsH1PcK/5yuYrb9dqfN5xl1HnP35SbrxvIbV0lyiyrSiU2a4USHomoGrZKKEQVzCY
pIBgSkE58xGmWF07fbkZn5NybrMxw6N7HXMLEmcFrsPlDNHhRj5D4MMNmFgZjmP1CHR3y4KwmkSr
phsZCSNMaw1wl4E17gDrNqeDb3BLz3RkowrSuha6XaXeeOSYzTtE8BraDs2JxJA9eKg/WWck5k/k
64udEBcKwpzXOVb/grnht+BDl8RikIWhIbp6J5j2TFPrKs/ns/5M/3u7iC9exULVNP2lGQr7lR40
pCY6o5l2X6+b9sjuTrvDK2vUVFQTTodPBPhuS+8gKQDNqxxzufRAmtSCeoBdeIEEodEfar0nkRch
acZNbuy6yq/NGX6nL68e6xTCYzbi2bFdGvLgL3g1vyBq/rU/SeANdANEUw+KiLWU0mPtzUItcJ6E
HyepLObfD0chZe8ezmBM+ppmgubXnh+bAn3u/mgnwxnnGwhcpsEEoGkZUSN66/l3cS5ioqx+BuDO
SoiFImp7p5M+rHEDsvULiTgOfnDhePxOqZFFHPwe0apI8K4h04lWirCuYvjxq4IyNO/PKbr8DPwF
piLkJom+J43swA6+uLrZ7iBl05uql6FJcPCDOKjOw9pfeaVJt33qqCxksjFhmCGOH1IxR6aJpGet
kopOxY9h6IgTi8U0zji75MHanXLPwFD6f9s9L3c9CFeDdGX0giMCQ6OCX+bjgMuMoHznHwb7+efe
lqLiUph9fqsrfPmYH9p0G/r6ntYTdnFbCpXMQMeI1kn3QRMauX8G4nQtmfsALvIuipTkRMQ81TEG
eO6yI5xBl1ttdd8eopJCdQGUCC3lh/j7KoYf+0gZD/Pej6iVTHDV1NIR67+ql9DdPR28h8fcxJBz
4iS1mSqzCt5XWjgAHHty32fmcjxUIrPwpekrZb2hApMT20hLGWCg8sLS61VPeqY4N2UJbWoEsEKq
+iVfAHVnNipe/3wP20/c5rGeYl6Vpz4JMaKhOV+eRlSSNG0NJd9X+EUhYpsLfxomu1Q9+CwoJI3y
8hE5KOSleLCUOsImr2aWo5PWwkZ9+Dyn05Op+KZnwEh19Ubp2hcToZ3FoZZq98txWcT8N4gQj4OU
aQgotoSrGPv/qisaMNBFgX1HMVdb7OEP7lJMRZ2RoIRlMYIR3rHm6PWJEMMbhOcZaBAeSNsYJ6QU
hxWPRiJad7WLeSxWOSEwuxheM1xc2iFwL9gfEUSrPlHDt2pBaFRMknX8FEUnKr1ccExgFEQG6gan
reBeMKpEVN3xgBfgptCAouClJCUpO5rqACBi7a4APsjOHzAr66C6lOP6cF4cqizqlwHLFBFXFl5a
V3CZ1tiuYNR0E2+uU/hDCxqndEVSSaiu5lanaCwXKfdQUgFscQjnCW9chS/UITJwgescwv0U0xUH
7cJJ+U909pz5Hi2ZoeOvoy82PjSeda8dZLwbqL8mdWvpTi5K+JOmo0r/69fDjA8Anjn/wGjC3LRR
DvD7bX1jhC8p4g36Tma7G25XZyTkxlobnUlkGPCSXDFruUih2sj3WloQjR6rvI5S6BUOSKryi6e7
YHdPDVA6epHY9264KX2NLBdqIaj11zjEepnMDPyjHYCXlg5HiroGe/M/ESgOe2NRWB5ue5oEXhpi
I0OVdWxCabreIVg8a9hTi+qPbVTP8gJsJGGvigZAnj+ZAL3zHOS0G/R9vdhv/+CF9fzmszTnGJSr
4rtCPqNhTG8mqdJy/bnxd3C7HW8rC9693ukyHeCJQgk83mVM7FSFqiYW1xrkJsEUV553kbwga+n3
hviHR15lQodKRREYVnb9NCTNB/DgxLbbNyeQib4PIncGP1ITH7XJq/1lJ6OaIZmGyefPOHRfh+ib
LTzdROrWGPCY1wYGYo+HVPATAcQlvAV1wK++vKnz39ny1AfQxisJIL6w+5K1nKQpYyqJMj3I3O8F
wWw4FiDyGx1FowiEfDr7ESy7v24ZJqVcqG7nilYtvnDTL0bMe8mmA1Q4p4kEQvPaxJqvGRgodgIo
3YtQagzHyVniWOUaModHrOdZymJ0XUVubwX461I8+ZH3hYZZdjkQlsZZLinPkVzUiGR3GB4w8D/T
112VpL1J0Dl1xEckWUDmPyWDAyB/eCKeTEayCFc3IepocDtuuXUprapAgUQuQXQVAFnnxLWkMq2B
QcnYCyCMkDe11Sxec19ZJ8p93VkxBX32CGP0/Ae0ha0O8it1WQtR2eIKQ78uvqKUlXChmZBowV5n
aulOKavaHM+3ByeptuwhAoWiIVuBC1TOXs8myT35OvuIdpmslpXvySZR5UL55/6qewEAXi8xP9dy
H+UoQk+MbvsD/dCaL1f9+dt+pIYh7Oqb0LuViHsNXU2TonsUnR+jy4ZhWI2tPHgCSH9rDyxi3wuC
NGJ+DW9J9ExQikR+lOsJE9SduJpk71biAUNs4847Hg/F0xgNfv5uV2rF+OgKmF4nkNDuZ4ivIFvn
Fln/kDeZVqz9qcL4iIVDNJkFSxc+SFGJldOGW99pcTyE/K30afG0xFGB/z1xvx9VsRxU7B0Ffk0L
NP/PYtxnuREKZ/Jy1xWazvZTe7aZbB5TI1aixuiyuH1c6KyiEEHPyaVuwkPzAVJUhXQ0tRSEXpiu
9FuA3hjCyAyOnHpRrVuakcrPl/MwROpPNMjcSJsUcmZuaGa1cGBtXrL6J0SBSaOctqwFFxh+xSxk
tiMeaooiWnvtEOHJKZMIYMxr6XA++q7jJD7WGSoTkYsSirmBG6Dnw1aO1w0XTSpxS821IJFPG5mV
To63tAzAVHMMOV4MbR0qfHcAvP29fYJO2lIWsK3Jpj1bMhaT0mSLacGtbCAXLo7yuopm3MfuH7GU
Zo9F0q76snF8lThxfq4T0cbqlE/uo54ZpJ//7CnM1Qb5aOWbs8mCoTNIkFg13UqoZDnR0RWsfQbH
T4yrZT9fn/yarBpLV4VCHm32Tw1/KsFx+hYSeC4GyFAJl6JmpSCSV9LRiA+tGZh7QU83L/+uICpa
J2XIP743SS0SEaDuaosXPFbLbV6KVlgmJZkeiYLfwEuirh8wXqfy3L3Kly3TUSjPgsTDfVyjmg24
B/t7j6n7PQvTgIOgUuW/S/6UAp1RISC4+JbE7ucqqlkoEyl83qhhQDwKgpzXEoXqh6/gB21I9FYK
0sOcsFIaeRpupvZaw6W/lVpoPNduHIsw/dwokQ/eyB/uYgNhHip/Z/RMX6lTpdY2EOqOLEdjEf0h
3RIosMtxqvO0Pajd9ah+bCtn3kBevmk/rodIoSZv6Sbu0rQvEqvi/tvtacGfZdBy1QW+af7DtNWv
e1r2ETpYSqm86y1EzWiFK62Z9NSKSWkCGc9yBdKRslrkpVYVan1rxle/Xn4AO+InVD0atabP6bSB
c0/edLk7/Rl8EOlL/ZY0d1HcHyxyyG01Zr5qbiGLSWCvOTh/gzCgiLkysr1SSYQftmHBy3DlNMIE
xZhLmyI9/8dTNIAu79jgpnOeqBQmqnY0cRsu0abYEpA8V3ir5QE6TKKDGL3gmIqbKSP7+7ta1rgk
52NqOYVIdpbSla7dvUFN0zKPVJD67hO+pWelZGuSYzcmduPuNUGAkGF/R5I5grtUG0AVu4D7jgOd
L/H1BogYQQucNuEgEaPcmN3Qkziq571Olwrijf6tsrT8p5rv5c6iFpUEo86sKOmAvdVKYKPwfnZ+
IXWTPYhk9p6x3tnwuBcbAZ+23kVivoyOBQupxG0AW73E9QGhTG5ZvNSThbRieHIdGTzmKTsNxgZp
TyeoBpJAbeXZZPjl3V+ZHO4H0xUVvmL6YFi73eTkzWal8YlgNqlxEjeNciWOmzTdu8QkfjJQVKYl
f7jCYSdOlmsxBE0XDro8j3/3hF1W70J/+FaEs1e9Kq9oRSZy+jYrdfcQ4n6N9IOcS0J52nf30hmt
wkrrGPoUE0qtILhAxvFa0KXaobPXbrQYtE/uoQ+e2+KpSAbsoCkyV4uSNaupf4cLexZrvHNBIqX3
bbqmkdlaj6b5a+VzzczBkysHDSJJYrGpWa3ObKegPokEdb276QFxZruuz7YYd1Hg+Bw4Fex6b6Pc
4RgfqvBLZiUbMt7m7GO3iA8kQg41mgT2lWMHcjBRXgXBcwgWmr2QAM5GYqqXAgqF2VKTrhuboxpG
PIvzbLMSjQp9mjtrkHsM2FtjfSUHK6uBKlSsJprMT98AKTqTLY5H0sv14QOMd1dJCfmuEaWVbohh
pE4EcVRydl3yQxOJ9rIapKlMTB/Jt/HPqhveb9eEfoKCXqC04Haj7b3y0QEy/GW+TYoL+y85a2bv
ISoL8sg+kMIUl81O4/gmKNkS5dBUO1VnsZ/3VcwJnwT385avvOkNJrTE/RY4mOZUlV0geOOPS4gA
O6TKKRwFM//WZZFwI+GqfK1hL0Du7wT5o4T44ChJhrm4YhNtEcuM1KsA/TgAU8hGXsw1RZc56GjW
/qgRS4hD87YBJUzFcohBTyO4RPuzDdWnNNAYP32lNpJo2LGOdN/0UUvag/qG2bcJDqZICpljcq0I
g3KXa6uXoTh3sCfvJV9Kj7hAuP7m4IbVuP/B2V0ixcnE/La8WccjGev7AVdzRbR/bbqkCoMkNlvn
ZO8rFOfXfz4mqjLKnGit5nZ6bjY6L1D9ozbjdIJNDHCIIGK7j0YnvCZi8T+ckT9ZX/9MIh6xOlrH
cfxT4GRAmCUxtbvySAy+k4TLpkXb4CYC0T0q9i3iXAQO2ObmlCQkHuS09hU7zEvZfJjdOHxNb4cR
TaTDutfJWc/O/1qdtBxmxVyXMw6gyuKNAkpXZy4G4UtXDhjtZIJMjClF2Ctg0y2qzawnJR0XgrzA
8Pe5yolFMbeAgb4Kgx2vqsfDOycZPn27WWC7vmasMyH3CwyFHOen4UpLSYDcRUlHBoEwWzO+T/Ej
GBsvBEp96Cgex2NlDhR0xeqg2oyaqwC+8gIGebf4hRMtamwSdzubCABUWFw89Z9+gzNEzqmbDQT/
gnflemnHRB/2A29TovBejlTVxKO33mQyxWNFWY43z9oN2u6hylpaDv4jPA7aspFmiHdeItWJ1AOO
XwJ8RennOr/tGN5JGQ3QS7UzC1YDtysDcbrDFr9LzmSPM04b5QWeBKvpwWdChsf0FGaRxKKrFezv
BwBwi2/INaKyeikEMJqrIzYdwDqcIZJX3O7WzZjaDisgBGqvYP2TY9UOcH5YnYrWlPuQcjZwKsyq
lEgKL9lbd9OtuqvTsHm/M4br79Q99AJLFCoGKU5raBK7U+/ett1UQDJkIxBVXfvG8LpQGpB7HuAE
YL9MwPiIvm8aInCEBA0o1/8BIF8oKyi5Ztr3IDNIr5gFjnYqoU253KPcm1+qU0tJbnvw+SqnvqZz
fOYBI2bDlrKrKuHc1qejgudrP2LbvZIuOFi0UI6o4xO8KJADUP0z1zVZ8b7A+ydT7K2zojcZarGQ
FdEfTzP4uLcPvJD/W2jXHL50bfh7U9TTkZR8GjACxP2K4ZkxO7mfF+BSipSlEJZBJsHU++4aJ/EY
zM4kzqAn0FOrSvUecPWVeXz4O2uzUWv+HmCP8jfd7h37rzhgkW0KFSFSaCo95yoX9GQyVLMb2n3j
qVAkuX/CwYlZf5bKwQ40krVn9SfmPQ19MMu+LO1N0jVZpfzm9PjqTIbmwTpyy+JwrkM9Og9CCMAA
WH/ovqRmlwvkVjFYBmFjf33ah2JbB/XKLJin8JBFAVB8f+wr5r6UpFoIuyurJaGb5IMlcwVzYLST
HtSbt8Gib+OAg84b9ppeUn7jxgIisTi35FmheCNaEPecCns+aMu47AxXP3XTKnczoFvbiM3nIdIy
l5YBimG7C/AFV/VgblaHjH4nKgski1Oh5ivnXw3kgr9vVkd9A5EtGFppQ2ZJ9js4/wao/AhXkbjQ
PfKhwrXmd2qGoaDbG4wYThujGwJ3xKttbMnktarSVA+w4ZY4Xt8nOJpmJmr+F0PVSFbFp+BQCWNA
NhEllV2WRXSmaFGWQXX1z9hp1Rrzq8Ua4I+HmGoGKM6wTLbnVfvbZ9PVVUvkkA5RjGY9txgSxZzN
R0JXP3TjLzzrf7RX5CAjmPKv3pgd5XHdtkEzONOKpcfrtdQlX4XXh/rnOU2jeyMr3qK/vCZPUc71
ox/gaCcWw6aBSVBgKtgXHWQLS/mGbUZrV/zrW3pSh/lcpg+Iht52SOF9+wbyxfmFUy6XI/xV8bin
e/MQ6Or+8BiJqgrQwNcafmAF/Xu2k0NPPIRNhSy3tg9OMIlMpg7MZ/M5qBMkV7xOBzO+16cH/4w/
MXKxc/OlI1uNFEwcRwAZF3Vk1j2lGPg0EEi1XRtLutYxAZ0ENYU5s7SER5tnj2ZBCaxCA7j3QZxZ
ax/IYCsDaK4H0dPFukWlTjSUan6ukdzqMzrYrqpbClWnza0aqz1zX00JtIkVCgVecoBpBXYLtx0d
D7IzGU4EnRTaKg1FiH9kFagOLe3/FgqdrYgp7EbVraK3qi20p3RSg4gLj8wWYVu+XXweZ0EM/05S
JrXJhqT4fVFaF9KSZlo8YV8SZbjPXTslvQC0ggieLpz+skLgnd/cqFc1+KK1Ea39UxG1O33LfJBw
5rpBw+/ymCV4oUUc7PXoQboFwZXZzsORz/u5FIl/K4d2zFbY4rHk7R/mHFAzYTKucHMDFnT314XS
gSL7MOy66g3aJZbQLtSOJTjCDe6MgxqWBHb+linytmXn5Fp35b3Bu3/BQp9C0iZclayCPxY6HF2V
oHg7sV+JmMhS7lmQenWpKbRMxevBuoKj8otjDMzD/w4R9dMKvn6/BL1kKgV58sOLSqosXXlBE3XY
rbP6furCwMY4iEOYvqYb0lp58FymtYKMpxqsK2p/AfTZgRkKlYWCCN8akAWewF2FV464vE82w2lm
1WOQ4ckpAqQaCAoiFolDVXnZL3vq5U5yKGruMsEvmuHFD+5Ugq77vLI9MiKpoPaeqxwQ36vysPwX
/VwVpD+JrMHLAQ+I42oCYBZ/cGi4Byhq32NsRB83t1VyffetRLCRuD5SGcKjuMJs8Gy9Tua3H48j
he+icYuA4Lg7C1wDo0d8lVCKZ84NEiTkUa4gKFgjP8Tj9FxgTl5emAbOiSE+HAYnXBOhU6GVo12K
aNEKsaNxqy8xCCzH16WDzIB2QSOs6GdGoBLFfDnf7RU9jMcj5PdpW6MXZF3RZGGmVL9fvDq9j6CF
cD55zJ52CkVmJO6hnVbWDUYlu5nQonucEulY6XX11N2Pu2Ax/FYkaGIZ2iHsxhahBJ6H5OJEnXmR
AzwYrwH73PLFHlS41l0u0Ntc+ZXNlhNQG1sh3kylzVN6pjj78WKSBDtXwjf6lWClYvdczzomrQIf
5YExJqng66Q8pvqSlnKoadWnlQGhV6QHgIz/TwCxc1qUQZ84vEPJ3boo1a6HuTDJpGpSXiL368SS
/Y+Fh3sQVHspARSTkp/0aj7ouXB0EGkCRkgm1k1D58vGxn6XPVLFutlmkMK2gW7FQJFlHKTKSVVK
5PA6ZuitTYwFd9E6ZPrRJPAXwKv78ahfPMeqr92dbCB5t9jGklyMQPCgP2JbJiek6HSUAZ1hzTk9
i81KbBE3xgT/45ROI9P3Q6pxsHf22YaekO9Ef+j+SAR3itOZ50rlzWkZ/U/qUISyyTA3pnvPRA/f
xfK98/v4tms6SU9s5NwnIxRfkaEREcAFETw9fBYD8CJx31AeT80C5LYOPKOPHlpTZUoxmrWbYCk9
xNFrigK6yd37MTSMcMKtECKFerrCjAZnPA0oRsiQjPZB2jUU4dhJW5dqRKzVEnYbwOzNM93WUlXN
LmkWDAr2zQ8EuaUfy2P8Z3yG0YKwZkrTTyqQCUlVWmT0LlNdCA0tYjP+myN15npVQnUc2Ns6Xnvo
O1d7CpxBFhmamU/KLWDL2WDOXfZ1/5AAqWXspSPHXs14gLanmS1h+ig3IS/ZB++Lf0CgU1xE5Dti
w8PqyMk3ieAmHpKlBJLJkz3i4q3IShvHW4djnl65ZkDbRCDhRJAcMPIB6hhl2NvRs0LgYnc/0xuo
3bJiUHrbOcGY0RKwbLieA4R7VhoGiPdOPU8w72sQ/1E4+bsfi8Ybxg6iMuIOkEukCaTj99q59iLK
mCcCs/MiFWpzQgN5Vnt1RQIGkvnWXYgpcPYdB1pKwF7ZjpX3ZUrK6rjCn9Kt9SHXz7FEBW0EG3Zg
WcEfwWdp/k2KA18Vui0bLsz9U60z+Gl/mUBCAAwU7nE+xLYeO+leQ6g1jh/txdGv6fRt52gMlHEw
q9kcvnJeZeuh0dmynKzZghSiFZ9pr/IEHPTjWYCOO7UdDCxPejMHN7bZUwZcAY+zyfppNNVRRwZZ
2qOGWpD9fAMTVRcTEDsLZDrlOpU3PpUxu4wslezjj6TzqvhCOdvl/uIc6nbq3BmifxNbtjj65UNe
mwvoUMftGIxp+5XbTE96ipsBwpjJGMRGh09l2bgVRr14obZs5S6vsTOihcXH26J/fzZlaB670a97
yAfWlnCkt4KQcY1ogsG4hs+6B/jPTPZfs7+vdnRAs5gvBtIAvS7+oY46tUu2M4loONj58rpKbWAR
ApmgP1le6C879bduV6LHLfPTgcbmDrB1JVyelzNsuZqI5eQAG2G18iX8wAN/XIvywjJQdmbULTUI
yRN95TIP0QD2uIKTPFrXZZUn6FFFdJVoI9P4/5lWfDGDC90D2PbYKLV2BK+1MXzdSX8ZgDojLNtc
Ri1S5m8pJZlUwGCkges4NsWpT75E85HrahRw7M1FjcS+S2lFrfA9TFgcza0b7yeT3/re3GXOb45T
BSsNsTxkG79oxfC51rE4ACT4lZB8qzoex8oZEBj+RZSgyiLLSSnlzGpCiu+a6iIqsGw+w/2T2EYW
L0gzwmZyFGZma9ieTMriAbCgYTRdwG8R4uwzkj+/yntf8kQ8lxJXUwW+wsQvKIKKiAp718WI6nie
ust/s58RvcyksUPoq3N0PdsvLot5sWGhX63kkIIcEQqAjHHL+9kU39ui1vbKz8jwBQ4JeB2PHCCb
i1tjMQ63VpcDM80FzWzd971z7soxczx3Wadwp83E79HrA/Oc0h1ePMAfq0NBkLRzCCYCdKGK/aI7
UJ2pS7Q2erTxryRp09xtHz4B8HlrsvZeISFl2+bMH9AcgbeR/WeKg5w4Fz84F/tbMwjB0UdFSf7T
IR9cKcNKqblrwH69OYbI+bhuBrREwSeOvJUw9ocF5CxiGySABMVXo1i0cQgJXdUjG0rEcpaexU/w
78JWwmCnv1FMkgFTCIgPFjvoNed84BfdGHXwaSTjTjZ363DhPRSt750bhqXavaVRHce48c4OMEDu
0Nhl5Ng/0gYqR/L/J6WISckigizR1HJEkiAHsRK0WEwNYp4oZOxmiXdPjfNjKRKGczcNGf/NfHXj
hpyujU9hHdDEhIGkkK2OGvioL7rOgcwH/HdhMkwZmsHFZ7s+S8h2dfraHKTFJl73CLbAnqfr+SBG
7UdvozxF8RM+ElxYEu017hNSvuAwHw1pPwQTBcNXINhzcksH+ivhb0bq/X3zGE16scDTwBc5gb/v
P2kTXEJNAvF/ovs3/55+xtvpjm3rNVy7hLWEU88Ch51FjRc89+ZPkUjvlzarfj6E0kXQc1hQDuWh
u2i92k6phAQ6kRh9kMM6rjClyhg1qrjzxLqbFIeQUwlqEZz1DClX5hjI9SVSP/5oYHzvcn3z8jkX
BIrStjcB4h9oLYSoCoj4JGxGakyDPfgmDdWH7+SdwlglRboaEAUvQAxSEjKlXrhQbrF5C2hr5zPH
nCB2EPHsWDre3AHoskhxFf1aBWWhBSpz6ctaL8EYTzPe2JOMkjk6CJt2grRu6GILR4beXD59KxxF
GDDD1ORSMyf2pcsj0P1g+ez/nGYYbqNLbvcoWGftaAWNU3VpRgvr5hT2rnm02fwqg58EQ1BhKMgl
/+NogvVI+kbVq7YC/tFvVrG+DD/XHm9fhE3niEHJuWGuVdEyJ+VKxUQl3568jb5jaQmOaWgyyotr
oD2WLutRDQOnooKr4fTq1iDLPtmvAx699PjyYayn5uCDGstncEWUGZrnSiBhCN5bsqiyDGLo+Jpk
2EgRWh+3YuM0xXlo9djY0eUM5/52iLmaG+uuuQ3MNEVrDd5WAQDNyEU2ctPcH2wQB6G03EJB002k
L5ODUL4vykT7A7bhWvrgLT1k2OW+GPbymAHn45/S8/byAv5sM/P7E4S1V4oXMsb3WCJU2Blv6Gzu
rZSFUTbE0TAaUsu/nR62eSD09L7N0qbIWp4MU3dtGMPo62CSXK9GRHZFx9bQMiGe2LjroJu9HLpR
IIBLW0o5ysg8l3W4VNyfe+MoLf1OxqEPd6EsLN/guEEhMpMMlLIc3ZmuTyKCZzUwV9r5Lxf5f+L5
z3GaIl5XrCBG5koGetg31sPUAHykIN/jfD+V1+CVlt3OaOXoM+J915YW4SMQbMxOKXwPyUKYn8iD
CDssTTfrBF42M52rpKqOChVhts3E9Zz7HaPl92p4tuAmDy4ZxXkeKu9Puc2RwKIxhVbn8w2rBy6g
aj7IsOOjRsyazkZHpF4b9vK4zAO1yfhI6PqvitsFU0I9WJLhHnU42Kpxpecu9wJSEsnGLJJtu50E
x3cElYNil2zrNov7POKM+0T3qJoo05gnuTatV/NqSp1VdjF7YcIA/t5FveLEr5Jso8/MYAKanpl4
zBPImSTOQEXZz/4gbaaDcYwYTa7bgIYO4vmni7jiImxYljyhHFHJ0/tbiDHfAxY1x+J8f+n4p4E4
fIlAe4STnWaIrqet5+idu+WHTlm3ecDrJx1aHkoMNXv3rOAd5DXv4845/JSdQgApOiG44jDogxcl
5/n/5r5RUbUQmepS+FrA3odllGiqNuR33LNk1gDVfb/W3Y+jgtWWvUylvIf4F0wS0IyWziuv9Kkc
l+9XrtY2NieSMVRU8OxZzDbIU+L78c+HDXsVJIuGfQT8AKaUvGDArIK5AKjLLV0hlQLkFw8/NNnZ
Db6sAwBgwqPbwqhPGShSjqukZLNyHjILIywx9D9PgYUs81I8EAVjYrphtvboKXH86jewoMLdfHgk
UU9z/LWBAvL3p+pa31aA1gXVQrt2z3IyTeBgIyMmKUTKux/q6POaUFPODuDJMJ/99V4GIZlvaRYt
Bg7QJt7AYBSTeA83ScoiBtUeJ7sRHr1kUJVqaLcA5yy7OeTnjzbkNKhTSYcWY6MxKHf6gWZekgVZ
xrQxkYt9XRe0VFYKKDxfYaOfmqA/nC2DyFC6+J8csKGXdETnH/nLIj5ksiT9l5O9sMOxV20TxknP
/sEoGOipoCmYZtbzV61s4JfbHQgqu0s4w2fsasdg0D5JJD8yRLn1D6odGwDE4upj8QNMGpnuGazt
7H3IEPnXxY98uq9zoDdaSIAEsYFn4codX0xFyRyXf/JHS2CVPFHwxAjOeE38dcOjg0j7PzYOegq/
nCVlzpiomdpnT3vfg4PiFDoTJn0MLhCweBLCO31fDFqMPlY6u1BdYmSD9NquANFKbJqDWf5fX/ZN
IyXNVJQ78YbN1qfb5cf9zOIuEnEPR/NzWDg74FCOwsLeMDp2j1Yu1rfY02tHAaMWoga+tMgBDDV5
3yDgK5SLKOVGsihIZVy0alwXLyPBDcD0qolP9PCdEBV5YVbTk27GWQBeiPZygnEiA6il65QXta6E
kS0FQNlLZXVEHBhjD2KrQkmZ+vij8YLbwGgclRJNr7Gi6gCzaHmnu27UxETs85OUYKCRbcBEr7gJ
hB8jSzZbkV2Cadvbb2ClNxlXxqgjka/RVh48CPMyYAVOA/lhOjNNhrC2eyfOUjduj+UlJJGxyfig
TfjF5NSy7iBbA//C5fjtI0WTf/nHoZLUHZbdMdeoVqWbUbYz+ljAHCXJCA7qdh+ROmeWN5dCnIa0
AdZtL9QMCD58+RhAAR6yciWUrAwiEjpLP/Zz4ErUvCT+zinrExkgVJb4PCd38xv0djCDOzO7O5Mk
wo+u/IHY1j0P802pltvIq/JPCcHcJHEzzNx/9JTIDji8nzhleIK1FUaPNd06ElkyWmBMWJAsr79N
q6h1bVgMl5dhoV3ySHJiezFKcTYq7Rtfho7ss7TyZfKK4n3lpu/nsCe7LlBmgya4KVGX14xZwWu9
yai1+tPfQy2StG6AjClo256Lt0QbyzxnEHfrFnceC+rhrSGkPjgugwmlGiZtFzgHnVluE9AMT/cM
NhI/EmfQFieKwrStwk+0QuFay+La2Cvkia671VFoqzwVlnWeFOVIOozbiVcyfJ+lW22ve0F30C8+
TzBKV41JIp7J6uvJkRL7G5Di0yOTO9pCDd/QHKw+Tqkz+QBNjw5QX8CLRkWWh2etJDv28o918LrV
2OanKYBz+3MdRHw/CGTYZy2MCdXCiJMmWfxUo8zsw380rc8NXL7kMn09ODGx27UUrJCYAys9qQXk
3nj6ZuEeS5UZI+yUvJxVwutdJZiewk2ORc2zhQdn+I7JthOD6O6yOicLpnfCDBg+LLrU3QnOax+s
h/D9R2A+aIVwcY1t4GSU5wc9iGOiWmj5GEQSkmyDsqt3uBl6QWwCQnMSUW30FmYoOiFdEHzMx7uw
Dr54noMG72IJR/sYzwWfbYrIIE5ltSPWoUuL1a3UHhwg/aDlvwdN89WvMnPG4PclzVFdyPKlRZVk
LUKbSAUgCrtyVX488xqFaxQdGihJs0ezdwsm3N2+9No7icZaNhEEZ5Pz5bLW88PsG+/UGQue2Wye
+pBISrIqDCJh8jMVlTjGVCfVwIrrB/Zq+Sap17KJ00beMBDMzKbU5g5fnW2z7DWp43/D49mKq2Tk
1u5mNuTElHevtIB23JphP0+z2plmIJf3/qJGS7mBzvccb2Y2ptDhS5ozitbobQwJSc4sX1Gg0fig
H4qTwi33F5W7q5nNg2iGaa0/db41Newhg5EyXVVvig7P3HAaGF9corgWf+zhSKkxF/MUfIgZ2iM6
42ZsyG/0/gw41yXJZJny/Vzm7jo8zUZtFkCwVU05aRZYoNkXOi+UKJI5Rrp7/HKyBLu2A97jjKt6
py2Z+Kr5FuPSRe8os3aEhlasHzjivRAaR1ehCsusn3KQYIMlOamQtx1cYuvaKd9Allm43wBRXpjQ
Xs7ClHr+rdmngJLCzZoRYxUGfDOyHYSpIhMhZoiN7RQrij7+y7F/tWKAlpHmx+Bdx/wg2+13CkJP
8crcrp1VViULo6sgjQl9Bv/YWuDGQmoTxA/ZxRs5QVB9T8OO2bDwP1pAdl2qmVTlvmoHiUBZk9YA
KiR98YSa+z2w8iyZVCelLj4LRbrz0KSnqwe1++/wMsCF8PcV41NyypNCpd0E2pkSBODmaLvWqDVs
xhK8XGicPkVPaoTGhBUdEcmzUbe4Hfea5DuWMf/rPFL4wWoqkSulkfZKlhADry/nXv61yBbArOoJ
tbORXng0qyEd1KbA5GgopKvxRENUzlklc7p3A3EpUdkyhjAPykcN8YaV2rPIctJwvFhvP5Fey3Fz
IimnSr+mQJ8S31w6u0XHlIk5FWVHq5cwZUP1MffcjNqPAAiPg939q4o7rauAynBEyz05jMijNt4l
L/hyfajvv3ifSe1cbIdeMYBJf1+b01HPPYBIMXjjLI44/6xzetXq9rIm3bVd/b9wnTNME0iGxP/t
JqelRQe9YGgKJIk1jtKBUVxG7dSaojJgUPrsE+5/cchJcN7TwuaZWktI1GtmVjifqdJf+qGoOfcG
bjhEzo+DlTYCVVPE28tBxKtmS0l0+DTdGxvneMU7RsIZTvOhaXOzffvU29iOE7Xac6rock0qHnL1
41HFzohmvNPhb0IJsDCZJmmOJWp/grzJFCiQbESSCRoTpbQH8ZK46z9ZgyZcH/VOwSXLnbVRqsKW
VaN0IZD/e13GMuz1VTg0ChcuO2S9LYN3OqmhIBMGEmuav7vw2Hy4KINPlNfaag7S8Auu2J2BGNRy
ZmKHCuLdxYQB2vQBWJ8YMUilCE4PQWDHYdqV7vOrKKqXdG48DbrDn7FX0kp3HnyRLMiK/r5sSP1r
UFg8GI2A48maIMOtMrxe4xL3n53XeM+DtnsNvxd9OjMV5kGv1KxKk+9To5kxjK3cjWtJ4e6x7A9k
OC60g5+ON9p8eOtdbGEquTXFTWsAT9Wtu0s4OLQwqMyKlHDSwvJobJqIZPScr2uaWJNM+vPArq7h
F2nmQOir3gDmHkv2Drf079fH2jlWuOMlbbI3iOxmsXf6/kprmUwf+O6jWeJ+cZHYddDXagmwIm2o
FBhoPED62CC4DUigMmg7sAynkw1z0gU963nGIctNxFf7K5D8u/f4BKfmKfcApuL7PzSYU4lmfLsD
ad65xfXE1X3g6mFQN7fXnIkSNSastxbQ6k8pANnvGV88vDwwukx2hjVSk6n5MvM1VahqXybjij3k
0LdcY1sIffUY853xUB6MWR+mdxpK1DhzA1QB5GQTXv/U2EO43273aoEQXcFiQZVmhwPwFNXHjy3A
mlrlKx6ATRD/MgNLd/vrkBx5hwkZCbMbvJKbvQhT6HCz1uoAKmBKFHNrWs+3sQ7xkiiD0PtkhThM
RbeENrjyYO96LxEBvvWfxgBI9xBSh53YjtdwQ0rZFB768CrqF8oyX9GOyNHrLdq9U87qVWKJfxwN
6n1daoF8dTtJJI1v+cVmllJWrAFxvMu+hIpenDuhzveLhzLOb+k8UEDWmPzTs4htU+eYpvqRVS1p
EM1hNYMaAGfmpu1r1TUB7Cmsb1TeIBPJ8cu4QkpGWhFtgbPN+MhnSBHnh6avH6PpK8Vqb4jMVqiu
lCajpStYD0ET5V1yo2OzBHeBnl7fT0qzdXcRucDXyUSWT4XP99L/Grz82NaT9Fo2cpNqyb3t8chD
xoiwXgXSuT4aHqwbu1j7ZNF8k7iYGS1YdlocltAs+gkeJhAed6ozMg1kXqJMMSiC25V8YmYiUG7+
pNw0oHprwhOFHSeSQWQnZhdwVSBFc65Adm5yi0oMvpoJTbnit3y5l9IsS6wcPS0h/n5QvQWLcaY9
HW1s09366E5O5/eaVoxoL00Xo9I2PpuyuMV/h5PyXMmzglfrVKSUPdUFKIGajSpGZjQHuqwcANAP
FAEC37X6FeJzuKCxCrh44FAY2rHp4Ju5cuCa2TrWIybui10ypPT2A5cLskoOTV3PW3ZdCdj3zFDc
uy9RLm13cqW/wsQ7B76JePGxI6S8V+qTytEImE3xfKlaFNYRGR/8Iu+J9f0mhTW5TkoprONgnOJR
ADxDxZkC7i4+FMeErFvcs4Ou7fQiHKBppwcbyrNo8Ig0F4rbxFExCXgMpKa/J4/1axAUkyEX1HwS
nwtGebFhe0OqH8Ofmv4vDY3xl77IwQIxd9i+pDXXsEAEX7158y3NOphf6R4hcxJOLjY381in+PiK
C3EOTFmFixu/XRMcHTveYy8ACqnlyVbwcusnvkbLI+cxETDYzX/x81/NJaCxIi1UYSYRcP8pVoBZ
J6JM9NlOpPnKI9FatgJdwj7U0ZduFtd9BnN/EyOoaBPfIRRYV421UxDys1hSY9QzYtC8PDvmLen2
boyehscUoAFTo1iY+ztCtrUvqsGBJWnkqh/GA72BDRgNkZlU3XvYNKSWLegbvxfdsnxOoxsl8bmV
8QCx2VrbeXusUiC6y8y6KnMb6wQkDoEndAJt2oS5etjUJ4V4kJHV/8KdXEGKNno/JfRfAFt/6e1n
s4lKnIo+u+OYM/gMob2n7C1o7NTZ/KDjtczI+Q2X3HttnwKr9vfVkveQrnhITpkwKi9XtJDn2hqC
30iDuibVgswTqkW44f3OxxGPF/FlVpsmxH6g3wm+rQ5uiCHMdYNMdNrFHGfRrcHF6Y/6E8DHWS3U
wUAuBkYmMsBFzPxU3+wL3m/ACGwCPD88q7YiiE6ocM6OG1LRQfgzuZsLYxCWqbMV3scR2pwwzbGA
z00RguM/CkQb4jpy0upWrmnncPVEdWuAREDOBAWJ4xPAGUKGpGxernrl2bjlvX2NMf2uTGSkAZBK
a58vc2Htlz5RatLQvI6Ik+6B8qATLHM6//gmg59zJ65+HuK9bDznuCxf6NSaO+sTWWBusWrGNNAD
bicap1GjclSVXQFswHUxQnieUfF8Ul2dHe2qt2SEY5qI0OT6hR31wrbdYJdvi+k7NU52Wok/Prcz
lFyIDhIEYkNXmKdDijigmL2FE4LM384WF5+xZO5g8xFiKiOK94pXPLwP619Nd3mra4P661+VGtuD
4Ly7+m7QKRrvQQyY84j4MUONXaUlOIFjJEC2ED7H1VjG6Y4iCwCrs9Ts+h9XGZiAZyYhrfiVPiKQ
AbFAXDx9bOrCSu74jkiKRRKrw9JL/x00eZR14KANAsetOa2mHLegtbl7rmxURttqj4l9iVx2D8lY
Prk/KwZVzYumhqCa+uy0t9iJZTmHe1khgChD++5jkXA0SAJ5EDOMD17lQtapafNh+YDDiafo46ll
tJi0jSvn6gTSu9pu7XiQsaBLeAnjMHiG0zAWGPs3OnyEv0Cb8L31EcBMsfVJw9TQ7F+7Jlq1mCqR
Bf40FgwOy1WQqwBJQkg0Zio/o7pQtCmYNgUa6tMBK8I/++IIm8zea04hdRWhuow2xAgmIM30MNuv
sTB8n1L7Z30G5ZvYWN9HBsOD8l8NQGJvYSOD23fe5LS3i7IKkv8jIhafy7azK24MB9V+dlLWrALB
xYiZmp0a+HRRfYDpHNSPnfj/MqJeMLIX8yPiNPOUYOfYEbc8Y0oxH0z3q5TbY6tH18G6VXP+5pDI
ioZ337dKbOq5W71TlKDRtHDDUfqRceTOVqF1VAT4v6GYvnw/qYnDLuesWbFIhmvRKk8T3eYUZYVG
nJ430BfPxVslcWTHXkY/cYy4pL+cgXd4fuUfq3kanjgmgSl+aTSeJ3l6kXc2CPDgYn8O+BfOdYxq
cKnUU2BDfLm5GZp05K/EdiNPThHdkp+wUv8TkD6NL7wqyl8zb2BSQrffmaHnBHmrK7WqluyXhvLr
m5FtTBkZarQyIpJLiGQIBh6AfOij+Pa9gKyjoJIJQdLcI3nKDNTxcQKEwyDmPFV6XKM6Hdl8uy0O
UIxG2MkGeCCpqEpN5hteqc8+S/+KpLlL50aOPMUdDjeTP5rRcm/xi2OmI2EsT3d2Ke8IUmcJ+d3A
poe0FT1pygRR1faNchGaUkGo4etFrSlGEo1tVkXExZMS85NPxISs4ckFRUTsh9TY8XUYz6IpVFGK
Q/vtCe5XMWi4kzDsice/Xpaukc1IRmsQPF86IXE1mP3M3MBhZlbF4s8FTTncG9R9MNR06gmWphq/
isy/HSTOqjvAv/Uq76enUS9qLB3tsfVb9uXuytleCWHsW8nB+sZBoGvUDxPA3RZ4JJnez1izogLc
QOmrtGvhExNN8XUntMn83NOH9XYRxuyEupajMlzcT6qiFAfbY45mTAkZ0kVJW6LmGAAybKhUuLcX
yagCEdjFUjriwDclanmw/a11pX8KkmGTTz3d3NODlqU03eKWthCH99MrtRrPj5+KOpHVJXsJaBzv
5nje3L987bO+GcNGl1ahVzUwqElxiRWRBgv7ThK6CnyDLdXxu27yY9DMjiuGMABUhLSfi1uNcG1h
H+ezC/ImUGP4cAZpTqLpUciEvdN+zrPzutucQSVMOGeSfN5z9Cf/0O18L0V9F58KU2VN9nmxygcz
kqhKUwJbTAZA890yat7WLft2jzWpYEeNyeY5DK4GwGxhncv5Tg049eXVY+lXMpHosv0m9tv0tWao
4gukKIC5FS1W5oVgYGtMaSwh7qH6L+OLpzREZVl0TWg6oSV94Dx78q0JMOmVaDftF7SkRXeevNNA
WwFyBKjlB02cr3qM17k5hZ4ONPY4sFSxnP0P3Jm95Jc3aOjjQpJJ8TaMVOH1wSfbyRrqCriSmq6R
LJE4nyzys+kkYHf9Xkqpm/0M1xKsxx8nMHlwjgspVyxPqIARm2qMYNTvLw1dUSF5DIjEUIiL++2Q
ZkyqAq+q/9fFl4vuuP9GxeJEYKbHRmDsJzR6KR1cSlque99GNAeLIJe9qY/lyzIRzWGTGsZlfnYy
TUn9OY2mnVJ40ExIM/wKG+JClBGO+OhW5roC+7CrJXqkwdeyF4PuFeMDWsDCCL2qlg2o1a/jPFfa
wHnVuefIi+GVqq1pXNe36zzOXnCIBZ4p9G3A3rHLp6Q8EGCyal71zPm+7XXcc7LMG4Stw79sJrfe
31bnz3G8jr7JGLGkt7NEuBqXxijLl0407nfvFjcXwgQk8hibFSzxeZJh3GMJE1XmCH6CmGFgp9eq
XZ51db4ztFDggYAIHQhwWYO9TgcQfq61hfieL4A8yh3PGjVlyqi/+0j/RVxxD/NXv8guutjJaf26
Aw0a/E4FQo/0kGtv6CqbdW8EjxNuyuWStJRqXT6bQXOdRJ2de1ICvOm7YDgCSSiNdSIfJ3MBC6Eq
KEqse11sy/1hUS6MHDUbtr/UdOwXhlHF7kEOOeOo33VL1Ct1IdAuWhe2ROI/og5sDyb64F46KTs4
WFB6y+YsfEqS2OnKyMII+4fMniXUpMSy0iZFOBAVJ46FOpOWXTzosrceRaUk4kLl9COkpA8KiYGc
ansuCreyBDFh0QZJqi1eFirUN4L6vgYTT25WzQ0cIy/J4PnbRfzAZRQ1/jISVdJF8zs5fiLUDlBk
+3YfL59HfCkCPzRw+LNf5QINAfEfSMds1aUvipUb4dz3TSTvtzRC2b9amQCPNKl72c8x8bg269D7
USdDKESfK7DS5ij5GzxB9PyjTesfIBv6OOqO0ZWcC/JdNrCeR5CgLMAeQrax1aaGXt/5iVQGZ5es
F0HVsNRTuch9Ym3snayxCfow8j6NirAba5+doWM0Rg0ZpxstuN8guIoZXg0fpxpulS3Gpqon9EAa
CLwIABtaV55YDOYKlzJP1zVEPOOz3TgDmY/3IRZmPPutdNQxVG6RvGCmlvR21dST/5suL+UoYqMo
nQNJTnaDQE32BQVv/6ZQqyio6Pc4k3/2XuZxSHz+qxkYOT+PgvLs8zZAtZKud4V6EiG69ZSx4mzH
Eqjt2sG3IdNW1G1Xpz4goUwQvJawnNB5GScU+s6iJoNcTf625djcg3j0mY0IAlhxA9fYvdYnWnSg
uojJblVajGzGzDL+2xdrC/FeEIS4wSy1nPMlV/+5MZaEholGU2IcLMkAhL1nzlCq6wncMNGlEXcd
JJiq1Rrb3TnpgSpy6m04cWXE8X9H+kXhrVZjDgyViP62JQrz/gbOuTMfU0ZWIHHTwISkCGq23c8s
GrePgstyrWV6L9yPRTT4H/xrENRGntWrMpKsO2y+lMOQvM9BoquYRozNjWeKjBSH1UJMU4e/OMfw
qIbzXDgVEaJgtKEypwPI8BAvuw9nPaBim0OuMkXnKXbELpsZ8CXGFzP2caHmGqZNaPtiaBJIvlRm
R3uOUZfCDKCuWXK6JScynzRoAtrdRNA6QmNO+R0Qzh0ynfh3J57TyIG8u9phcZ/maKjB6yFx4Kye
jkANI2/asavAKdmVHj7VenIRtaAyZP7GGq+e7CRvsdeW500s1MTmDw6MITSmWMXF3xv7RI0Z4qcX
Jk46gJ3fyN3ppTLt3O9nsRVmS2YWlEPITCBuexteB/dAyvEgdyrOyHDjAlh6YxTZ5vuIwd+8edr6
hmWTSIWMoKPh8eYeZ+3UFfKf7zCzmUoesm0DVftQ9E+WCey0seQ1T16wDunYkzzFO9EITy1s2d2B
bg4lL7zel1ygHQBnteRWRiiVUvz+WdLOue1YZfMQouHs7z8pd+IO/CrHYvb9TcboC4vN5vr/YIbe
reko6aDMXYLWfO0e1PuZmFntAApjh9xh9ST3kpI57RDsFjkzurutdH0BlUzinCj/lFLyn3TRdEEh
HylnMFTbPU+6HMi5UOY2Z5aaD0sqPQLjoawWU1wkcVaPuwT5HqOSltkh1m85+XUl4fAGdM/TdPje
n/rYE9YdElZQnFo8Mel2P/1VjxseGj4EElgKk6iU3C31KdYejqXOxlryN9JMGQPfaCf38Gj0Ras2
lmO75GU3Y7vv8Ugf9pWYD3OKx871zaw0KFPgAuV1NtLQI+XyAPRtmcbFUnul1a7jRCqsGqQd8U1G
NguU6YttKAH0PNblEeyDU5M087MiJ2cKBAVURhoJZpn/US7ok1Bmhb0dpbrsVgwkYgsqIZXEi9Cf
Ew8KqV4YkuCnS6/TlHi+dKDVmdqxKmHRyqLzjgT7/eJ8j2UKxoCbElnabngZkVSfo1FDwqoHyUwu
3bePjydx/+La676fmapOemb1d3oQznfwMzz5zfgynAwGN/OiM752a7LsFPABPHxoSluLCcN7JMI9
YROANs1/YYtLf3b33ScSmE183ZPFpqC1TqXmoCkJUWikaTFo0ZyfNmAUhWSoaAis1Fa93DBtEreJ
x8u6dSSwGa/nT9Qk6YoJtSWjHtq9rjjC1wCXzy81L4ADksudGyrYyqBvTcx2lbvFgMosTEhrux/O
SJfRPc+A+zkRm6q2enzM0r1ZI+0XUN2FfpDiocnjeeKXYG4ueguunOuoQQfGCfIz9n/iaN9gsbCW
aXOYrQ1CkjxyOvNn90FGmoHsIxpiNg4PRCmuOvD8oDoSmYvzVrj9yRMLOYY8igMM18t6RaCWxO9l
qbAeqkTSP7HnUZmzzSzmBoKV9bcJat5Olv6UtnJ8eO/t+DP2WDYloJtAvxGGBvEKCGn8tD9UWU3/
0ssh/xG2Ia0pzGb4imnN2YdgKcfKvoGcTZ/ZHx58S/6MgAZ51qVYkfCBQ7rwkGzko+VLkIpYPgMZ
zRKhw8JeX7K0dfkRZd8dnu0DwF55+DXfIgY0hNndbur52xcSH/sF2xQe55AChrabA+5ehbOF5Y+w
tLVyQHuyj9kZ5eRxfgH2h9k+9/Z9FGk71kAL6FZXZG0VHnAsflBsWF7Kkm2TOjM7zgsziONbv+j5
gBXwGfhDFQRbGSytxLO+FpSnLLczoG6HshaFM9HGOW75XFLXkhpxie8DifwbgsCzZQdJ0cKGHOb3
sv99/u6A8rlaySSYJdY7rUeRh+RkSbI3NiQpWZX+HfTWn+2ObH3xFyehP9yOBxUb2W9XGw2XwzJG
uGWrRcJio/ZOY26KsCjDS/yBBlHwBzDkrPjUYyWVknh8giScG+GfB9vbiEmYfjgrd5P2/pyZGHte
Zgv9yY1NJGl3KRn9mk9v6tfqf+CPnRiiZ2iBRdbQ95iNlLZi9YUYglqA8TIMDZeg2pJjqsZ+TlXJ
HAKTGsmLnYvfI46HVcwj56lEJ4BmlRjCRN9TeWZ3Yn/3MrCyeD1jdHSZx44vBq/mNRC+e8rTg28E
nXtClD4gdEe7tPM7FisKqxaNcfe631NYI5+gFU0gvePXxEAyZ+3UWplW3sTvuympG75wDgWbVt/A
O0rd06cuav4V1ryHVF8S2BxcCjtupJS5uJ/KoeJrBGwDHCFLzmX4UBujeoVb/fCEFxnNkhl14GqT
Tkr8Duc1aYFNCE+VpPF/SqxXcbfGh7EsHv8ENdKteXGSZj7XIoQ+MMUle0xPD5q09u8MFQ8zWoLI
y3McWvwjt0bvxSdsdQRLuBD7y+yyIXg6gBbZV2EGyz1UPxu55hdXdpvZ36sTSb0icF/5iguAyzqs
OwfmRJdmubH0HnhcjasFD4fI9yOFACN1dZnpfGiD6CXYO6+iGgwbpXWuCu+s2R6i7Cp/z0XERsBF
uk93d/OjpuSVK5j2AZTq86/0IxX8n1kq4Shq/BSXvAoJ2FBZame+M348fg8jeq6ZcgdIvHw2B5jm
2zriqX7WFLP+r+zGluuA0E99olE4dWVVStpGjYMazFaDMmsmc5TfD7acuP7KLz51Bw97nKUYG+Xu
/oKqXk19TAXWCrgamw31utlf0SiBxvjLL5+WTy5LiwikXobzPptN9pMyogi6otiLZevqzW1XaRZX
eSbXsh4ACSvPXZkmaCEVO54ch9bPnaXV5wo2zpzUxY9RhQaPzBuvwujGx1rfII8kudqT9vINUwSR
Fblxeg5/1jYGY3PXQFjI9z+qpInQPkr84pwsqmx8rp5aKoZQK689sIodzBsiJ8fFhNS269seZqlu
ozjlaY3g9I+3gNXoEh8XAxAUssxBacgt0gsWnB+g6Aulywewkh1tLu3BehXM/8UVgD3RivRvNy6P
hNhJKJJgbkQ+/GEBhscQafyNSutY2juHjcn3PkmCjRyDOY/+zGKhP5GaLd2kRcEpaVD0pM7YmKnE
ksKusQdtsBk3rt5uvelqRwpEwROixmwDGdJc8Pjst7cRYJldtKtM6QRk5WGPO2cEjRdUvjMPrkXV
30V+huRsh0ihu11SO7VH0WKUkyryfLok4gKysYJaMypL11IoEVAn7rIU97OTMhNqnAu4/O9wIVtB
VoddbRDtGYRVyEn88Dhkxbbl7aQ5rGL9Yx6gtS7qSeFbNz62ezEZm9YHu9hW82BOHGVOSFbMxepV
oWE7yOWZhNIPB8EZg4nLsSUQw5+v2nU3KUyZI0arXIra95l4LUjEmj7piTm6q6L9DAtREYg0P8sD
l4TbQw+les3OhZeL8YE/s1f+v5J6quyhBI49xN4WEYiALo3w4bh/R5VB0Blk4QxCsPkaodGzdiWL
0TWKW2fa5phbKnElD1N40uKUmpVitXtn4/zXfd3rZggRLZv+g6DWpt/2iv+S43GhtF6PoNrj3EHH
7NyvmVsTbJrg3ckqbQd5kCBVR1qS85fifEZ4lJQd/LmzeM3FDo64CNPs1Is1TQ52hnlLOMSbX00E
pfJsIheKliPFUrP0S33tTxNjTEf6z+K5ukg+t8KEC4t9LR1eyM0t9nl5eB8JJ8GtxExamFBRZYyO
SR4CmrBFYt9jMUz+FWqut03kSo+v0N8C9yRcSJmyjUVIGGZyqj2J9H2LQ/PkS91tgh5+x7Y2+Otv
wi3pFIPeNd7dE9VHpLoFL3/AS31DkkM+UewNEDxfBxw1eZ+SkbLpp5PvTRm8wg3taYr3g7VqAt+3
b9/0MRBLfBEUy82FIojLZEcGKvaUgdgCzDdwQXsUJaRz0e28MOzqM+54AuTIuTStagR4Z89FAtUH
z5no3Iy+P/ecjZPKrplt1yYtoMiZ5/C2xQFOWQRk58TriekVcz9tkl3xSvsqIJZKPRCWOVxuIGEG
+Q8SnuGH2quMDjL7t1uUhXYCobXaIvz6klxecmwrYig7nG1EuIGkKYZ3OItzcBdfnoUfpx6jNuZf
zKIiZW+kjQ5GFhg8XeXd0gEEehFpSM3nzFizkXzgTy7GIIcG4QycVAkiHRFQ/npMlYO1SgrxLcYr
LRwa4xdWOjfwdkRwziVKBndTynbn2BoyWR5JEFT4QyPXMsgL+eYNHUGpUN8q8o9fcPaXSyuS6UQz
5RJEJWeFr9+A8KldQLiP8u+mNG7KrepVXiHnHAjQFOpFtfsUYvvXaLatbricbTG3ii647OqJbp5C
XLFcGNYsFRN5MNzfFRWYlZXUkXajYVgmJ4L+oC8wwUJLIOwCTW0hu3PWNYSbf49Dll83oYc3aFGK
YO8NXj3SY/XxhEHRDTecrVoPhhD9BJg8k9XXdMbVecX6PfGuW6EiKaaUOIkIqm7vkM8oWuQZOH8c
CPPXfykBVu/e6tGOllYgPXRq85GSApTFgLgB41JUCQSAVbMHXcck+AoCPxWvYFcxdIdFMHeYpoIn
VvWPZ82xGosh88qm8FavxtSN035GEytQ8F0tpBPsoASGPrt3wjRk6xYOEjyfyQXGUvHGW+w9AVjS
wTyc/EoaFT47E6NcED2rME2MfoGX/9IfTUj2ONHYMnf+vGlL0EF9G4Zg2JuoklDiXdp/OM5dUBzX
TS9nI8/Xrbk9r/v6YzMDHzLnojhsETPv2mMlwVMUDvocb5dQUfD70lQHEP/OAXFyVsSfX449vXB7
SW2c5vYeyllFmhHYPt6O7lyGhgkA2YYP88+YDwU2yfcguM9zSplLJlsaVqUsnsHQyYrRLegVL0Nr
louo1Wy+Gqb1mywpVi9czS1vNFCnwDXdQXCccH/5G2/ryMgHWDed7ypTEZr1unzWX0UAXfHVAs3c
uM5RGZ7WD5hvD8HiRrUXn+aUd2tSsUwqy2DaPK8ZljHhcBZ4dLTM2NvC/gp02DK13AJyfOuPxZv+
uanw2bJJzYd44ieq6IOQIGHq4YtnM5rcotDv3hyHT2vd1h5tYtLXg2BNTaqJEv9yYt1D1RC0zRm9
eyPvJDtC53vGgCSD5TLqLyEo9jMzWWlpewWfs6AwXGNXEBTRMJfAvR5NNgjD/LIF5Mf6WtIYW3Ek
vFAK3+tSM4nATRN8uPFRwnPjm46tUFAjDA/IPyXPrxaSfMKJbcdAEl47jqHZXhrRaL/gBkEpdp+X
G/lXBzDk/5TeVdjewweJNqKoC8+fdwSlbFXVJskuqTRRwbu1CPWJcPjrODYQyAKBjfTSAfRiOdZU
D39LglPHbgil7eOf9lz4d7ig9GYmvkG1knd7We1tKGu0M12kmYLZ5fR0uQB+w2YLEInyoeGd+s5b
hOO4lPrv8B/sgOTpar3xO/8UoD49sKbLMUMX2DQHclVjBkyNoRxoPmII1FPBk3Rd/0bhacMwJBby
E3WtaPn+qOuRaTB6rKR1BWrnvRxN96DgrCc+g15MhLX0NWDqN6oOb9YBaiGgcfGzW34DE0x+cG2u
rTSj5OeD6p9imC4ELzobn2kd8mblMbKgSx6Js1OselEYZdtZP4veUWrXM/X7UuWUzD8OwzIDHjjG
yAC52honvzu3GKr8mZMFHAJ0boyStZmQeK9gyzkXf8vvFIx0BiIVN0iAYRLn6XEckbYP5KWa0vU7
VLKSOnVXzd71aDk0GayDZymCjdtE2g6jrw1VFz5rIUpmfjEeFsNyt5/C6N/6nBPb6uXTEOILasp7
BBiL9Yv8lCT5C26lb0hP8ndP8ozL+JdT65xpBGTanW5cm9MmACl730djY4+sWHyrWNmvHi53UKc+
0Jp6TefKSJNqrP/mtC5ehvwMIi3Vh3cFRwqt8ier8zQPlNB+LNeP6E3FZ62PvBnyFeHzQO7du4kd
Y3Ggc+mzaVgGqJNzPrBRhUjyOfNosCWALdIyzpSq7WNWWd1HGyVdU5O+yueEflPaXKty+of3cR/M
s80IS07nHHEVpXMS5/E9Uw4OybR9QEXdHNGMGhU4gkfuutX1z4VKK71m521Yy29/wouUclVbJ5TF
IWtf2yRILDQL6Oq4YwMMXIqctallp0ICp6ff/kLi0n/wudNns1PvJRW3qhvQiH6cJtuws/SbUnws
bhIFuchSMVokkeDjZsPSAmBWnLEVQ7j34R7ahy6oxfheIBEcPSW8rZEW/atouYRJ1h3f+zR+FtCy
hv4YAUZsR2m5kn3u+jLDf4xFmMcUPUmEStsTNNKMwArxUfditC4ewyJIiYKfzSrRQY+mmyNcY7gX
cJrxcUj+a1g3DAQZzcOONcjWwywrcsXXTATXhV3PFW2XU+yL/sXX/2D+FPhLsj6cjeiz0IxBaaVh
1O5tONKu6Go7TilEiBX74+cnewAKhRDnK4lodlL960DvLgRWQ/COBJjM/RNrPZ50Y2McgDiOJLSk
dnfKQueK4SQdMEH8hsGKfRCvFD/1S8PNsBJKGmMK8B+LA/Qi4NNyjJROYxvLLfLDLY6RssBKCeSW
/X502qqH+6+MNcuIHKTHoSG6JRF6WFRY2e2RMowGlt2m+bVtyUsq4mTlrBZINsIQei8oHqDdMtVE
sQGSp+xaTVl1AtiJKzSZGoSWEiwOk0Lm8vKemyiuuevy+Zxye/Musa0vMb1FmSLGqVyyEAnqToxC
58yLt34REzzDZW2rwadDqz3Q7kwrtO+xmoyriUgpmptbZvMTlcIrgYQFAjPQZRJq4SY+6elhXCGY
Rc3MQh0+1AQocRrPos03ugBFQm/RLEXBo9sThyEFPDLkNBY2POPmFdk7cgXgEexsnojZ8YX61Esx
ZzxMuUTavJNgBx8QwwO7glUmmLJ0dCo7vSywRx3VeX8jK9yx7TZCc6G7bWaAKvzna+fwn+AX1g80
8JGXfFBowlH/qWsxBMsXSIIox4mkS7J+/d+rfPWewwjC43umHBIWFYX5wGbBXYR2BcWbtcqI9vLp
H3w4fpxzbTVKCVv9KqohHWlqX8uHHSShEoLoA1HcuCaIW+5x7zyxW8Ws4ipNnzQJOpM9n8s5iOGh
atnW1sNi75LiuT2QvJk5Dt9Cq5PCKI9ddAAOaMTr9ZcTWHEK8mU3wmr3HvB11KdkVJozOdOuaaXV
lMxdnuazmayEVJVSgawTr9qqDxSoRQuHzsLgLNATD64d31Z2TYk66zP0TP0hRmjME2ZQgNydKq3c
QtYj5dLs6MODXoXKgLUtvuJ6g8PjV1ns60U9TPZm+tuLNde/v0UIwrsm5d9YbGw5l0xguvzc01rj
i82NPgI+NZ2q7TdkkFV1NbNxG2Pkc7/ws4BVwToOst03ByCjDUSvjo5Rf466OU1NAawB/x9fipC5
H904okphhZjfPJvwPlz1bBQwqZqp78p4cL3K9HSkIuA6EICEpYpLe61aYm1zbBuQCoir2tbXeF/3
SEhF1jhTrnx9X3EXW4IYS+gBFb2OrHdsO1q3r1xGmj3koyOJOv7kbNs+qjV6AKSnNc4wcC32h6k0
j1ZhyfZxLDnwqy5816OycVsAmza/criizEB7VgovixLWKNoQEBmu4mOoQMa5vy4GbCb0y1vAg8oj
4cfubrNNRGzs6WiSgbEgkrnSvwl2eWd1XbFn2mxozCWnVowRhu+zHvYLYSzi/QBWfIl0AV5UuJIm
9SN4KuYNccGlSHGQodnMGkME9KfviHvfTct4dOdWXEarFoeBeduUVqChE3mxHQLV7I5eS8s9QYFi
oHIpT15WpbsMuu4pr+HuCRXbhXcfY/LBpU2bdyHr+z25m2KwGhanJMJTXbNfKyQWdiHtpnLGs/wf
LsKNaoCgcDeNjhr2SiBqtkUrdJDpbxbe5M4saSI3kbW+Zjz/WT7/pGEiZURYMo8IPZ5Razv5BPnT
/dqE7sF3o3kx4iOMN7bJBYSBt5ZpBuUJtVv4WdLPbifqgIba1v/1SwkLLJUONdV26Z4r/4B5zGYb
0nJDOLt9Z6fTXjwZl3tab2H5RsJGOfbNrBoxNX2m/ZXZVoHglnkdZJVFElBRjXRpM7J99TKjVbCn
3KomqT7Mr0ewyZ4G8gDATc8ClFsjSUqZ7HjBmp/TtrQWRuc3aEz2s+dxUUJS299fnOwiDU3sul8y
yKkjAzJqj3jsxmLg1bW8PTdbzymFN3PasIYwkSYfA3UDYzKqfmCTO/jXmtHclWQnPRCBesen1DS8
b3Is/jrwjiC82YIzUAlhW6UC1uGy0dZTgjlVEEbS1idSVvGRDNgO2B7kWRiyPEmg3LrMerEmNoIk
snSRBFdZrkHmFRh1iCS6PJP0SX8Fpr3P7SR0xmfdkvrVgvSRrz6P+W9N4QhRXi38ANGSTRbgE4S7
nb7Xo3v259DzFAQUcRzWGLfKEYdbFrwBViRHK4ePk+7K7AVeTBuPap1nbtkUeXhXlwOXLBtbmhAI
sK7+1B+rYnv+aXcz3fL/oKjLXIL6pGwv2PWmYtCJ7mnQ7EYfN1zok2ce2qbo2lcswaXOyXU/uU2O
3D6ityAOge8dOdzFuAsmjc7K31ZE0rjH43Zrmh4I33Rrj7R2vyORWLcqmC42OSztvYwNlEqjryww
VJGeSLnz78ukbD3/Xg0sd4P/WeSkMeikOXi84zDfWxqrDYcrFgtLH7qD4JZLw/CV9cSl5fYRDQxo
Jg3YNK1PCHJGMTahGPOqYXx6f1wRSifbYhoAMSrvB9E4IcUTCLvjWYEV5CS/BfhQaicZYaZqUfnU
cXUKQYHWh+9EW3sy5MYhc86byJvuaVuSrPyc9zSxijB5d1Fc+wB36tguxkJIIb+L20m5XJpSAlRS
IQ/rAfwYachVieUSFvZ9XQOqFsYlOOn2vI4ufK1sgEiAoVgK8Igd2+1tIEMJVwlqodXZSjn7bvRI
btK4/8LIvGnMBcOb+5nHUEFAfSkEF7UisU08IZhXs9ZIknvsDLVy9XJWDMZ00AX4W3fCtoU//OQm
TCQlQLHLKHSlnvlvYaAUE74SE8mNz3WlBb50yKFue6mfX5pS0Ei3yQDQsZB0G15+SWVGD0BN7Sts
yCcheySx0I4wifGELNYYfS/w4L+EyiHvWKUhRsqmiHFNNbGPjia9hYLRUM7W4iZXIKaRfZfGVvln
bEuqftwU45+ijNu91pQzmBuQYxVGg6IFe2iKiBkvOX3cO+iELIOjDr4UU7fdpoM4NqOt7f4bwUv6
MlaKlhmAWqbRWtHUL7Jrdu+nC6jCMOt8JMtGItxf5lJGa/+okLs6sQ79Q9hF/CmvUef0vNGx12ZP
K5NCJVswqmrfQ8rKC+/diKc4tQdEfJbyfYttyWK5iaZEMpeQ6XUAep8dHoOtDSf9bIKw49TC0Wo2
OsHhwFt+DBsvPn7mxXCXsTk+B6l8Gf4vYed0/zWalflHjihgxJytloqM2qHIYgOAoflr2UX05L1A
Dw8hAVWoWkZJp4hm3LoXT0fuiBJb/nInGrWhEgXqWYc+uFGgOq95lrYXtrGhJvWWbuPESjJGam0w
OkO42CbqQXbULRcNoZtcYxzgDHOBGq6Q9OxlvKNrYxdzjkFoVAnoiEFSCmYZVQ+4Jao5IOhKB8eR
1yesnPvPQVaaJCNT+MBjpyTIEswqvHRD0+tVdRLFlzpdD/WgNV/JtMXBPKFoNPtxigCh51VtkHxS
drkJlOZLLZ+9P3E0F+oDnozTVVmpr77V3fnRh1Gsdb4wDSJEAQzOWcU0IamvAFuT8ifgHIeSYDG4
UFBeAmTnNUjS6aWHdUwGJnS0Hk5laxPrpJHz79OEzKVTAo4zNu013B6BRX6R0yOmwU25I3qt0iI3
1EPLGRXEPzRpque4KOdpHVcFfp1DEFfu2pxbSsNUova23qap31JKv9kIjXX/CEx1mv7yqfAbQkB9
fz27Ooc38kEvCMhGHvExUf8naF+m3ZBA8E6ed5IzQ7lrKIjU9IvmBNlHg9PSGDHz57Q7B833AxWk
KIo9hV/CROJ7Lc+hpc20o/TWnEVjVhhB5e6jriKSthtPhpE7UGgeq2i3Hhi3lIVIMxiAArPCdXfg
1krEcbR2jM95wdS9QjlJCAWIoCV12Y2u08C2VJ823KqnQu6YhQJ6IOJ+6iM6YnrKdB8WQ6qZP3MJ
XeZdt1ij1h9IBEt2iqrHk5Yes+Zr4CPkRFQBGhnQajZqKkXlX+RJ0OrmeYTTo8gOBF+ucsO1VHlD
OspSbaYTwIWYKWLJLUewiyOzqqzBpdSsuU6cB5ErOwwK4QIhJVUZ+a/CWnHdUdt6b19MR4f6Kjv5
YHyGzCtU+0s/hRDzvtovK0PHTU966E96Nt4i8RzocXJ4UUXUvRkh3lzmMVSDB1Lk1zpJhtTaop6X
Fis0GbPcB3b16+3A9yQFnYYPWtk/OZ0z3Fv9i1ftjdo3FrnR7B9TXoTc0iMEs35Ib9dQyKtfzRly
Tg2Gw1G3oIrr7faQUVBbAJBQrlN5p9FgiSJVMQ0DKr9gWcDGvGQGYuGuSVThP9jrVBazJgR/DsMW
FMNx07BYxihpu4uxzcjsle3EAIE9FzZ5Yhuiut7s35CdeiWVMae57lHe9xhfjSxDMOEEJruZwov/
Z+JUYzzCauUVyx3NHBa6DWDoLDRuNr0GFkIUYaGkM645FfAZ63cTm/pj+m0/YG5lXY+R919ZL5vq
+9Z7yQO6WbZjHQGee4eB/U1RH0778VYHtNM+HZIF294lk5lkbfIocggBeuTfs+cijupobHgj54RX
2D6AvN430Uk57bBhTlNgA2eeVvY+lyhUCrcx+78GtXQG1S7T4Auoti2FSvnaEmigzB/y1+f4Z3EZ
p3NDVzpeNX1B+vAr8YODskWxJzX53q6qdAIHIBYv7HXqGlg9Is2e0+nxbqlQg4+A2rUWgyKIZ0Ra
Bl5/R/4iHFldNTfSRpVYoUUkxO32e05WkBNWY6UvkmbglaGg5kwR9/uLUByAX3Gmz4zMv787H3gi
e3vPgq/rKcOba10E+2Pg00tF3jdEASc9dgBE6XLsfQ3wp8YqTWZ7eee0gSHUaqYJi60z+d2mjQsB
ctnbgPDJ3S2UmEETKItGm7FdztyBEz9ySAD0Pxt7YLL5oq43gS2cKyIfS7t4kEofuGZYycea6dqH
VrZA3RWDWilLuhzlmo4cMjXb//A6MBY9/Bvc1CfI2ugMeBUbBHPMe1sZsIS9/7rIqO99+jsK25Fi
A2ndq5DMl3YWfFJrPbBujmpzFJ10xPENE6yBf09Al1W2VNhbGpxpsoxV7KmZZn2tLDTVpY66XDEJ
c+SAoI6RmE/O8IGDJ0vmVaDXcRpAIlBrbkYw4zhxUByLMtu6pkkwxVpzVPU6lubCx3qOTWusJcMN
bMoLtCiEn8a2JLzgXTx1hWV6KsSopy3CWb+oA4J+ZLDjllB265H6EvMCbuVbM9OaVsvzuQdL18Lu
aiRHMgRz92yNyIZt3QQjL1JYXUUhOz5vWETFmRQ+VFQP4cz7yD9SSUkzSvgmSfVVYR2fUvCayMVr
pkrDn+9CfKi98atoK+7YVheuYuqUyhk68TBV1JZh6qetgT0RYuYkSucu3QMe4wgZbpsUOADWwURi
RsJurpd5BWdwdtV7SJu2b00wY+3N8QIpaRiZXV4R5k3CKc6ghI8WGbQOcAerMeMJPTaQJzPecpTH
UE1pYYcYHM2RY8Z9BEEUo67AjvpYSMAI3NY2gLtQ+9CrZnVKSM8LstHsxEjl6Re4WyW7lOAVM3sa
6wyVMttTUM/mTvRj9earz9Lz1kswVLXSwOHteLlKWajdnB1A/N+40IyqHpi/EMK1pxUsnXsL2SHs
VSKhrMHg2m6Z+d/12iledemaCXvKnChP4pdKefWNvlkCIjsYJlcdx7l+4/UnUXzHpCwjJaRV/0Yw
NPvu9vrzuiFRyoApn/HfsZkWa2SFFT80jAJiSBD3FVFOSW/j7oE1N3BVmTBcDehG1IeUV25yIZ6n
AsA2ZQHysh1u/LD3e2ZiT5U9n5Pw9ZUhceeRVqseEf7OhPVrreI49NaaxrGYQ0m2bSLTNbxujSQM
wROICGCBtA9jWxDCneUapz384ew2Y7UOxGR7OANlO8Of57D+y6CXBnnxCW2VyeXbh4XWeQ6FcFuJ
5xxSlNYmXszCALA95tpG7jujYy63zk4HvWxaeuUmlx7YhKN/0pezO3zSY+jIXnyubAKWyK92blbD
av7Pz1jCBdE86BirYbI7u0g5hXv6w2agQX1hGHRKN4e+0CJyKNWk0EzjvtemPD7Q5vcSIwCxOfut
d/yokHTU0oDe4w6+kEd6CXB6PJq89xxZjbWr2DT8Ht92mDUWyHIPWYilWajVUm62X1Fry7SMtivi
+7U06nKfQD/4t9aOQrPStxMQbsnb4w1YF8qq0Gn2rYZm9ymAtGNB1wmt53/VgvDg5myNFJC9pzpR
PfbZbVepD0juS8OBwHRY1tF/iA0xsTO6A1aOiOBndYYcjv8Pf/apcUAIlQSh91apEtCvCZ7YjglI
5A2899iknrx9I4xPRt/ErXguG2IYIE8BzD03XobMIhA/cUv7HCy106jQWa1Zhprb6qyh5dFo+CQ4
/BX/Om8UDB2/85BKeyoOK88QrkfpJMK27qJVCBEwBt30koFAOaON3NNbmn2aG25SS/vZl5Lk5QDu
GV2tc1sDdqbu53qHIiEpccBWeMrDY8aFmCB4gOMCFkxfV+Qe/9oxiFTzZBdQeAAHFejFeDslQAae
BRhD7mRer/FBp/jOIQr5GdWtx3GK3V3xI6VBsSY3Ko4ejzJxJYVtme4YHV2s7xO/KT6TzsrlKkZH
rHb2PaolcRXXnW+fGD8RYaOniNvVkbAAXL2qiabIYDef7P50zH3Yo/gA70L2u7scLUC8SLDH1SYb
0SYPT/OEHsgFoUwi9MuaeUa90UW5BasrZElSTJA+GFblLTVen9AnSMDXMtDhKbVil5QOxM+whwdr
225pRwIJvwhdJnl50uuGDcY34E/4fhJ/gakqWAxPblvdviATOaied2xyMSRm8GbpcZyiwnCvs7sZ
A8ZwZ9/x/Qrx+I9P+VuW4H2p+p0IwS5pKNr1YUOUKX2zvujOK42zXOnsO+s8O6AAeFVPJPcFIY9Q
N0lxIpGsXngLRD2VdLLTH5pIUKxMRXF6IOFtjDC9tTMobwZDCeDYpZ1WqJ08Iw/qS3+87/TGkIZZ
RpHPLhuIgeAjyaakAOxyvIcVz+md4/UQCFB/Syk5x8kilgroZQrhswl/5b3lt3rxfjZXcC29rVaO
soyMexXuXhFYydVC65t62wy2RO41BMS2iMg9AuTU74k+uHv/TU+zuZW2yuwGfvz2KutPCzWvNq7H
LPwn8lLqqESvrPD2QEATTU2VsgnHm63MQlDksQWBY0CP+WstV/xggiBrcJiTUNKGu4ZUYfHe+hJy
JrnTqX8PfZfdVTxD1jCHCYXulyORILP2iQFnituDo6iZH6TVwIdkz8T96/LsIHpi1ctANDYFPxoU
OGB2m4fRsOVLDc6AyNm6CllLBGVDCPFRStPDBMoQ2jThA+SF+vsk4FbUHcPGn2FEqBLpOYERJDin
j5oXtStLm8yrpkTv+MIss5MwC1/7htPejayn53fCWt1TMjgrKz+lS3VEHuFOgaIub7a/gTzlPLX9
BxLT/oADfur0l4JqZhO20Xw1JwwEC85PvAzKODv9hpCzgbFD8D2IgWESee3SEMY73GxWZ3GrW9dV
igOfC4dgb8XO2evij1tiVPe+1DJKFCgGMf3TFGLb1zQthr9MuLYLCEZSXNGrqgIlulbO3nAc+1al
MqHLJph6s7TTMznMIPKFuITW1B+CpwEhR6vuSnfFRsVwHk0Q7C5gGIwWx6Zc5yyHDygXExdwyGQY
Y/al4QTfyqEtXD9mOu+3Ijb1w9F4jTOO87KF7ukSgE/ifekvP3tKDsVJnddJmwOBd+r93cYCxt5q
+dNiRd5bP4+CC6zh5IlAjk1sb7pJ7NxMQk5iTB/nfH2Kl0Hoc+6+7N9MQ9ZLjnjt6+pyJKw6+dO5
QME7GWRhFfyqULHtA++AbA04OZ+brJ+2yvCwkpoXS7AA67WfAtWBorOXejeP6X+k6gZWzBwHP0pc
k/tyGIDGe40p8ta8v+WN4XuqGBw+ULub8Z8rp8nc3C7Ay/iZAh9bqj3j4zZIAgdT1tjbx6BGB/PX
0Bu5K5ZZb5kx2mNFyIE0k9hiV2eZvPlctsXixde/h1GJO8/nrNvjiCsTM8PzMIuU7aqXR2AgNztv
LsiyE6OXQYNbIBFaPxeIfivfD7aeqhQ3K02sy+58LaZC07tL0eXK3NUSSyqXRAQDZdEbYU14vA2Q
eILABwOcO9zybJMAjNTajmB3Ya+AtS9TFWOYcg8BJ5ChNyYSYEt99EFS192xlblFWRN4v9ge6/jt
OViCYZ8RTYgZnI8ev2Xu4PgCvobn1zdQiBTYFnbzEAT1ZpKVsqJkfx5F4XF5Jb9m+acr2YW+X5wo
YxR21S50vI3JuV6WXjX/N3Km6pmSf+ZPLHTM3qksY7XNjA0vJME18voscRjjqgbkcJp/70ajQOvG
Gc35heYGzFQqtMhvZVUdcghy3mHZ1al4aCW+TTrpnGaqbcjIYRTQjhLyNB6LR6wJr+7Rojp92fGR
fc3E4dCtHCAQ2vehL3WyuYDscZSXeaxmvyFR1pthymD1obhLtOOE7+YerjlF/L1K+vZuA9X+Ofr5
hl61KpBbDFfIAwPzEJXWPlYqsvTPzfPDF/Gz+HrBSWsljwR7jShBEvpxP/lgTbrQXKdVFeX0eNLe
1MAerFtucm0FJqSrBc+yA8VNFesRWWsNmrXVGVVufqqxck1FWxT+gQd/F2F9Hbeh/2e9fjUvNCn1
W8jaSqBBy9rB92PvOdlNM5ORDP7DD21M+XIRuYAliQOrfNtR1m7rw5ynGx/nVehIguRGFTat+yjP
fgReZQp0i5iiXPBc1tPoMoeAh6R5eL8+s2SiUOk8L8uXqAfRHWeRbmy8lFP1HxBbTF/djgYrwljE
hmIoCKxLEnHewvvAcaRwCB9z8vwvKM+x49rwbvyoUT1wWVuPh6w2mWBDA97Z/b9odWvwEX5PoRC9
yYftVJmI5JWzavcr0Hfn9YZC+U7iEBzxtU8vY1Ot4eMh1lgKt4Gz8MzJPYbQIBO+jJmNCPxjVKgw
NkKzpR7i/Jb7kAzEPFqUgQ6cE1JAb2AgG73mTDafPB4LMxpGfs/g6Tg9rBtOIubY7DzbfKhu7MbU
fVYiK23wQ1CDQ0TbaX7i8Ygm4Y0T5fkloFfaAETwWwl0/MusJK+fwyFvVmAuCxUDF4sZD+aSlzn2
6Yr7wsq1Tsq3n1t1t3w3q2+2/r32vS4g/ATCLBTn0ZHY3fi1ZT2Xkkga0/hEKOOT8WIvgOaLlHOg
5lrv/zVlIGfwWOkNz4+wtbG2EcSo0RfbMRRoZUzoHwwDhO2uqw/h7szhGHumRZc+uXgWxJUimKwG
xoZNWDhFSUfvQXBzamZRnUyUa+NQluhjJrqVa8iZY3U+KXcMwso0jCUIBTAmSB8lecdSceItnGA1
1Teuofwanx+vVdsFXgNEpZla8p3yHpOHWmAICv6BvI0Se2J8eFxrUxDORY73966afAEOJsK7jCDo
AE6egL//aG4dDkt+v7yEqVkNtq9CuyFdN94hxs7FdC1PaELwBIWjEutAdh6NB6BG5ikAX0hG+Lz/
VUvYd+L6HnyWxPWcoGoYtXVegd6D9nUjWinz0KXlXroZLphDOGjYbyp+ZO/WHilm5S2VAr7rYp5N
QhHbpPNrQ/OrAd+4j5JWmEagshOMA6KcvI6mLilTzbGlUuefaRom2YOlb0W6y867vI07xTMuTqds
XeSw9RCSTmaxCCM9BwkZgLgDWqvYQi3uynQdYcXoAiFabnlkvLt/6cpX+KRa2H8CM23TUlyr61eY
V8n1Pq6vPbyDSmSC2mrOErBOq5dIP8NccyiohmgeS2zZ98tbUVmDFzDiTjBgJ5dfYnu3/VHimcky
9QrM42pcXotmA2TbRyeShbyDWH59J6OJEBURzaBZV8JWvV6RNa2JqHC2fhbtLFZ/Ok1HnTXqrlqS
5OcAtmHmoxdayQB7ZXEu+qpBhzxhqktqDX/MTopu9HTArgFkgYwJ5jb8DpXGNm7oA9/Dh94UgZva
MZEFskjWx2ZnYdl+11T3N5vsNuJ9RTS525Kce6TUbrF3HucJCkqjFH43sn27tJhAlufwt2OLPbay
3Sng1IMv+p4aU/+2MIpaMEQNPGmZauwn+FSj6g5QqrFnsVVRw6B+3L0lak18ju5gVhJ0C+TdjoNz
3wzBiNIow70rHDMnzzqWnYcMdZTVJrUf5GUu58Az+C0welAj6H39cKfndc9TcjGNJdluhnP+bIxD
dxcMFvCGpSe6p7OYPHskP7hyvBJhctz+lWf2wSgcVtd1rFlWBkF2qsdPtbOnD3Tf79KmMC3+w29v
JbUnlgN5Y48J8fLX/cZqfYNn5a/TTQSHtgwBigc2jN10BFE4heYDncc53qRof+0nY+QDgFmXkO0M
VYZnbdif69hLnr2os4gPd7ekmH3ShbbB7SAHt6WxLI5wm2sX9bKleL8jGSHXlf+glTU7YlAjs2Fa
q3tN5bucLt/OP+o62L5tipfgWwfH3fgIvtgdkf9H533vjh9uY2S+oB/NQf41bBOiNME6oCKvoazU
tV+XHFbRMsEBPp/0DLwdOII/lCWWVFXOEfTdq0pcaq+dIdRv67ruvYKH5M9MXPind/17nYgIZ++u
Ds7vb/TSznSGQmv3c+alP9HNmW0JFkRsO1CJYuB02yzViprj/Li1cOI0KnAplZlxPLpaAVkie5BQ
+bBUz+Ib5B9yilAbF5f3604oNZB9N5SABbb92Y+2u11MnAkllduDvGtlhlBRnGqWv1Wu7VfRSDWC
s3OrI7ibcRRBRHBU3f+6rUpPMgkYszwCclLiXy0S/9gwZNb6yXEdohXlwyubI67FIh1gfA3UCqMV
JLD5+BGRTnr5c/rRPfO21FR87xsZkTrmkKGMFV6VPnUnMs4mog2GHCcRE0sM1xDFxG4P93vGnox3
j3Gi2b7Vq/poB90H+roR1YqnlQkZcPPs0RZVNdIU/UICxhm89I781q88QciwTCT26fKMbnSr0EFv
/sj2f+NVAeIvP/S/MlMzz06G9/Vq4edcuTkGdjbnNwxdMM/B4bvKnjExGibYl0GTR7Cr2FKDnX5k
nY5X/z+L2Air6OYcCpMPV44oLfGV2FtoJz+ZfLYXOsmxy5yqJbYv7bsBmnCzYz5VGNvk0N+bg1Px
/MwjwGWvvE/SRVV8RvdTFMEQX1ehjOfxK9P/S1XXl017CUK0FcAW/bHW5/1BYegCQAlOZmBxI8j1
Xp/kE7N5GuDD6kRVEbKl5B5VvlYJwHor5G9mxqS/j47u4oWk7o2XehLagNIghQyn0VRmt0ycqJpi
7S+Pmr0VLTqlHah4qcH6uHfKLPXDYM+dRpJcLVm/MnthnnPZDMAtcByohSk64qJYKKhjQCa2+72+
v9x9P7SNhgbzuYppNbpXvNe7tDCcIrv7hQeP7l1153+sAVjhr33+zp/8dVdR//NqIACHc7Xyf5yB
jNEVqUAV/lAZJcA+etUdRGlpZXLktyeySuV6/JzQw4gq27O9U7rNgv9wVOfGvdfqwpeEILPhBqpE
aQIslTBKrnfduj2qVP0R2Zwdcyl14FQBLwChPhBNz3dGr4fBLOjZG9Q14Rj5FGS9jS6CDZ1PNRxY
pXmV9rfkCPLHpa5fcMHPXoMRlirdQEkRmKP+Y2LiShCeyHvAvXT48B6/j8OaKshk5W+orDIwx+5Q
kl0qrycsMwr8Rr2Xd5E1IzaOdaRyhHECG+MOF0PxBLxPTz177ab2N7wdcw2cHsDwlo81xTshuhQC
LCjzPyuHh/5hIWpO9l2GzzYgMILDzPBD0uI4rHAToDI5Ac1hu7Az9M1c4R9JSzzOw+1SpXvnxlko
1LjnbqH5Xsl+Bv2ACPUaoSEdyOchZWg0YFwX6WnOn12W8oNapRyAeec+TmWHswtuhNUaCyGUHPSh
1eWj1AewayDU8lHuw4VG7xtw/r505Wvmd1ydcZaKQXBjLiMZvtHN2+iDFxXgN6lzY9OjQ5uze29/
q2tj11Euhg6ZCkVbOoL15UjltvXALCE2S7gKGe2w1XcFfGikWVqSYsL6Q7NOPVThLFv+79KRVHil
HCdWR/TSHpXWQVBcQOxttzhsmv2OHmtUIjUoEjiUGs7RlegfqR8frgGVb/B91yNK+e4uAmZCyQw/
ns1F0BA3manDOjUyIusBo0VRxrvvox1e2kZ5jg/uaTT+Hpsv9RfLbfRiGTQ9HqC4pJy4q7PEHHT0
qxv/+rTnCjpnHCs8ko5H1mMlM8COjM1OUFdVromNBb65eS/PPuU5NRj/t7fiPWiBUZcI+YRVdfX3
q6atcvkuZE/9jLEKxATEHflbFrvXa5cA5Xr7/cRMgxK77K9AFj2qKO4nkXiaq6c7+lGp6IjOmEez
4ECAnV5e5tVE3nnvSVxOlYexV5RzcqD9W/nrZ2AdK/EtLYvJ61G90dc8x4Z5p+2ZKY7WeIDuSmXC
Nvxw+kNcewTtJINpLWjGk4q81xN6wZIz29zV7KRO3X7mQAHii5WX/i4fkc8AWEFN8dM4BboAGXS1
2GghN5PZEYtzOKUSGQcC+9vpfls9m5TMDhTujsMI4RGbr2O1N7foMwp4ySfi+jKkIcsdzNIq+FEH
TAUBuvXF0w5HxZYuGLQON2vpApTpgFWPxCgbguK6Kz12OXe+fEogepgPTSiyrr02ZuaFJgRuIvW2
hxT5Zrzb6xLr+rDIW1ue7JHO/TR6CfW1wP8+Q/KOLChzlKsHuAWoEqEh7tJNa2OljYCuRqN30kWK
s0YjUundwUZxvdYH4mtfK3xbRG6D1OAYr9kviHLknfLDxUlP6tD/bdRVD7IdGECLdsBhAYg80ih9
Q6MN9LWXQsb6imaSgQfR1bfVC8mjuTbOFZVhue4GE215F1vj4oiBh3ztw5c5fKUjX/010CHSwvh8
RUoBcXamtt+5YKWWP0PGyxl229dCQHaaQ+1C75Q/3wNDmeLDeUptTcti/EBNEo2tpQBrtIB5GL34
2Frk+lG6of1/AzBJ0IImvsyFN1MDyAw/Bnif35NyTcOgpW7uaMYnyH8Xp9rT1o4i2gsMOjZkPaCt
7raOPIRypuFEDKPNDE+AW6/uo3/65g+wf3Ptnr0FDXwpr7axaJzGojcHX6A8cct7lGTgC+EiBWu9
t3Av1ouERUhw0ie8kkzkoxNy1/2tMHQrV3Fw0ZkJuF6T23zGH179mvuhzFG1+TPse1/kFrL23JPB
MZpfspxVNvrF5hdJH2xJvl7Oh1s/PA2b4Ow5q6Hq7fm8yYQJ9FaaHJxoBkfb18InaRVDU6wNcU/V
jDyye3pRVqBE+PtPyD5cYb0dKxUNgjUCvtkO4g82mYF5ACikF29Qgzfjz2otM6+xvd6WzmAUVY69
bis0XPyAvPBg4WToaoFB6RNboXV//t3ImGzNon6hLqLViQ7ZXl4pWs5NdYaoiLb1DON/6hCgkgaI
3W0mUyoHfzI69tgbqxDVSREL50fL7YeSvTCzQuzyGBdXR37Ge3DKWg7AXRr3ECI7pp+mxa7CdMay
0w3b0Jv+Bm+x1j8EWlIp5qTkDk5lYmdwnHfEq6zdX9IemQMvZs6sJjbkn/5BSWPOav8vVvmK51K+
SN50kYai490TAW6TllvtG2kmi9qQGWu0+ZeIi0HHcnA1y+cRGMPb+ue7nSqlwMo0bbgYTahIMb/x
mkbq2d0d1WUWj8uR6P+WSVv8Ps+PLkf4gKJCYtSIwUyf3zGxRyiW1v8fA3mvfebXOJCHgHj9KFGd
x+weAOW+I/IhC+n5dho5dr9DNKPvtLJW7UF8lzr3Wk/bV1vOIs2t4cOfVWZqfuukB0kGq9/33Nfb
/7ZvAyMayo/rGX1NLZSegAfs2kUCQTwCXYNGSktjKRNe6sEGIF7/x1rqCYv96KEIIcteTQHALNBZ
TsUDL7zN8+wYor/FofeaYQOrKqAHLQyLGQkR+pb1XCtyxtuF+YWOu8p0dRTF8+n7ModcpPftUAQ8
rudnbPRc4KJjoAxTk/0a7rDMvYPDBfcStVnWP/YcHFndueyGMRY7a3RQFcXjurNR1kWFMYPtN9AJ
/3AXDNOImg73yB9AMTc80GTl7m51ug8V5v8SocaECTB0tV560Otis3UOAHUAVx7LTx9haqh13Tt0
o5uO87nBW5BfNHYixQUxtx3D+VK9WMVQGHUwUJYcShfIEgDo6ioi2LtiP08DFDzK6ts3G6hB/ldn
bphwFINFSK2jBGBWAyP7fZs26g2w4N5JgDveRrA/kwG7K2S9L0MSUMh73mzFkXQF8QKoHXx2DnG2
fhohCIhedmHzSwKI9wRCiqE9v6V7REvuFkJ6AbgoFow/QV7bFjtBlphjjlnQDR2TdOlH37yGYMBI
JoxMYGThGpIYmUdHVxnBA8qhtjdFHr64Knd2MzOLJ33l4tkil639cQZ8haEhXCNrOPIBLUWvPk2Y
dThPVLA7san0lCz0mnGADortFxF4RzAsX7Z00SBYq+aJoc0GYSNdPloiDj0yUTY8l6zBVcTBP4Pi
0mWPvAzfd+Um+5xi/VpwLCHRabRGDQAOlZLxFqWqWdy13HLsmmISHlaMGdBWUuVWx/8vn6Re/1fN
3VwnhT47vgj//X/p9cKzD9+FE7/h8crtrO9TDchdXboxW6w3675dKuImxXlt1eFYdmuOdHhtWYVg
s2lSH9xvKqQ37OEK2YUmKxd9E9TciLyfvDzNOzbQBG3jy4hgt94ZdqTC5J7HZRyzbHrrLz4Wisf1
PxX5qxC0lge2KEuNlEWt+tMNJ9nyijwsHXHAzmhKCNZ6oQDfxz8J3qtUEnLHhZkv3fgbRR0BDOvO
negyk/zTij8s299J72l7o0ZXXtLN1ftSpW78A04y17Idu45rGzOZdc6QtWW0YWbz2w8xdGLOS1Gf
Ggo2Cv+J5JDhKUm8bxGcX93vWYOVte7Nr3bAq88QnZPH2G/SzNGAGrOrILxqqFbbwTIxTcLOpmTi
3RwEQw5WUwY5Y0EwHocV0PrIKcSa6XUgNKbZBt/MKgGKUpX7ZLAcDRKrgpOHV3ZvqjTltpmJ2sKS
9K7fBDKikA1t+aZZxAYOb+B6CrCOTzU9M/GsLGxi3+oES7RRStPKKeaNwft5FhWzgMxDKnoERNDx
LbRJ+S6C48wEflFRYy1jpLLzFBkI0i94U07Ds3d+1NdTGFU5itSKBbh4JJXMXEUkZcIQaUFiHCp+
/j69TMSYdK+59Ib3qL9VDcBiymjN0SCLqAow7lyvhXZQgrr0lYPGi214iK7qp18HYo8aguz9bTbJ
h+T9SwTISZltWUxGPAuj4oR54fGcbIPnnbuW+jh1HYTwur+UA1KJuFMnDsaKdsh70/eCF/OvqjWj
6dCiHoN6zG9O3LR/ODfR1NccQ+VPLSeWt0pvHWbjg49Ibll6SwetkxGBGnUhI+rED7DWwgyXscd/
FkFAlgXepsJYHkKMeYK9l8nqgeyMYQpKWM7GPgj6PaPMdAoMwlc4UFVCbT8Slj5dMMjvuxMR7rnM
bXHK8cfAyMeCOMeYoPDiSeqXt0gi1c0pA+yfPkv5uiE6fG6xeA1crdmdBR5I8HGHyCtR6lW58JlM
oLzAshaY9b0uKTUsFKK+02h0hKcRlr3fHcqD5vvfbrj0qoufmDX7KeMLdbVbG0yXMt3DWRWI89XC
aRmvMB5zKEmKxQVidLaNfzPLBK1B4J7yIY+fMEt9ErHpT+kRU98x7dVyzLp3Sp3bq3BorQsXamx9
Yk9uJ0cW3ExucBwUGbaJuVrUS8+kU12vzaE7FjjcjLsJy/w3uEN1f/HmC6OfrMxEpWHKWbOwK4UP
TcuhAY9H/DImRvmN8i51CeBzywipfFXf2ffQTDpztvQyi/AlqANjQvpyz71agSJl/h1o9eLFpQ4E
ROXUf2SxCrgyXfTKVLT2J5W0vleBVvN9AvoXwj3DGyMBESulapzDffBax+EgJ7olKpWFm1BaunXt
PMeHAOb0WBRo/Cm5452Z92Nltf0vmruSr0LNr8T2jMg5a/9FKCunEc0A/VdCGnAzbVP4t+2BoJLw
Uc+CVTssz3fRGlePJl6OR4QqRjRt2syX3BanNbAMNStvOFAMms2hwU6xEe2CP7QOeXzjJWH3+RuD
Ugon6SkH8ijarrv1ogVJiyGbLjTOeBHycbhiR98idC3djpApzoS6SfwWPcyg14tI90ECda01V7bh
hi2MLpKBdKYcf/weNqhRCJY0sMkmJsYZ1DgxoNaG/jOBgLvlRTJjIefQtgvYrq5amYtNSpvPzuko
TZ2ujJ+bcec11pv6Jo1G7IsJGsC+TR1hawRg4Z72tBDxbr/42reY+TT7EG2RJOiBW5yXWommCLFz
wl4O/coREfliRo4qke5SChmPkGwdevSmSVl4fC7x9XMpwEO+LqJXRYL1FelnBfBF6Jsy5Poyh945
IlnGmZLP2+wA8GnaI+87AO2J70gEkOpSlY1M2ZlFQTcMC/FpH1u99Vt6WGwjxiuZkExEne9k6/ND
Rd82b+go+IlKioU6AKRoFsaZ/seu5Z5MCIfpH8HbmKfKa5Uqrz0JhTdZau78/GQbcq6SlppGGzDk
gVpRrSi/+wYbEgik88/UsC1DMOPiDUDmYRjkWY63k/0cMCYZhvuTkJ7bh2RAB81YZk6ILdDmfhEl
VMM3y0O0wyOMhPs2cvmiWFC7N9lPTBGThmbdhAvnf4S/2NxIj3z3Pr7ahlx4+oYixjxUTiu+dWxu
WaofwKYJ/EFRKlv5zO07Iuo5ib/1kcsq7rak+hmap9j067S/SuBulGHMrV6Jw5y4UZC47gV49SO1
TEPSDNbwCGIZqWtGVKj97SkAoNjgI0IHCdsBh77KI/0d2oA+JFyMVmj18GOfP/BdOLASbCwL7M3G
492ROJTDZi39u+Y+H8WAMT/+XvfSuoJbpyR1BQQbhUdT9EU4EAf5GB3i3l/K73tp0PgwtzaPiRVg
2W1/QOWEG4lLV39g0X+CmWItNFiP7zAc67XXrc21Jlgee00nEsKUdpnpA40FI8tQWB61Otdo0sPf
ajkmzOxqgN+aWcakoK5061EwJ6MR4Nv1unZljHLTir/JcYYZqhBwJovl/kOkyoypAPtJkL4ntBu+
rPyx9TaBv1WKXWd2dI/f59uc+z27TjnA/eXAR+t9bTo1IeOyLHzrH7HT0D/g1NFCOqwdBWdf3CpL
nClZGndQ8p/0TSD/r1STmtNAXI7FIcic3sbxvQ3WtG9fh5fnxBgWCjZtQbRIOHXz1wa4P5aPAODI
oYhObaHNVw6Jt0HMN6jNkr476TN+25ApilVYoFXbs3Z0sn5uKvd4yeOJtzir6Zz7F2azfEm886yO
vbBKxndM3yXut0us4p1EZ9xRFsFzblCr4GgQ3qHB23Rj2eAS9VBO7mr6eu7BZ9UYbWCzud7AxLuU
4eKLzVw9bk7f8aEloelpAWxw2dX7lRXGiGjrWLo5KsuuM76zSgcNW1mze1HvDtVudAjaa933j82q
xmoI9SyADXdUXk5GvjwK06HwSeF/nQizmpiYs27TEaIiR2c4d+FZQhtWFSIxD7kafCLAhxtPiMup
OCv2nqpcp9DgXqyd85YAfzUFWBQKl3k7zSpRn4mpofSG35WrfsJpW3UKzr8EzGsCe5LZd7bIfFFh
Q3rUCGta046O44oNIiOsO8ZiSa6Sm4zVDKuXkMOU0IuN16AsyOBZchitJuoulwSDKj25D/C44+YB
ZSyYWA03PelRVp1L2YCnge7ud53Awinf77zJsTQ3TlF8g+UfVxJ9xKM8gLdMoyQ6Afx/OXAZadxm
Rb9TRIE6DChSK2f6K7rPx8xSk/0qh+uYO5Gr+LU58zJht0O4CKY0wqywhXZG5J58UQ0QSordtefP
TVsGWSHoP85gxbP3lgAhkEsN3yOdZ0YLBVIhmGV8wlKOYtetHwVg1LdrFawiGnINyV4Z2SJg8oAf
Vqy5lLmvp0xkjeHc3n27jBM5R0mpFjdj0IREoouxmNMG3IP0O1Fmd/KkkG5sdr8/igUIVaVuGq8y
RWQFnXDUknCXfPuTdC6TJp6vQN4M3GiwS1alpoE/7k1V14oxXCopBPcKL+Wp9sdVkUkbHWo9XSgj
R8pQb2IFZTi2cPQ1+SRimTN7f7H23RFU/EFZZJQtFS/7lOvohtc6zpnr4A9KLhaQ6Q1lGN8WB1PF
hu0sc7rwNLlQFpYHkq8v3kl12uM6rUlCdGBs39IlweyQd0H1UVG4ScycvU1cWnpEGm3TyssPyjVx
T/WkszEBr6A46V3om46JBS7pJlzdo/FinciqYRwUpd9B8Gnd2FDzeE+OkGwMdRI5tRv7ucvjvykm
bf6kiNxZyOCM7Fln18TSGWEVpPCelKmqE0jHiGs4h4BQ+KtqxYFGGmzxftpDmskAy9ByjuLTFx5J
99rmrRPhMpKT08R3arLxbDAVgJ28PbttiYfiUqUsXP7Gyist3bcpnYfUoVn7RdB3Nkz2kpI41pEm
nKGXLOt1fGHOJaXliLpXaFV09Z6BXFhoPeM/9D8N7iWtnqyKAiBfonm/wgRQmcv4XUL7WUis2MIG
YHT9XtQzM1cLXUCHRF+x0NzN8K/OIYjS75CeQgpqW4q9Jpeet5orT47k8yxmuBkRIU5d/pR5Yj00
OYSrj9e89Gz9NOlUHFjgHoRD+ZtNGMml/tKknFeOQ6QnXGWyIt7bhDBLWdg1QJpeJzo46N92DmTU
lwl4Ga4fdte3N1k88sdrQfA31RrQjtaWsCAePSelskIrY6fPaX5SuuFEN1nf3imLR6cl746gucYB
roGJoPBeuEUGIjP8Bjf5vgiWneo8LGOGaeRvVBVLwb3vdFUIZJhMFVxYNAYTuMwi9MNVp4i0KVO2
5I0Dh/X5lsAXACg4HnzEUXVI23wPuHQdNNuWO/2reiGehTKiqM8K2lAmV4mEo5e9q/6FXWRLQJrg
2VNyFXVfSgXdPKgdrv/RI9osp0w7XWonXtJHojPZpN7L+liDANqOjs0Z6LMtoUPR6UmGo7Uc6wig
hcJMKtdQNHm3H+BxG8rJoeD1QH7A3kfDzyN5aZ9OfiHThzMyFbZHYA0TsQcR7UO4C/mu7oN7WnNd
ivgGEq4nGVYqkHjjI3v714B8BknB2RqN0vIymJqWXVgAIab0OuFt+6IxxUBm7uRd21rpP7A+niml
cXXJuhWaN5ZBKWdZ2rPs2x0FmmdgNbaAM2U98BtaCd4yHsxiQE5ZW4EUtQ0khy/rk22qVsY5ho9G
mMzfvZCBEmbw9TrqXbknEbq64VRSVOS8iXgM8oJPHP0QV2QWn4ZyUpwfeVNK/H5i9xvIOQcFJV1T
OWnz+7gCdG46Rjvpv/YFG7ikBzqZh/A33zl0mgliQIjZPqXFfH+ffWc8cChCVJiHjLoRNEOlDuc8
TSE+q6yWtZedbGUnxX9U9N4DzKSls2MGjZzPdajJESrpykAQQA+uGkgs7XS9jeCWFY6pZDzFDEf1
M7pSVCISQlHylmoKlksUmcqIOvE2pSGVuTJlAZcIxLCg2ld+CU361q8G1KviqANkaZNNOGCPq1zH
xpAzAc3RDuXU7jlAALPXSitgtAeW8CD6m7JnyZaOGTfCsBdh4bGnhzuj5DeeespaYeqKGggaUKJG
aJgbvxu97vheIQtxwY78g4o0TYWidIW8R7NP81epjRV52pZ8dl9II+10o6Nqi2l4TqJ8ivjjgDC6
PY/4cuyZ9dZXhzRi2TJAIn9d5ftXtsaAwCf9bMoqiIsmV/wYzW/h4Bcg34+8z1nBsNX4C9lE+2ZF
QIklxCi8Z1i+G/sZFijvZZA3T1iRjSv17ur58th6RP1K6wnf3geBc059hmq5o9SrIZ5Hha5n+wNz
FXVyRP45YiE1+Qvy5QAMKMMy6BtcAnazLwYRZ6e4PzkZc5YcRLO2iw/+1iJnLrYlqRzhViAewD63
cTDGQga2lE9izt0qFwMSE3ceg2iMwqBonZNz8e6NE7y/zPcGaOagc9Wf6t/p5wZ9EYP/PFA5WlR6
MZoZEkxqNnrpyJn0bmsjKbvCP7Ex+IyH1A/yHYA2cVe1f/xC6notlD9tnUhQh98m2fwOCYc2ZuoQ
UAMImxLM+JcVyWkibrR24jUaNhbaX5VUcGFPErucoQ/55KmhTRTKQN3ozFisXoB+k1iF4xNnnDdf
PC1q/8n8VfaShTwOaGeqH4knLi9HGHzVtQ47zrr9YzgtNDikxWsLH1ysF9SCrwcfivOcKFv4J5Pg
avXu1EY7TD0yIJF1377Fs+UmxrRM/eTzlnlzOAqg8V7M4uA+OrQ0F9hLSmovGJiC1vlvF8nkiUlC
ooshr1qfkJO6NCP1UUvQi7uMp3CMnz+ZBHzUMqbZwFp25x3Par2whbe2d1QruPb0vGWs5FxcXw0M
1i1lfJbowVrdHypglDipcG0JlxUMEoEZhMcvOZrCUl+lscvD7f5sFlxnyKB2SPW434GxBstDlo54
y5zl1ijkUduvjexq8EfQI+uKzbtoh3sYwDwLqul4U+4Hyl0DB93H+zt/wxRU0Mz+GlNYf8e902l/
DE4k8ZkfQ3olAbgHew6PgLuaBwfMgqFu7COUgmK90jxL+Xn30ui6gSA5Rt55157pEcFblJ6XYpth
F/OKK8kLe1QUhxyDaJo4HI0/7N1sSDQmYb49uMlN0Pl8DB2psxVR2U+/qy/WVVAWZzn1Lj1UqoJv
bHhM98VLSxFIV7cXxNC03NOsjpq64hAG/HbMYclp5DvCMNkrj09ElbuekekrXqo35bV5TXeZudW5
UySGWByjJP41aTHeg1MDymzmSRX/I2yORvX7OVEPyp/GeJPXj8PP14VtVUInNTfpAm89s5zVXF1A
Glu6ZnNBEZVigJB4JJxx23BPQERORzDXETQ/Rs6mN04Lma/qOfIF4YRNz63tLN5NgGQoBnrQEqgB
Rp3GI5dXjevyHgOfkc1+cGCNSHVM2P8zU9Rj2UHtT/zKHYknmU1irVpHSntQPDIKEC8/UqLqdvB4
OPmlStBqJPCZYswPa8MsStlioNRuhxyl+OYf4ufDaLIdNYj7G+I/N7Ulw8jR8Lb2bIs7VgFXCIAK
umdZz0Qb/c+wUlUKBvUj/BdhYzyVfgBxSrStNWWMd5Tf3efTmD4FGO3YJ3Tc9dJ+ZhdF+vAN3uhN
UN7ZnVCJnl3QcWwf10ThcyAlQgosrRyAzVESiwi/qmX3CVrT3JD2aRk7exIOAcVote0pO81KUu33
LbqteLP5HLagOD8ilLfOWcCNuRfElUeRflmqag54vuQ+SCGvkjAMRyXlOkjXfj6WTQIAw7HIH1te
RpX9kysxe220ozXjUssr77ZA9DdaIjA3/f/uUjg3qquCiC2QZoEHlF0vEl1b/hX5F2yOjX2oD/W+
hchTycpBPjzpdByC3R7BZObDNCEZ00wxArDrdaSwOama5T7Lwhb3RikqHIsl5IWr/hw4l+Tg9apo
oGiKiBKixVg04U8wa5Z8TQU0LELwQvaDrhNiOkFRPBgHG60jhtFtohsa/KSsn+Vwgt4CWCynKyXR
OcQ0XX2hJgkiy2VTxLx4XE7PPz0llLrBh4kyQvZSdcDzd76z1TRufRtMk++TNjlN8DsX4HrLyWPi
JceWqynsfApmBS1D0h2lLiowRutAUUzuH6MVvke9AkN/Po56S5kj/2GltxonBqbaTB9Sq/lqzsGv
NhD4ZqghEnf7uy4Og3AAAZAtNGGnCuk121+hl/Y2ayYSufS04gqpYu6vCrsHKxjISg6lxzkGorer
wWx4IzvFrZZCG6bQ+EHxsdYgvA7/8OlZm2R5J8wyBfOOz47V8eNmw53dqmToEojKlv7y+M5t+fum
ObY+HRdK8f+nSh5NcLc8HfJHZyBy/RfwYLZ9l307m/9dleiNlqlPkuz3ppBeP5zirVYxw+cENkAK
XlTZCo6wGZq8wzNUHcM/5DN7F8/W72kDsHyWLGBoWlDPu+IGOlICX1OFihE/0repaE3N3kqEMfhd
FbnUZ+TzQAGwn21e0G6jQLB/+Bc5fbKU9NE9Z73Wwh0EJzibXQllpaDvj9qT9MSlxqXmOO/G7Ale
Xo+KsZRPDJV+fWh0oePckKM/Fxp0oPaFmjZB1ssBeufl7rcgpWUz6VAAAifKMrEtso+KtGiPhdoR
mG1YSWNqZSh7ETIlo8BX+vB6V9jxpS3sT4KsI3KAGLJFbvBgazVKDY7hWgR4VZNf8pf+QgCp0tNZ
JzfBHpoRDyL52OT6PzWyGghsufjpA2hR5DdKh5WmciV7XY+ngye2uJ/aaJ6kysSKEX31RA3c+gWp
7Bu2rxzFcBJKgzf3xZmufN0jTOEX4KWALTtpO6O1gE3oQTskTkdiADgfgU14DordpdH5+rtoWAAa
dBGKrbX2hOsMGqllKcqzDsTr74THu0Yp/C+AtdDX2JkxBo1V1D4RgwlKrOD9BbrDR7B0p89J9lLT
g7D+XM247CSp+hEQHbcplotFdptTkya5DHjjXbEsqvkl/IP7ZCCK94i6duRODL8KWjjCnWaovkoN
ETx5nrjVKw79oIyBRJhIz3TXP+aW1mEZa3ZCtVlH0XILwLfFk3H5IZ0iQM81AhG3aeSaJ6SDw8xH
CkPBntIiJrNUqrVKVPC9zzf8oHDHTt4c0uTdtGMJ7eik71h1yOzt3Tlb/+aQcPiHtVHpmuU3CIMt
kjk4kjbdMttaXaQ4+52Gt9Q08t00N/sXJEo3DTWJfMMwado2DI/QJtOIOPfJJelwsIaAyW7HqhD7
S6uVRtDWT4LKV0M20LbOkammqAaUpBT3HWqa1Lzo8Vi69UKcDagK4AsJIu0P03DaxqlP1jSjxk+L
7wuvUKevbz8R/OlkcBeSkxNFKFOaaob+33qmEI9blKVJtNIH/2L+xjLIP4/rEi+qHJdOgS5r3jZZ
gsPY0TxzTp7hK2VW3UW8r3EKOX3Dw9JvWSaK/taWUrYf4eGeG4aOqSWT2yFlpl5F0w9jzX1/3+fl
5Txrbx9tB8hO4eDDRUVRRNMswG+559j/o+FsWRcqygrD1n1yun5PRLBdBKjYFM20e+yFvpJA5pfG
EwSKKeUqbryU/SBpEIAglW5oGEQi1FOmTWgu+w8vchWJJYTsnWBfeHqkvKnBvBg1xvToGGxzH0x5
aTBUSZAWFdf39RQSvojTx3j1qVnfdX2z/GX+v7WM42i2+MolsDzOdOg6bvEBBC8lI9K1pGdulLcD
fEzp9uJrSFVMkF9ZaPBc46KT0/7Yp5WNtrWNPLjyuLsLmd1ndEs0A8BAPbwCLS8VOvKFcQFDd8eQ
CHYuyvycE3eQYdi2wNv19OgLVs3MO1A+FaRI9l+LdNN/brjw1eC6MuQWYo4xoLrldhL2sYuFTYBV
cpuS8e+zdqO/RMixA81OslVLjUveKTlyQpC4i1Q3oprAoIkpuhGreBPL4FOK9IbjRb3mWKBvWm+3
/A1DGZ1X4yaRZ+fyKqzWOAPHFl2y9DglGKNnkrHCiJsymX/TufF4RuaFHhi+YA4poXPp+8SyXAp3
dlSC6lnZeDU3R2VzYWyGHSvz/j4Kb0SxnZD407U4WnKYa6gggASCo1xevntprRb8bm11LG6SModE
VmGFofcwkzqQuPG6GhntkPZgfWVIaGVieoMcr+ZL7+J1P4WLcDdBHAQqmCM5fqYOPl5welDZnmwE
C13cY2Sm3RX9DP+JUWmXuSuhJcG2hOk7jjWN0Hx6flGDZXCW22tVPouwDSx4umM4wpVe9Y60p4mU
f28J2yBVEC6SIt+VbFAksOuaQ+5PpQXSaL77/tKyt8S8MvBmxLNem/LU7un0r68M811Dl5ST/iwa
zuJbSmc56umOw6iLBUsrIh9r0hPoYam4DZeyAdHUvo6evovXHjKept14ETEhJZIojyP9boCaLwVD
iCqQqcpQe/hBuFwKzCg1U0T4Y9iOOvDznpGiFunPPNa7pF4p+wlziHEZCrT2SEY1vV2f6hA9aOpO
zOyxFepSCDCmhL4rjAJ6y0r8GDAUYIT6IhV0Xua+kBnouHZ0zjcVo7yY1tGhCHEVUknc3ip3eBHS
fQxh2Io7UOitoTjQ9N1eNmVB4AXEHiVEb/kHqKtLrmLUTrdkOROF998SPe82meKgPpvIxr7nwGgA
9MFj2iBhGifxHQhJAeCpxp1CvuuY//wPzVMGCr4hDGo6LsbYhgiSrdlIOULOtY+b+Gllm4IOHFrw
Mgw0aJzeRtFN6glPfDZ5ayh4ZKf6UWfBVtpENYGbIxHAB8xbJINNSlHxZGfGE9QwWKwkB6gtPx5T
1BP9ysGDAkl27QeaIltxUy9uNTzC4Cjp8YQBQTGnfO2ybm4/rcj9L/g4ZIZt30rJjsHDzmv8A35x
R9mCzup+GEew/ZvhB5+HQ3Zh7/Ma6hEqH0Da+spaJbvAGHX76/E116/D2soqFIyF2DdxK886alts
nmXG0dbFYuB0OdJSFu39K/JUyor5OUc4QSbBk5qo3mOoYN8esUPrTxttSBYSYOQrymuequ1Bkaqr
q6yRHWKRlEXNANOUAvj6m8JohiEnSR5HOkY1iyAG/OzpInlWkF/1I6YBChGTbGnQN0cb0yokFXBT
ZJvH/sg4VbWPQpy1H3G4m20WUgBfJNmhI9H7YrOhMw/OexuHdCv1fyAcdvmO5JSW7jgI1A1xGc67
nL8Y3N2MVAaaxbHuo3hi8h8Saq4wk96LKmLymJz/xFsqbCnmPokNP1oqizTo0rE0rwRam/RTPgyT
NsQhwb9vjk7zaFLlRtZD5I+AIAe/IDezlMfKgt6wgURus0U+BuKMCAybJDCiii7Nla9BI4sPt5/Z
Q0xy3c5Eg9xXPgcAG1SoNH+ufBi8eGe/CdvSTW64QfyO8ZDqCNsKdHJny2X0heKB6ey+Vo5/OsNs
Xm8fKsBnA/NBRL1vB7gG/3y05tGAf+nmGxE2YrtfC8dVVIWrTtYhylpcRL4hapHCTrIEDVIDCEGU
ldTiz+jhlp0I92nXNDMU8SnyzZS04POj69l1EmguCLn8arTRvVetMBq81I2/NuDTQHUac6lqiQ+6
wdbZa0b1yyXif+ceXgmPeivFoTEGnTtnv13Lorj/dLxE0R/xGkix23kAWMxOkVD4T6RZySX1nzbO
GhBZFcAx5KlLVQrfG3FBJrxzoCrVtE2LFP9J/LEuMARewN7HLI1cH7P27uty5/LVYYWE+FiUs2yM
yZcGDg0nQgREOSgoxyRNdt6qrg6WD8+hc+nnlqm/uMfUKPvysXgP1yBs7ieZQIXzx2i/fhHHe9i4
x+Bugu9gQFlXr3QxfeGOvXz7QRNPeURdvHQ3+HjSeoUYfdA6zUGMx/vIMHu0nER8vlzg3bPfZX/W
/G8iLAIPzBtQKNoJMSTyT+EQnJSsYRsP3HJQoVSwNm6yXTPX1xLOPYSi9FhTZB6B5J6ePO0tYYWC
U4OYuo19IvT2f7oli90m/elNiB8Yg/PzPKaEfE8hQIN/zLCK3xWL0IWTDrKYDKyj+2cJq2IGyM3y
i8TE4BOAWfRI2DbBFTsknYL36TcElgYYKvmmvGdz6M461U8iW7bMtNfUeoNTX6P/4N/9XTxbXFbI
uWQPQkIRuEa5GLZDyDf0Qcu9kDsRm1hsqIhQQp6IKHNFWWQryP7H0R0+ijsFTDp4K+Dq7q/jBCgY
LzuppKNklPxmEkwT/NIa72hHwYJNHLUwJ1XafRoR7rOyPoLi8QzV96s3IyXBQxd4rQzjQivxKiCH
n8BV/H7fWu+v9Nkt44QIhj5M6Lr025aEKcd82qWhQPbotZI4wwh/miGqg04RFN8A1052sC+wAMnb
yD01n7qnRE2qRPtYxsn9ae1Iw+IsR7xZBInmTRfpu7CCNw11/Q7QWvXexLtb9+OXEtwVHdPcHUCv
aMuycvzU20ztqMzUWKVD7aemx4TENsloYVaCn9JMP7LIjzkBWA2iQBGVAxIIM742bEkkMuUlynzr
HaCbHxSJMsjbqTj1fhganETIODp5sy8uso2cw2w61ZhVvaaI1lgjdjHefLFBcZN8xQ+njbgM2LEX
5rE8opOWw9PoaOch0/Eva7vJFRitzp4NHrY5DiVIFBVe+paGaaJ9m68bUCwlXuEog4Gb2PQTHR45
1l64RbGN3yG6KL7pu2wQ8UXJkvxyihUxJfeJqopaJegMOBizqgGGj7/EXgX51b5sRhZhEwQhhoz8
R1EGlQfhp2AQz1XjRIwJ1AGqK7s7rQzxC4h072hSHWTYuZ38btwlckjJPOLXNUzg1KtcVNIR8YjQ
gsGBYrcRmUhNG1hqPgmRdIEQLLALWh1UhqkCgvlyq0eR2r6/Bb0/ZDeaataUI11mIwJuGneQchUy
v+ODD6jCkt7l6nd5WuSqo3n98PiEvOdxmAa9eQ3dgAVNIq/4yE6Mj9jGUUZalICsAmKguBDkfH22
hS8jqzPskwR8+bILhbnyT56qmvP2PSjf97ltvstqP/R+KGSqdtmCkG0fWLfSkQHV0XW5KRFPzUJk
xllYBehvd6rJSgSXB8b59pnQNg407IOFB3pG+1+trf8nCPoyO3fBGdbsg8bVVOpsxmWxWD55zrDt
IR28c2u+OfwkBGU6BwsRrkJw4Kp1OLBazD2vV7Y9PwaLxgGShleolj8BICP0sJMputKv2oOQWiTL
iMZtH8w5o/gnIkW6WbOdOC3zjAPMCl1VDVyICkOXrQPeEIpFm4U/vWZQrwnbPBMKoFg8yr1yeFIw
99pgu1X1avOrGazFMtXXveKq4B1cgoWBXj9g7F9Ce4L90pSNJ4y098RRkbTnNXNEqEK3be5qbmqc
ZA4CEIuxcQ1E7ZG75OaTXs/Gur4e4fsV4hJkwgjyNcNTJ4bAvKvhpJI9T7PepBWouyYJAvwDY0qn
NrhCoQmp3vniZ0FU6AZaV8ict+epHPIkDbbQDbEarT0ffnlx6J2y/6hF+Hqb2WPW5HHPJT1IWXBr
TFupabFFNgEZyrtjWhnxJ/8OYHL/5FWdxD2BhvYBTJNOX96oYd8tcuw7E2Ta4zN15qDI1BbjzLSA
kY8ZseDjYm5qxH3y2QL9p69HxYFMUTqQD1tPYJJUs9Yv9akAXvmS8qv9DaqeJ1aQszi6hr2Y3HWA
DHSMSX6TSHrfQVbTN4g68B3VBGuZGEx9izVFlrM7C9svi4ffw6xxk0yV269kzy87HayvI37Dytkt
XOxJNkqcbdPbE1zZhgHaa94H55x/CUjOR7rJ17RVOmMUpsUt2cO0TcwwOdG5V+C3GccpYnynm/Nf
uiezdW61D+BFj0RJth3tr1CQLhKxQOKnuw26XPbfV199nrW4vyF4hRExbLhIk4bBFxbV2wLbKQzK
sp2Eo89FWrFsNQHkPo7nsW5KBesdP2DqmIfKTrGxsLA0gObKADLUoTeldDSgXh3wP6lITpFoAT3L
N9ysKYKmmrDXWGdEzZNVmXCszYFAYonAOk+Q6YiRX//OHgGP8UWZ2nB9LTPZdefrfUpYHl9U6dQp
wVxOjFUROxXgStE8UOP/BAz70pRizJ0CMWbuLUWe7ciPcSwLJxOjZV1BrxmyI5Qn3eJZ/YyxXTtR
qQ9dIR4PgCb59jmHW1RnuO0z4QQstD3QQ0zUzcu++Uu4stRnbBLhDCbCyiSNmrtb7aDxufwPcvFA
nOy2KyKo0UmLFKnS7SMJJqCsyrHvv3ucrElofrDnX2+bOVVsQzZT9ENH2hvoZvJG7N7ZlwUnMcsD
3Awe+HCSHH2FdvWyJEzHYgCpT0RXRF8b3lXAW/Ubfx4vzVKXf2ME01qMz7WnZIY+vaolwwEG4wsq
Lav5FnXxszDSc/6Tyg3v46Yxf4jLoqqosMpvZoP4NJLS7AjI+UQ+ZGJECdy7pF800WVjGynOBKA9
rVQ5iho2+yaXxLjwBFUKlTc/4K2PQngtk6bcz65KHeqZDv0chIetnpd9YD26MV+GEBgKIFSN9ScI
2xYIjX0dSKrRHttQAWkzRtljZpGOXCxrzH8dR4Fr2Utp0I/3RhSScmn94g4NrJg5XG8kdt6ybIK6
jH0bOi6ctrLbfN5OCfkq51ihCA1zbAzOcB/XeTOYewNN76v/IX6gHypEHKM82XMeeU+0KhAmJWe0
yYN53Nie1RAUleVisq5g2bnyS30xh4Wbm4dsgUaOvorx0mwgTDqmAodSB68Z3A9TQJ4MiCpwClPF
Tkr9uGjpbj4jD9VpLmnamw9FQQvLet5LRRxonGG1wJbBV5eGSD6Ltwm8v6u9Gphznyktf7x3P0Os
QsaAvH545hvpXlYY5VZGbtsGlI2UQ0u5v3GiHo+8MlEQRp/mZBarlF1la7jscq2VOvHoLg81MzWK
ZIcm6edGcmh43WPTM21XJDioPffjr6er7MJ9vfV+gwH7gtFu7g1WGFv+QJAkUrFjn9eJ1X/CroJ+
nB/yAPYpJDV/A2ASPZyqBgPSMLHJ502F3a42l7+XXpaBfYhF2Mh26w+x73AtEvdz+yIbpX9p3+Nr
MxP/CABjA99BbeMCNwNeqP5oH5iamutPetLeZbTAtXMChWyCV1icppfhCVtXRjcCPfUy00xD31zf
prCa46XZo/223S+hg5+kMxsViYMBplJ86Uqvl/DKjsd+2U3UQNuTljXIvRAcNWnttOt5+fvfONoK
AFcZBY1V4Xt2hrvRf+FCFObPIeWRnnYuLgq304MSfB62zJUAl95VZZp+eldODCz1NXGT32czSWRj
jIniubqi/XDxxYXxauBltI/XlZK9k+l7mLE5/X4ORAi3nPlw01ehBXoDbKv+3vqo3T/l4HII0Qd+
WHYJptFzjv83+k0wkaTZ/cjW/fyLA/CfY1ZlRCRefXNKri0TuCwQk8zWu37kLcVSsjUABW+2RtbP
jrafVKjizG9RnAUjAMWQI1TLiBxH0YS9ZMwRTWY+CB+9tMVbRAUX/yaqMc8YXuall9iSNQQ0VYrd
7Fx0N/4xASpdzfQvD16B3v7hOIhKuCrdmsIpn3X9B0XpDLs7pzvQ/YLCKy+7CixFGw17xolL9SE6
C2pC76CwKy4dutSD5GHhTlXL/+bhRvx0qdOtp5gMqD9TbSMmXgBqphD0yMA8Q8kCU+h7yrqzphhu
m+z9B0Rdpsv0FU3xOB8XkIMPheyyRnZw7gRVNbAMurEOyMiztT8QHCtunfXycFFWsdu+x6HNoy+l
ejwH9ZNITDH3tgZc35pM5VdzTZNVLd6QDt0rvgxMuFpyczf92EaWmtYZb7sP1EI0pme0ehGJg5U/
Sm6GRQJPGAbd+wbA1du2dirnPER4JpqWoQvKiD4WXvbqg3XgB26kkS8oHM4pkEMgn9SED3Yn230c
/XeK4m3lC93QAuydHTzAHnwY9AX5AsS6bQwaTnnl0FIGIO4P+eUDB4vbU5JC690roX+lNqlLQ4RV
O40JbOiA1mtEMQ4MV99k1X0P7cz2HdLpGQu6xG9n2ZMdzX+AygmL6USPwHju9os5FRB/e/YLfAW4
II1CwSBH8nSBlKb7ZwP92PiTmhk4ayTqi4Ut2mhvFBf/z4mZRzHSZmi54ITW/WRMRamLdPYkmwnI
xsy+DTFrzJolacnQiHRbW69hkVaknrgZqnW6zq9Vn+TC+16mHEUWDqJ5P6d3Oy5xkyFj/hHXt1A6
4SdTyoAEcRlTlhIorqPUs1XwkYEQY1m60scdXqem+wjv5HNoNs/3/dn/5IsWQugutc5xU/7vy84X
hBvTgMOrznxWXEk98zNBovWrAPZIVq7v/AWzA9D16y75EDJhBGPodHuixnvGJxHd8wysyffkrjKt
GGXxltMKeKDbyx4W8gYfTYQE0qtgx7t8PLlldezAv5fz9AppqyqRkixUvf2uZP3lssw8h6pU30vX
jALiNeAmx1+ZXc9LnW7+n2WBFcDYtzL8zBaHDeJOt3dgLZaqUrvgDYBUcXzcuTfLcnDCNWViuJCv
ZQAJqNO/iW2iTzv2+6q29g8DOTH2GoAmLtyPiWT3ETPHsBsV8avX1fi+78C2U/ouRFSbeTxqKkQR
MSW79dsgiSYXIpikFdkgSN+x8+xympt37P681UtfYdpRPN+c0uQbM/CKsepn4YEjS+dJxIa56x73
upI6ugfoD0Eb3K2VQTeJFPKrFV9aFr8QtGu4VU0GUA7VxXkaiBiveXf10wDUXHYRoxhObC4RGcU6
spDFDNCm18L8/tIUtolW0raWqMgFO2mBPVQACJBVdUzB5ZpZ4M1y19Ed2iD223iPvymm4FDQ0nbl
LuokSC80JYnPjwpF+JasRp53sD4aKJL+UT3Takxy2OXj+jg4CK1DafoAIpMWDDy2JVCLZuwy7V9r
cIvRPH/THv3QsJjDH3ebbhgUvZRrgPm+7vKThKIIcp0EgIjqE4WHUqR1TcFdodauN1cPFn8eEQNU
FzLdftRErjpl66x1CNsVfLINcTViEv28P0RGaPFolV8D3y5qoZFC+lMD4oEC5QFzzn8+2Y89E4P2
y5x3b9R4WQM+GEO84TcOJFS1Yp6jQXb3i3W55uneenDgYOeKzy0dswXWt913NcwhE0bRLmcl23dD
OcVENH658A7mICRI+J4ih9WWWNikOQfPd02brrR1TFNALCy7jc0CtDnM39QyUWJUNlr6cuB+hlMA
rqmUTXxqnN9xXAwXWAdCX/bhVH/SMKKL9EjspVCDB1Em6/u5IsZ6d319tKPV2pSzjVKdXfJ9DThL
hW2wz+BRaIXnGxXQLLNSf8BfCMdsnHj9MHZV1ONfFQs3oOo7lB8z3u6Aiu6ZjUgFluLTRFTYDsKj
5+Du2Vij8BAlrNhFI/wSNX9ISmPLjB6ZR/Ap7AhBWCW1VrHV+SoVcTk2jRoXrrzzp2GjWn570Ssb
YVlqnpUK0j4wOhb/xz3a+2c2Tjk3yxLM6r0FvMGwPEYe/jI0n4mHAqnm7kVmyCR42Qns0Le1ebpC
0gQCnoA3aGbMw+Ffkgfwf8OYFRCuQIwQfkEi172c3JjVK8xwqX0NWMlDwLJI8C4ch6K0XepwQXqJ
nn9rzIGybHecLNgNNymY3zfVzK5Tsipk22Lk+JnCB4PzbxOGxbRkABgFzlOQhYnPepUDlba+anal
KwY6ID12TmTyl5WgAayEH9PmO1XgO1ivXwf8mdOHwenj7YdwYYeQWY/hJhT/kvIeaFkeklyI89Il
acAQ4lvFMuk1Ah6ViTHNzNgL4IyEiDIH6ME2I8vO+ZLgT1gnqh7liNaPnMeTZ+J2Sq5/kq0SMh5c
1mz/7337lVh5VnE+o0FewT1qcMOognMD2rjJmV5njcNgywDPbFaf/tDjZ+ATjaQJFrWXhAFMYH/y
EoOTgGt5fG+iCeL1+AUvpb73gMOyXYfVqlyKiUVN62RUP98kij+b027n//dsfmTrD+KHOwOMrI/O
OCSLAKUCoYtvhZhhcyRpsZcfHD3Nselycd0zUU0XXPX3EX9JEIA2ljGVX9foh2/KhlwLpqeC8u7I
QMziq88/0GNAKsq31/wxoQndR6An4Imk3kLqig0+njPzP/Ww098oV3JJf2xL7Rvp1y20IMof/VCm
XZCBHos4DFJIfK8Pd6YorAndK8nLLXcYAWTdgdBmDLyh/ofnjA/s2ovOUAlwQR3RcY5o2MZXRKdY
X+OP8PegiyH4aICkNSzhnpu0X8rvi6EeKN/Fm3tq+oZU86ZysHh7Z4nXfVZuHb957PPrOi2XeScR
znF4OfJCmboIwoR0KPagjfuAJcETqJ9heC3j7BQhOBnA5GLOVAE6/rIc7pHHkrIZ4SNUF+kFVe5i
jlAIeEWsIv2sYHDithPwh7eJVbTUQWoilkbb0NjkqZr7gIb75U8JmrFVSt2NkQ4pMGUh3tIpInYV
PeoBwoo+CUH6ByY4VABJXjt4VZDetP5KNke4BfxHsNY7bRdvNNUC+MHizQlky27bD7GLJcTBViB0
3fxR4GGszEDxVYf7XSQr3oxJKsUIINzy4pDq4UMn+Yo5n5eT3j18/RRjbpafLm+YtKPxX/KgNDqy
0omHzRkvuLr+RdZWI6ZTIg7+Ykq7HOJ2KAJTta8NFLzcX37VhBY34NHO53G97NlXwAm4VwrzAFCl
amBA/vq/sAXq8tcBC7wlB/j0OZTeGtx6bL6q5w/5Qz2QfULl/si9aKbXwBzvVvJEv62imzQBSbFB
r0azGDS4/odED+WF7ZF3boUMkiB3Y6OSMNmeXlRl68GYMcH14bhAL5Z5XER8i9XsqafUp9E4wLyA
ESakxZn6fUlD+IsON3z2aH6fmWu9YyK4X3HXb/mDWK6r0OFG2aef0nnZOEelrhl0HBt/2SlTj/Or
FPrez0hWMBXO7s0fkfhhYPJ0mkx/3OQr21f//O1H8qcG7O7vvcvRajgJJDucGSvz0B+k+LbYZQgs
GhJ3f3b9NDUjzP4xOk1bvoWtGdrWdzb24gobSGmaQ1ykwD+GH6Ed9hv1mpjZxJjyO6iwX7GgFSTt
4c1Mqg91Wh/8fOB5WzlXGev8ytoWzduvVJuIOtXJ9HYvF5oVFCb0HhQge4Gf9ddX9VflQNvey1XO
0M/4S9hdHm9t2bT9EP35XLidoSbE606+eiVN6omLJzjKP0AvgvW8lRVbStA+MVgO7HZ86MeUhiqv
Jq02tXY9TyKe1v221OkjII73sDF+WtOTzQQ65mPWqtlTjZO+926/SUAtOOvu8x+wfN7ijd4/mycr
ZBAHIFV3QbxaHbZ0z8w7cxBZtll8cu6jilWDH4QIll/1wa56eDyjhniWZuLVrkvM8PNoa9CPTah/
o83bi0E03lik0vul7N4lkHkfVZWPtxlIq3/Oby4rDjrgZghd1S0cK5EMN32yzBnzo8JnICAPPNz8
si3W5IiZdTGpfeXRSCoDOykElM/DHZDIm/R21dCsL7ttu+tqKpQvtaxRlKDkKzVQOIgFRg7mSzk9
LiiHdweFxJeAau3zWDvccqM7wWi/ZW7oF806uHAiBwtHUPC4UPOezkesYEVhc4vRWE4LotrhlOnD
sJu9vfnwjiyDMTT4GIrmeLPRmrHNL5xokExTQ1jRHp/CF76ftjMuewulvFzjOxsPxMAkDFbDYkeM
JsVhDcPW/rqLGeiPvrVZQX7LACvfGXsNyMHJbyiR3xQahojSto1XgumPg9wh4dLT5k69AcoK5TWn
2QVdq095t+WcDWRyt5R2tdnNQKG9OUbLlRihk4mJ+Iq2BhricwniUc+/P2dVOcQNlW2HtPyTqZav
268p223dgvm54sQVdcABEvDKCWi5+l1i5nusrbKmxdDs5upSuYTjqR/IXGwPqVa5mUxjLfO0FSc8
Ozx9Zj7Iho3QxZOrRA7LZJCQfOuth8cbaq+qetwEPb4BauUgBzt/3ulFvWFVELUbodkm41zpGOdb
zjyFzyc7Od7X8tLCsXegoMQYCCL2zScPrMP9Ux9qwBQ5BL/B9EH9VgA2uYZ3u+3YbLHSfgBbLWyy
hXKbfVEqThAzi5ZqgD0y54vFE7TwgzkQw4wVAJuE/CM2KbZSe8TBparI4k7dz9MI/UuBkygWK+fo
hbGP6Gtrt0otLVDrfVza8AHIZS40ye2xE9rEn/oMCAAU4Lm38A9/HQIdFbCgRHNmOfuFnYlU0+By
JQgYAPNEuCSw2Ocoly2xeAdF6eIpAXFHmkdardoZfpO2J6o7Z5TrymcdgYPSFqw9L5RZv092HMFr
Q3K1iwbzJO2oh+i57w4hSuQkJmF+p653ImCLvb9V2YchfJDYDR+p0p40WrS5vANGE/Cd+vqnLTpE
I7QdEvCy8k953+ptd/IEGYWDs0OYaNTfgXbtdGcIEunlM+QcL8BohiAEP0JqYLIh+rg8ae3CBeU+
ZYpXoR9xHu7YwJ3oCWHbDRzPKWyYAUDdf2bWj5DxguxW0qIyLBpVeDX2d47HCJg1ug10Tl1AkzH7
DOmV8bDjXdH3GDn6z/w1IGSN73HAO3y03LPEHsJqpZsorNQkKdHi0Ucqi7q46pA6ycOkkIjoZMsD
NNko4Fb8ndrYscwBP+C9e575OFr8GGzXZXun7mQSUvC7DGsJVJMT8WlaNj0XZMhuAmSlvW1dVPop
EBkuT8u9MMiOfIyfr7+R3Ga87RVr/LVyMZnUu4eAm5gDIOiZBtNU+1JVUE+HiVC2yhluPCJes0d+
HO3sxX3FMVEyku27PYwK10YhC22C6yuBbPmC9n212q44XtdzUe/OG5Xtunh8wywhwNEdBycrrGBY
i4FoIXYpDTDEn2DQa+nCRmavNSCSUZ3MxIh/PoTgl01hE8NDaHcwGNoZU1WfrvftkfJ1oMjF3Rgp
UZpsfhdSG6d9aMgSQRtdmWVr/uFa2h87O96sqQ7Wa7GQQdDB1w7LIn69RoDuR51uorii5wFi8Kvk
La1f+484pfEHckxG3upukF0DOJYACJ2IhHoI0e1pwtZvkMaz2N0/e7QRvKyKKVhuwZfnTjkaSzGK
Vc1MvtKFiAa960KP59fQtrx5lTL76dtQK5WVXRy9RKMuNVxllaXQDcbdkN1DnLfwf+MMf3ZtFaMv
qGeMte0EzqdymRLw05MU5RmheKZ39t9sO4fhZlp/MCKDREH0yBwmdOY0MNUgaUQpapN6MOWBvI7i
s+bfEAGWn7S+pI6SS7YkhFgtpCAhP0hOKVCDJdUeptJXPlBMK1cJ1wRlxyQMad0j8uaTOXEGBw+g
zOGbY0r4l42tzqMoDQB5ygiyiDS2hGQEVzGI2U1bmgmCQgaO8FkSqodP5nur5emGlx2a1c/jC/NB
NigtbsI3Ky9WcLOSqnSvTxyut8AMuD0mdN0WmovRtREHd+zayJ2bIiMe/05ljXbgXZHnVR/7Y7VT
E7nPm45DnSUeFe6PZfpDncWql3qc9tMXWQbR+ie7xcz0q5g//X6+z7ctuSmH4/59G46iILwdnFcO
8aTBMQ72KVsvvzF+P9zj3qynLIZdiybqZU0ILAs8dD7PudYHck1K2edYsqhCwiKiaBwTCyZf5GGu
86OC1EHToFaGBlsLWie7Kua4LZvBdzmQ3Tw7EXRNv2d2FoZ74iFbtd8kGtF4fUDFHjckVq91uHyI
AO+E6hPzGrkL2UCbrw7UfDN4AVzxNPThgIgaCx1+SAUbYazTrGJc/dIKXb4ekve7uaIYk0gyphfA
BVCp1nEnhS6RSil0CELPucZ3QUFe9/3Vrea/1m9c8tRbpTtboXDBTMadOwcWqug5aa3L7n5cScFR
oHH5VfyOckymZwcnmbukJBanpr+dr5Ntwu8/0n7bOiO0s/84arXcbOLJGKvj/wQUHNhgiAPQ0Dn2
5T98yNYjsAmw60yAtYK56hcvXZo5kKu3Uz4U63T4AczRykqaNpzF4iuAwwVksQWXGiKVLLRBmI/Q
fYN7CcUaAsUS3SI9mUXsWdh99VjRR5V3ttcyr8FLGVJjvmL0kWAlMcPVHiIqOEl71Jn9o0WKfHKl
z3gMbFmO0qEJEzrTovWWTBCv6tLtq3VAWRtIW4z+dnFhUcavcqClF/ofZ1flcLAlCNxLnWfFfwvV
E+1cnm8BkmGz6d3pLeBWvmkdO0G/3hutwDEwte2BsSvBy99ylquoTOHJogae3Gpi1+IWIQGnIYdx
dLMKXMALDolsq/ZFwbP4b3zGjEjait/p3Dc9VfwRoTRPBOnoDmfimNXRav+olxFnM/ABdBCs144l
y8mwseH0T1K78ZE4KrYBEMeC9WaTyKIT8n1dtqnIqlKrwOMq2gJg/zjqJFrwRdh2zZRuzA3JuRbQ
9TmxBVcvgByxPiGMt1uQL6ln/Cg68Sg0lDYuNXGOrOm+4nmWMQz/XbuK1oWGV7QJarbt9g0Xd7s+
cjvzjV6L5wRM0K01rwDYU78gp1JjJncqy088d3N5a4esuAulSRghaxlMAc2hDeepv4qDRpt1JJRA
27KBEdwQLmSjsAA28puncfhlmtQzJcjnrE+dswuE/klf14IWUhtkL630/Ocs5Nb+AklEgf1bZ2Be
OBuPDANtPPgSsYpZeFdHcwybFV+sEshtFrYYTGa6mMScfvxBvU5pSaEK6HYXseF6sLnOAYc5k7T2
0aJD7TS7L0IK21FaSQWKv9xkSuJw0MUr1VlXdJY793O3AcmxntuMBlwf6ui3Z1xp+vzQOisUg8ez
P9+toSsc/3gDvR05JuM3nltNvxrYXwLS5gZdIe2/64QhQ63xjoGg4Os5Uf5bZCxVMTmDxnKl5iGO
9YfnPRexECJfJpxHL9AJe18B3cPEbdMuNur/I68wMFH69srjIGZ3GAnJsAa5FHLMjOR4a1DqfUJr
Zh9GM/QGqOpWytviKR40ywphP6aO/Ah12zmYuuLAoxu9rg07Eq8M1LNV7SSYQg5v/iYwlmNv48iL
1UzdFdXh8/VDv89S615CkNldewT6HnZNiTbhc/lJtOK6xDg5Vmolln7Pmu5+xdRpQzUYsNWM1nwu
6g+mUmUAEjYbS5whJhgdAu397KQ79Z3/Qmce7N0u9qZ2Nu/T4vfsD/UjyFC+wp94/A1tOyd/Rku/
aJClOM8zzIptDuoP9Ol7s77Wnu1ImsNTTwhw2Q8pJzYQM+jL3QfhBQCzCo7rloeSDiYZW1fRIU8b
hoqIulfqwwC9rk/YDs4K0xe2AgsL9yhLIic9MIzrvqh1YKUwjonXhE7505YLGQ9P3GdZDqEg+7d3
DDoOxvqmnF2bwk+nP//M2X5MQG1gLbp1QEzVRDj6Sp6i0vrrfgfziAj1qXkfB9j/L8vtUpyuHLKJ
oAhQPwH1hn1558IUU/BdVG0cey5Y33KcaG6ErgGzCt22i9tgXspxhHmb4BaMuC/b8GaXAfVNFdcc
ivK7l68aQJkhstSJgnx+m/D8A5E0y6c7z638v7wApa2wQwXocmWQ5ehxoucGnifN3qn9g51n2J2R
Baj14X5WZKESbLwpT/d/y5iHACM4SNBlyjOljs7ATldqGzMaaSGv+OpWjhwc4Nu6WYxBEfIeMW/D
DOgTO9bkFdxWLhIYXRFzpHlHOwcO1JgE4IqR7aO5y7yzSmc3hLNFZefeqJSotKmQLkOvMhnTdKqN
UPCKSFmn0W3Fx5hmsG673T6p63lae3A5dGYKNDYt86w4nUVuPMw2D+eXGbQDiJA8QsMZk6DM4NlP
tu6jNe3sBPsZao/+l+ZRHQnEMFGfg93QEcc4Ga1oNY+5mfQb85w77ggHpAn189zAFFWTEvZphkWS
Z6HVtohJ6CGANt63D4nVxZlktPY2HSr70/7yzFEG7vdm0LLXbFO8H+BFS4CDLlp35T7riLDKMoBB
QXBZsJU/QEbvIa1WzbG4JjtTudVAW8f/6gGMwTaNh+ClppY6HPB7+nWvCMF7SG8y/6sL9ODRk/cU
FzkMzgb6s9NiJRQUMfJ+pKfktjD9rk/IuZXRXXxkFMCO/zlsKNW2h5xd9+Z7Q9Jie+KKZl0rVYTI
nUZncFD33ZANBT33j1diZHhe9qa9c6USGneciYZAiffZ6tvZOP0f9+JWUJQPE8hTg6OH/8efyvd3
rKkL1LglaJjrQTKVvfle66uUGQrHcpoPciRnM0OhWEBLs5dLVuBuzOkVfto+vxZ0F1c5H33L8EUE
S5g1/HHblMpYoZWP0jVin3J7M3ZWe3npGhQ2wYvcOBhOUQG72BjR4YvDIHzxfTpiLUNjERmdG6mi
yP1qmiOMDCsLtBA4InSuKjWrk9FAu0cxSueomPcpcXJtPV2roomndPPHshbuWKn5jsMOjuXsSwxS
JCElVK8El7INsGC8Frk054Kqs7H46QxezAL63GT0e112gKzS1pUVRp0xlUAaN/MYRTT3YQAn7OYS
u9/yKTJAfcqrECqOE6c7x7Cp30nyKXqNge4TrlMkg5q7Eq10r8uG7fQeUXnJF6wQZolFUg4ZZ1Tn
BmG3yvO7EwrpkVSgfp3IcxFAQfKr9y48g8Hr2XW9mdtOY80gbtXjPwzsG/4nSEkcCHrGmX4C5XGu
w5KVnJWNmVLcpRkRlnv6BQk108aa4ENprniiXoYPT4DFHog3zmRORhrMasz/TKRq0o4WmtXMTmCW
WvZmNi9xruhhIHw74ox4PWhfmMw94TxhmA+OtYCsZh6r+qYWPZqo7iwFDuDY+X2KPc87GOIiV/BM
XVukGA0FU6Smepf7QGb9TEWaV1QeQai8KzMagGs2XNGrUKyE5eaRNO08OxpcmlzM9qjJGZl5Ag5R
aNhWKLTiDdH43InUPHNiC6vnS8uViynsey7xsmdqWmgwUmLiFvp71upzW2L0ECefgA3ZnWlE3Lkp
5VaG8IAkTeYTyaLkVd4FQqL8jvBT4P0MzbLgsPPWYHi1B7blg+9rcv81kMgpfF1lT00GQoqSf6hq
WN5waxbZX8b/6Nmzkpb0+JLZnsgnJaT2tNO5ST8q2OmeZ0j8ZcQupKnZb73ki6IbTCSLlgL1W3A7
EbumSNzXk3yFkePh4AC3+B5k8kTZVAemhl46sx5tbTeNtVwot+N9oEwkXok2pe2IplVxeUZLawXy
s+RvsxUP5hBW4mqJXw3sUTpkRKOG+R7OJgX1DIoYWp1GqHd1hmOxU5tlafAEH3FL736MS1KwNOu3
d5yZIZvRbJrJ4iKVZoDMAamHmxQbzsHh+5gPvby/kqpMCjC+OyVwDycwB5a6BhBephehFJQtCBzB
CQ4q+ZBj5BNkM+77/gkAjukRBCcuNISEkT/mBf3NiLGnJgFl/qcPoXkj0L/6ZtX6Nsk9TfwnU56I
nYFFdn+cqb/kjQh1F8kn/xtnfcnz1qHkBY/iwmjMZRRqon+g0HmPR2RaQtZnG5VwOdSROXilavrx
4BJD+ipwKytxy33XpBFgib3s/tCQAtUSE9OS79WnHu+PbILHJUtZ9Y0eucjZL/3NtTB9bi8o7Sy7
eg7QRVtx7JScka9vUmp9mmjndGNDUCiMp5+LFG8YC8Sqku0wTVDhL1g+wQmKMXTIeZ+rwMoT4VsO
CtumLy5iiGKsr4c6Pj1kSlcR3Xm6/Zfmb8L7dI7S66NT56nKXtxO5uVa5mPPY3twa/NvFc14BuA6
CL77/FV4flbMfIonqXUVcYT91wWWuMSZ+7cSJqLJSsoVH6Qv9J3kmslEoJ/Z4KR+kKIWnWnELVAZ
dd8CeMaVQtvp9Mb37QrPp+/WCwLBAe8XpoQnwVmTOnr7dLGHDxEw2gjKauhgEJ7G9k7YKrIjqG2g
BeaEiHwHibpRu4HeZS6zUfHM3N67mya08blnt05kel1HrMFETqAVxDjWI118NPIJB8vf0L3Iy+eH
A65CYb6bdfVH3Xc3iAfTNsWgRWMQdNhawzA4zHMAc+rOHt+yLFidIUOq7ooCe3MG+1AYtI2Ys/op
pL1c1fT666oGrhsFrHKOBSLIKf2P4udLYbg69dM/AKibX4MEGMZwMqqSjqVSRMa6Rt4dk03kzLEf
iGKmzlPYVqZ14A1bz973je1F6zUWkZZavfb4sDd1E6uhKLtMESzO0oLrDWdKYnbL34ypPlbDToUW
PhOdCtdpi8EFC7zi/OHAWsPbTohkvU6r+JwOOKoFzuYy964BhLKcNgFsTJ33nj+C7UnBGTOQ4Iyk
Bxx32bqjMe6kn/tYIHRqYD9nStUy92+N5eqJrpG+SUKuocQDBseEc/chQzbRTKAQ5bhCcfh+35CW
gC+KBBn9q7JcEFTKP4CHTtfLfh97wi049WqpFxP6m2nogT6lWqQcm5xgC/CDddmZ1nLtug+ov9jO
Px3GoUUJMtvoaOiWxkdkFgi5abYZUv+npUmViY1ZbdyNz+SoZUrKBUOFUxKfIhcY4Wunl4Z97E7z
I24Ue338STRcsGDGd6HEmvlK3FlHq6tYDITfLGwM5NtBEEpxGHkj0linEYysAG4zA7q0ovp0voXQ
g1JnqEDQvHqQzvbv2kYknQvUaKMbuM3SSG8z98i+NyNamstS/d9xNQrdmzLEkVJJy63hQbT2I9bm
vRrp2i+O5DbBrGylyz1ZRKrHLROg+U6JsglldaVh7rA5iN80vjeRMf5H+FFRvTzRgYnBkwy/pblC
QliarDBf3Jt+rRHTXP0y9ip4j9MwMwgCwoOzPV3q8bbIrvIQ/kNX7CbRuvWszCCyAiKGVEVgH9jv
pJuMuekifNEdTotcl+sbaM9nx4EbJwhlpPQ/AtzzUu+kKnMan1aUC7TaoFV/yGozKxS7Shd413oQ
dEmtbAc/7avrP13Gj95dmaEfYFmAbFtUysQHPkwkwclglH8WDx66PsaEKSwYRP7cm6strSJO4EJD
zwXaTs8rEXSguuiO+POCGCJi/JAzGXMFLfDuA9pyOqYHblbVzaWCwjcGCAH1KEKNM7inpc5ZoDO4
n1FHqQZ7u8aUfKjyfaahk5RhDP7BZ72qAVkBRwaovk3u+NbXm5KT4qFS6hAmh/bzp5dLrmGxMJ2w
Mj8XhgPWuBbnR1OvzTTJTYiyensLO9zH00poVW5BKdhdze/fzm0R9qzVcO3F35ZNsrwy5iZIKK1G
ilugdvKKGkNXPtTby1Fj0v7VxAy+eprCTb/x/DGvU/JOR9CCtX8YS9uexIz805gwjGuALadxz/Bl
PGYaI7xidKVUVLWOp59hgreoIspN2dgWFiOlzA6qbkYxClnKLgEgIeQshmvaWq5KKAfwihOAxedZ
sBjhciyNWXtsndRUVr4muXa52fuPTqxG21SHj0jgHwM0OFrh5Q+RbaItGsJLoDgT0UDqxmmHFdMR
31HGRuX4mkIZc/FPwYsdfdir0Ak23ocdAaBgTaRuWfN1I35K53ZZDF2EWsgi5jBm4Yp3dsmhvfdE
jyi0lgWj2OafFTa0BYkwFvSN8mNdCOskni9jMyGsU1vrOcvKP/eF58Yvs7FUq21x8IlOiUBKsj11
Pu2qNXGB5UMViNzjr0Z9dFxU7GFIMi3GtKe7w1qbIqfIr9/2DIV9T+QWHgS66SGD3lHvpRL5zeG+
eC2/kSm1+30/E0iw2GzQAdCuSJy5W/Hal/o6TUESYxSkuc9KwKfNM75GxVZgJ9Wgk2590mDO6gSz
uioAY7vEeb6wdXXs0Pfy/NMnloJaxzv4Wt67TDWhhlU7aGeXeT78/hf25jHT9+rvuGgIV7kg+VI4
e5JHvzAcAOEcqUK9NtXoloc3IBBltmieag+RHzgPHgdZBW+SImPKEwZu30C50O1rWw8dxGvaAsgi
WjwBIxmN0hjZzEI9Irf59WB5g4ffJLFBpixlU9Sj+kJwOZzTpXOblTQiwiuBfuOsE1+SpJY2XgOP
v33VggMluo8EzfNKIFDzhMe+mESexMCwN0Mg/JxvteOuqHIgfl2Y5DgxOWQTQlOF5fH1OWVgF7kA
GqY48CL8jVx6miFfDHSvi5TFlwp7PcSD4nzmgz64mmI9Fl3FHb/HDmCcrsu6TphuDCNkkIo9OAGy
AdHp4WIcfkWnf/Hq8BS1WMabmYBto/XQtUmZHzXOQoyTuo6r1ItyPPQw2vkOKU+R/IFv/mMQnh2h
FL6v3i0ysCvfVjKN1B5YTmZIUCMRSpotpEy0OnMLFTM2UBqMpm1u7bcV1GcbI4NMYdI1xmAOZchH
tzFnBa97kqHwp10Yt9ZQ3Cl/IGiBWvcszT+iwCS1xnh1gPWOByhx5APq9PU7kV1RXtJkV5gpMi/g
b3QOQnZVFUaYC06h8xIkn5Emkc1cTclvu5guWLxrcaAWnsCsQ3jzx4bKo5ytGZIhaO+CgsNuRVie
0OdeCxkvsGB9Su6DGKnvd7fJrhLsR/cx7srzqT3Vw5qnnF+A55RQvdscQANZ6zsEFG8aPLuUAN+y
YjhdOBTZtMWlMgIawX/EBLG4yUpgJXI2sS+/FZcq/ST9+79png8f2Pnb5mJ+o1Oz7tgRvfRJOL2O
F5zQFn9JBdPWSld079s+2DETbmsiGUuUXaHqoBB2xk0pxArXtSRO52kJOFdGGMwp8y/J19bC1q2x
/wV6EoauMFWgEFy6Se+WEbbXHzMg0RSgyMkgj8y43cuzf+L8eCLh9QwLbZxZZljLcKS9DifiHC0A
FDLgYWLRXo4t+s9qqsIXRwaRGoDjmLTAD4PbCCCmONQ3jnWcKSXi2Zxn8l89suzZHRNOTKK2b4o4
WEY+5GpJsqWWkSA6meejbsBrWOJvx0XjR4NXYa285oSSgMN64v5K1T6pOjdhA7LxBORW00kXzTNy
Vb4peYAygO7gyAQZZwusBdtIVi72fLSwubq2XNsr+rftWi2PHWmI1Xa6tQlzBQQznr5krig3a9rv
qVQFE9qI+pDeytPu7SdRnQSmFKu13BsruLZqbujPCd3zE/bdL2LfEWqXCiQMlm6bBeRoU07vTi4D
k068EcqK0JTRLtiSrK6fu5ULH2bYqXspi/N1yZMrlMAQmQuEDgzrIWTpPH/sV5OqcoKoPS0xD7EV
I26N9eFJ+XGgZV2hXQsf08L5ANp5KFD5H8Ebe9zYutOyEvQ8kVUaG2MnOdvzsKriFDrJlK4pmAtx
L8upa7xuNNCZSkuu7SAxcq+Q7ptk+WAleqlSaIQ2b4K8/jaFnW5wfT1k189BKf3bLEehMLv2TCl5
YdAdumP9nxmMsMUbEUZmjQLQbSiFlhcVOSOOIycXdoslqIFbcgf0oxZi2ucBlaUSkgQdnF/x3TKl
eHxQm1I6pX+5jRLWipVwJYkn/8oJwi0yiYMxuuQhczzumaUj69SjSeSU6uWbf+7iJi3IAAksIRr4
IWeT0ujxgTmIr2mYwco9L3D+7ydtpDkIej276F8jZJbL8eTaicwaT+gjYRnM3FUDVxnyLbRgIDSW
4+n4Ix14kofhrBHZ01rFWeKLd39I8FRTmwQDM1Mj9BIucT+ZcXq4DTjOTWHevBMdqrLBzMtvss87
gZo4mXrUX/hljyJ04CfVtPQuWY3aYufdfjO8XN1JeiBZrBvsXVHPbRxD6DW7ji1IMtbtVeSbZc2l
4WR3ZIFpJ8FnuL3hoX6cXJpWP5PHeAVY48uripnp//6mZvKXtbvl7KS2akMQvJo+ycrmkOADE5uC
bRMuRlBGf/8Vhb4K3wRm7qWuPRtMj7dGb05+vpI1Mhzj0LuYnOWdSRb4KcWE8FPrVT2sHYTNv1gA
C8Vvj4tmP/bWI3PSqVK6cN8l4a8W6bJB4SQvOQGp30mtdQElHVLSK5XWeDVzC+N9BIy1ub7qC2Dn
yVy99XZMUgXvohMNexlNzKX/AiGRPcN2WOAQH4Nz9WkayH3rAi75+KfJmQtzuc8vgO0Jgp0r89x6
T3/7LITHLMyPabCHNJl9S17/wQdIc+DkLAcpc70ZvecZMpSpzLlO76YYuEU2pzEVmjp5YSGk8NKm
S/T5blJFxN9FsEjacIpLslWkHjh4hT4V/2v8WzWNGuZkVyGt5oNw/sWSdVMkTXM4vCttv4gd3ydJ
Y7EbRB2gnRfpyFr4bSiUd+50dkyUlpwj1AV1v401SX83PlvhgJilfdtNGFcvmACbZAX6GGnkbdrw
OraTV+CRfd08mnqIvRemp4cKIV4cwsjrmL2g3xEZXJFmXkO5XvrMQsooaPwFWNL1nppsM2+0x6RX
ADuA6ks0VUqFE51VBFpl9/0zLW5sZ5/D/TXbgwLt8Lp2NrDrF46TYSYZ/ek/V35fZBCivm7I+JqC
TciAyZkn0PVvZ3FwwxyQhWj/pAbWnO9ITzVX7MYjQ68/ZSmbKgMdCviPK4NFj7paCy4lQd0u2xmK
Noh4TlVGwGq+7vrdVX87iwkzmRp0T3Qor1gHJ6QztclupBPn3I8m6j4bnkiQM+auCUxWDFiEAirM
MRdGT006foyf/Xb1lk7MXTQ2EOGqhl2WEwNp5JnNtV0rjLNaQb4kZKT3SwrSluE3kfiKAQ3iqymc
i1hUm5GUHk2O5b6AVPcRCA4BCgd5EmbPdoK8xhhh8lRNFCldCkQardepWxtk4GU8qsRUpbVai5pN
gTCjlcKI/6n37j2oJxbXLi5lJ/uT2heus3vHGsy7jhNKNWvQZVaZsxkkH9SBHIX96ToAnYqoDxBu
g1TlFArwMx1ER4PEiPqURdJasagF2Vc/isSivzPrRrUfROX4opEL9RhcbBp9mDD13qjHxbIqYB+G
dFPHdRQ+THMNK9V+LKHdd73Qkx3YIhwXG0A+q8ESp+G62d1ahLrMSU7cbvoKy0yNlbvxECjwYCJ7
9fnW/cOVZUqWFlGwp+Eb8xO3B0ZPiMHp1wmZm+/V+OP1JXMfXRoW8nOQmuW46feAbFQoKedPvSgP
gdGF5SizQgbXPMaTONBWj6J/Ck3vVQvbTHRHewRSgu+0Ms2TlmHHRp+D6/Am7lHhPFw/IY/MbRTt
KbZps17xZF0HhiHx/v0/5Hq6w9dqjghdlPl14UsdO357D8DedGS5A8tskUi2EgzYku4wDQJAG47E
sAYd1wQ0gphiCsWwd7AQNCAlRp83XtOeML/t/p3XsKmm/ZQ3V2W+EdK0WIYAN9yJMcxIPLQrVzLn
J4PS9zWTwOUSB8FFta6MTNQIkmZSNb7qHmW90QT5V9YsYjFTXde5gKcGNypXoBf2wrKrUOeR8dS6
IChx62DlSQUKLhYXSQHUxKfFmYI1br83yH7zelXzmrpRwFHQu7koy7R4xWNxThnBsNxo7KsB7am9
AbL06n11W5dXyv8HAUpXqKs8y9ESZuMZX9lI97sTGL+EvT/FFCSWYsgF+3RToDI5Wmm+XKF7C8w1
z19vSDqtx7rWZ7EAWcxHA1NYjHXQR3vb68XL3NNolg1D2+FbruA3lZnzAslxl3wicjkjXAHcGB1W
ji+nwzir/WzSx1+pc/RZaYvGxIXTo80Zb0tElHrhtztGFCahj3v0HRwJiLQiWdBqrL7g2lNL2sIv
ZCCmYnwEdIt28voZEKB0pPS4hqNVcBdld3MjFwggyV39+HHno9KiUrFoAawaAU3Izh5XUfEoC97N
bcHuaNdPXdUDEH14zIog4xQCFFYNZ1h1oaEkslYx9TkRSyQKNE1s4Pf565aA06TvEsyaaafwW8Y2
d2gRWIBn8K9MMuDtmBzMBzJogzqWntZY3imT+alvCb0pfMb/gykA8fiq2gyPC7J35duFws2dm9Ed
ZBZtfBr3mK51NZeHd9n4D9KN/g7gDQHSuzvwdLjFEHcrDIOn+gbdGT3nvGXLbRmVjtJhwTyzK2Pl
Mku6T0j5yb4l9dmKVhy5KkisfgFKybpZRZFvc4cq1QRpmw9Ks1vubSP0QsL1sPZyDu5RTLwE8EV6
jf9v1MqyHDHLAeCSYHYPCvqb1Fa9vGiw8ufvLZMsxzuC3WcWHhbxzzW3bs+xvIjEVxDiEiDUfCAS
xLLuz/TfnvZE1rNfD+8KFf4VyriGGS0grfDq1bLVwh7B9qOVzbCrtZFZeX+cT3wzOhzunJPN1zGJ
zZa41249yJHpxgWes8mQOuXMfZmZ5YHxG7+KzfC3Pui52xzLqQ9D6/JE/RVIwGmn6Em2Rvw0nDgh
AheTjX3qo5OLSHqaP+Iw8l7kwipZLk7S24rs6oKEA42uEo5LYe1g2Nhp9ZMRVPy0sWbjWc9gGgbv
D7r8tms4FzgnU9u2dA3L/uitu7CX1s+GxgGOKXob3O47gQzYkpDj59WDjjoZpfMxq1EAhsmd3bVp
LkFPy4XA6MMScAE8MC0DpFS07wFFRtaOkpe62tI7ryePsgz+HJARgDOiFlhym8IzWNLj4gVCG9WZ
tOq0Zv89LUtlHHIozHxDiwIlCRa8UiZ1MwTLFcEclwofnMUy3XULJacz3RX2wEkEyy8vi9nAP4jA
B/aGPQ4oeLvs1CqzqvoyyROQVK/rA2xysP14gU80QUFqPRjdu/ASzOE0jRdkG6yEq1zlFjfzFZJu
M5Ke8pICl4FSRQmEc5RT8/NEaFcULHS6slJnLF8dAtatKnmgrHDn/0x89MlgYwXQaw1ovCFnp9RU
rHTIneJQUQGAUzH921ZAYpVgj5DYpYdijbRZ++I7M5K/Iov3sdIqZGENPDjxVaa/wRr8lD4aN4t+
yqX3yiyVFlr8zUKuXfN30siIt75VKR9hqxoegivAKOZhjXmxQk2A8QScMNMef1lfoj7JyKwNi9FO
xi5waLf7cjrTgP5sXEKOJDBOKgevTDCOnAXLnjaEDi165zeriK66hJnR4V1UeQ3p83AsBoRdOPUs
HZocoQEu5ev3x0wT/iuAfUC92F9XCvhNt1aTDrxOP2mJz6eYiygrG1KL9pJjl68yMYctyuabGswC
uSigbOJpd+4ChBAExkYZF/xj0GYTR3ziU58l06D4hBYqmAbOvjk9y3axL+NpjHO4w3+TZUPvP3J8
ceCuQa06MfIn8YyrERUDafHyjaVxZkHExiSioxIIJFAKxQG6HqIsIvPkJujdBDspU/o4cZDDr7uq
9AHjCkzoI8SKL9OKef77Tl5LYq4rgaeTBihFPah3QY8zFpNlJ7tzlYnik4cV44kjDERYFDTjQEWf
jVNY7Bh92uLH+Nol9ww86Dbw1xJMYLA+4A1WCUfW1NN7Oxy699LhYleYx0BnuHh0YhAmPnjlxg2w
7NaaLHiRMlh8nmFGN1+oSCTEgMcLdll6MB9KpOHnkCNpjcRdutRfiByGMIcTLSGNaEGssWLhUrcr
MjQ7GNNOn/a+thH+yb4uD8OrV036S4RDLoiMIp97mc4TZj1G+9UvW23w4aOtJLL1Y5JisWw+D5hu
irklWHl+haDATzHygQCLH4zRtDmnMww194PulCLOp7mxxSG2wYz9eqMSzVmZAZb9RNz9TPAWVLc5
MhGvrOdfYKA65DA7JbqbynaX4PmoVTPpTkp96ygm4QdM+Xp+vWiyjR0UP4q6o8JyhQsfIBQVJEzx
5rxdI3jMPEragKJimMIjmsZY+9nlGsTTTbM39keilFGHhahaMpZ1TUByg5GuHRCggBcknx3Wh9VT
zVob3nT/LWIfdpUbb4aAtUVG2kEiVJyrzlb2PnD+7NrFwY4Fm4m1aoB94GM7kJtKcXUMK2cdgzfW
nKS+6JZR+c1R78pQdodD/VWEFkB94QGSmmip5U69qfm2JA+WEdZ3i5XYANHwEZnlE9RqTusSbT7N
uj5SFKofMQdUKEwH3xML2ySBARHpkw73lptQmmBN7oHQb6VGs5LOz7XdugKp8ohAJpKwTUjaqNHl
iEERpedAv6OUuPAk9Ww7WPVLyDkYQKiJ7yO485Ikmv0JmcObgwweN7SZK3SMpEDM1cxeRQkXZWhg
5o87pKxwcjnwpKzOmdBlBGxMc3uqV1yTUqdUN8v1o4ZnG0ODyRUZ9yINjMdWncyoV1tMLG+prAAr
Lml6yTso12gvGvH6U3IudRg3ND3oysfn6pQPGA3kSVGMGO9EVpBsK173Z0/AxUCV0UydpnBhS6ft
SL01rB834ZhwdSJVluwQ+zn+wggBT/0Ot85vWOrW2jAsCuJDC+TxsJFbufMNnxL7o1hyiBtqVcy+
KoA8+dNlz+U5/chOBsgqorVYEMw8IBqcXZ9x9JmB8CgP7Iuryojky8XIFoh30XJVOgSykkN1PP5U
pjefXj3R3ydJLICLGdppasudRY0rH5+tsBNX33d0tCj0g3nZ5nd6fvnHxdlf/sL1zvJUhRLNl6Fn
dUisfk3tK8iM/eas2ddq6NUeDyN3v9iOUnDkPdYiGyT4MVkQCckgT3c60TJRYdOLftalPQvlZ24u
4o+6UBGXZZ1kMuJ1B0+U/9KXd6mueaBSP7Z/J7jn1AHws/DYdP7tvenyC3Sll1TB1Q1mwmQMYCT4
atX3xj9+ZPj9VPTd/l1KA8NRe3owlOCxdBcQRk+d7Koj+hVn5MI9F6TsIEC08f0errfAAxoylsCx
BiTX1FDN+GsquEijlPn1vJICgbigQBh8GF4UOPliIgJhWqHZ3+ar5NZN/L2o6SJHZW80ByzFBHjp
yJ4DvsSPuw4NOu3NYolA0FMs5UWmwKMtnuq6rXPnEk2cbFTwlZHLfryslcCBSykEWieTuk1h/xDj
2j6+F3dnhw7pynfQgK94br0kHGuTN9AvKBK74DW2qgbJ/l1cZj/YMnGQFIjb61+tfHJ3PKkbtO2f
1yGveo7zsuH1eDCqQFnj8V9wq5iPcE8Ld/TxmiDnwi1vn1iLWHVkqTrDol0zFxy2ZNftnAAgEoSF
0gV7NoHvBKa9DrvKsjiZ8HXD+6CVcimfK4eK47HovZTsp9JBoICmCZjwNL2p+YzIlIAcahSA+mTK
qO/E/BqHsCvjaRNxvrVcvhNHA0/gCrVTU/vk4rHX1nbGZpDK8GqiYYqhwZv2VG57kwSacIpPO1aG
f7/1h+NJEfK3T+1NM0X26J19dTw9b6Nnb8YAIsPYkNWWYNUQ5oZOq9VBE4ePEXkEX+9JpZosyWkd
liDzqRjY/C3XT6spTiyoQwT7IR/S7fXJqtTbRv7vBLQUREw4aCSG4Kl3nG1v0OWi6pXJIDmv0OSi
nKqWiFng3cdEz5ylVVixfr9OJOiWIXfVtqWn6hHsRfsMow9KOQR6ZV3ofce9BAdvhgGH2OdrsoMM
HncBcEoJzyzdBOTEgLz0RB20Po8PZgEAkpqphZ/6/KfxHEejfVOGHubax/wEjm1LIUsxt7vyNPE6
0P1tu2I50zmqOsfLUOoeUtaYqrMSkXd+lncE2Fi8dOId+CRHNeQye3je14kf0D9O+Wev4dpI8LS1
S+c24iJjw11ogbBz2j+0Kyutlm7MsXE3SD3nE8qIewPo4SuQYPpfbV7U04VVAlhbZVF6z2UwVjA1
N4k0G+0O34lDGBdItWqZHeJIfOtSE9V+9iRcSwghDhkhP8D0/UU33CyXQ55thJEVsmAwwJS+2KUn
w1YfSg0vdYud9qB3Q60auUtgyez4J/gk3feG+3WGpedodelPaPYWZCCU4x//VFgCq65GTy4AfYFF
xYy1f43Di/BlNSIGz6uwxtMEANeJpYxVxwX3Cg6DnIjyLjXpJ1inTmSLOeE+3p+rRxIBzlgYChcD
71ngAo6brAZAvC008vGs8yIjtpN1Pw+MSNiL18HEpjH6Zp3O+zFsSGc3WU2qSaz+5aRxGWNuwpFK
TUl7cmGQb8Ndhtk95UwvEI6A7pE3OhUJ61Rp/nAXOvqN5onzhQuQIVWmAkKuEm70j5r2vYGHjrjB
T0HmIQoBj59gTGoLaGVkxGuyKVG5eNHDuCNviB0txq9Rp/TH3zVMb76sHPhbgehPcNHJN/nGvG9I
RhASjO7aYt9+Yvkkgwmo9Sm0v36PhMKA02uz7f6CUE29/pqlZ4dBWirJeWf79my0sWzGcCMwvqtJ
tGR791jDJIJwU48almNAm4lOxH7DHhBA5J6nPoq90jTa6kgXnWgKKs6VftrMJB5TW1LiNIdlO+5T
k27m0umRPlPH6lgweX3T+fMEKgMTouV+IrbzEvlMh4t7KoNBhvny9XlzKZR5fNX7rKlaP5TVIFdF
dP/ULWzyNzIsNUEoeuUT8bhC3HC5TrRFE96cFXVHtx3f5vpg0SLvwYNt5fHmpxHONVR8M99rNwVM
HjD/FQ1G9GKDIYbzkBcmzyKSjfFyezJ93W+SHxEmBg46zWrPE7YBf0HPYkX9myQckTm/i+mWugnI
Yo/zbxFKuI6SNz3xrgwCRSmyy1Y40glqLafdyjwf3y1Ge3aNCUxrgRpUU69o6vGPeHTsfRVzUuV2
bHAY2E9QlWO8iOXMrPcuKmfptSN3ZTKKGp4lMjn8g/KqE0fQ8tDNZo5J9fFzBbQnJW6WpTY2Dd4m
s6ts8XvxteTyu94eQ/qYeL8Xg1clUwqtfoum+buCNdbBoglXSGtg0l1SMmUmq1gZjNbhU2MwXNVb
jKkq8mxHfzrs2WqdDQLpOR/03+uqysgPB1x3Il1+arru9GmcoZ+VJM5TFusnTINBjgNeBMUI9eFz
FPvf7DGL/dnKDKk880Y5oiPsCVVHVX7VoIQtuzLFolfDWUkR8Xj2a/yJ8nm7q28ZUvx1V7uSvvxO
g/NsBbr35O9Aw+OIoVb3KzNGxWuZu+aPdWJJTRlT/tc3/WTlxRNXJHqMQi1Uaf7Jbvr8cluFrmXH
YsK4Wb463vDWzRjNx9IBffDlPV7/qK1a+rewGNdGZpCZcnKDSVkDpwjKX0H94m5WogXQQxRALt/W
1K5c23vhJxkriN06fP0Hsy4jJUnU+zHKPNMfLYLJGSk2PviRBpdZsvpbFQMgfaNYgEk1oEv9+KXk
LqNV+pHITpMKntTWbiB55T0w7VE3ItAF/duLgfOx82TnS1MkihMAy3S+eDgB9liM26N/SNdW7hac
vS+ZmQmMvGeFAL2gUS07MQ+ZBBGpkwisUg5aKc2RTKmctb1M2eR+bYALb9PnZDWUugame7vGTfD2
mDgOiwKjqKIHoe3mL9ZcOoOb7oy8ZRzGCo73s9RgX6LUt7YgOmhVGnlcvAzacjCPmnddEkA6SGeb
VHRrNaomJMJYDntxJjHK/Ho2CDj9l4FndIWq3VH7QMMObbJRwLnngzjXJEfqk70zE+KjPDu62cLr
WgpuygL5AYVq0jZbqI04C7gfGoUvrlZ0nGHTS0EG4wYOpRNIHy8h6ry+F4bnZcvf7cOwWXnLGcII
M4ZPR0sNUvHDzR3J8vIyl2n4tid6g5rCbDU+scE170Hz3b7SVUCWLmeU0mvbNtNCZRGJE0EkBOH2
obWGCWIv2mTTFaYX3zGh1YvTOEThNaG7Gn00+I02AmI40SWf8iS+ld8kBW0am8JMI3OLEP9433hG
XOpVWPBmgtmYNczrLpRzPVnVTgUItioTxQnBBBf8imFODG6/FNcB/n8AeyS37q252yUryFo0Yg7j
U5UcTHES0jJoT+J/atGtSnxITb1IL8eV83UN/GHnC8bh0am+wFc0km5w+kiA9oxGWTGOR6Cy5ChH
cgpjrXuczDbjwoyQSd2SDTc2y0uqH49tvmbetP9zg8WTJUn/1Hk/Dpj/Ca1N5RCUkdA5r/yniKWJ
jpBC2ypqlTecCwjAQ7fJFMWMsGxcGq/cZgLrahSHP75l0LuGhg/WNmVYAA+T2DOapaKzjdi/uNpr
gIqk9N6EX4lWwUm0uuJr0QnaId4lgk6ICagAS6XHGtjfKgcHl2XOpMGyiG7coQTOc9JPTr/NST97
Byi3PXtt87BR7rUMRIeh9CLU/VhstKqbJVpnQb1C01mQG1DSM0YKTHPdhmoei1W/lYWjslVeQhE3
s8dH9RL8kEn4sEWqhv11wSAV4DIFWkORUUSf/vsdA22e2FwcrB4JxuAivSZxJH6xTN4OB3xOYFPn
8Fr2sQwQf4At+TwhNic7/F1LHVVf08baFNDVmOcVO138QLgRfzOXqJ2S/eP2P2VF1r5anIZ9JBXH
AipniQr9Uaub1g1WewkAG3IMcqsFJ72+XuC+RsLN4BxpTGrSk7CYKTFccWQh73y806VtoKHZNH9H
1lDsxagEiqfi+yK8sEnDXxc3Ll5ms1rEZG0QhRdbt/cNJkTFKrg3ZyYQVXAxfsZ2DTpOfdO231fO
9ZIQ9TY+LBA+owIfKj29EedsLh9IG54Ns8OPsjj+RWBvZAAhDYN87dI7AbOnY10Mo1J4EV5DdqKY
7VmgVP88BCUNRvXym1kWd22WMHd04Jbvb5QmxLbOS8PDTx3nbZCPMWPQpNIGajm2KMyHyMF2h+T3
aaj1OV/Z8Jd+mH6GraVPByfxtt/AFgtQnCBzrHW/+pdCoaLHDHo47jZgGkSQHFtLzebyIcrA3qLh
msS3XZsJY0Gztfh4qQ7hsIIC0+jKP/259SvwMFWOjtV5NqvaOks5P6QwYwJpILRDjTHP/nfWxDng
OT9sqCemQhEuoXz7XaEo0/HvL1ACEzzFUUP2RvZiL5rB7ku5O6eVdQ/LVQ6bHBAesD+1zfgCSQki
y+zaGwJR+BnkyLOI+y/DcL/FTUqUFl2eNU/q/ToFQfDALa8EwKsODByNJLvPWUmA90+CL2NK3T1B
MDabsGbz3GV+xveW1K8UYgaf7SjJgLVYkFKjssUoMXl0YB4CPvsMnjTE9HSAlNJvTZHUvDjvXskF
tyUi2O1hXENLvqf+7jQ8aPqae0X+rPLfhEUNXgXt+MEi+s0TwIOswRbB6sC6IGYw/BWXbC9C+MGb
1yn4u4EwUfX8t+NVQx80kStD7OGKOfvYnJX+1z1RbGq1ZNSExR2gF7LZU/v8w1KbRZPnsm92XiJh
1BWJqACa7EBQKZhsBUR7dkO1oLkn6h2iMg9eJbDRNE0rWLgBoUL9SHKErwfY12LY3o55Xhs5l/WP
mplm6UsdQZNSv/1Gs0PnfMZ4fwbKybr4ofaPDUG0dSgLDTqq+ZTRF1QVOrVRDdX/D96qZ51ijhcw
5InkFvSR7OzuFKvpL0+1KWVaGfbbWQHS8UHj2F5zkxo+0t9/Auqu5tWJO2GzhpiF2+AvNxSCJ19g
N1/cV2PsTnCxfqIhvEcgffedQoDeLZQxd2GCI49dBr3xBsXTNeW75BbkLeokI9TaQOo6e84lZQw0
ZFDKNapE6BVPb7kRPCIiGM1DirKHuVvRGTg9P0rwWqmpJcgiLZre0n1YIu/7O/Q21kSe4MhjkUR0
NA926gxSLPW/QRI1RmsNw6Rkeo45NQneycQhoIorbHtSuRJNDTNDGBf4m5xPkaJVqpKRUgzKhITi
SIkosSxMcwlFbLm59kYEoDpkdhYRwIi5OjZBIcmKTlWxndZ32UBWX6CmBAJYeRqyWsL/TR6DWRI+
7QfyVQU4jBx+QhNxrUqdQdldG5Z2NLBPTlfRVQkhAlQCcDidNIYrFfdX6FC/TLajaB9Z3/OpHKDC
MfanzTNap4RJcBTAZfzXvDITqpe+K5rQnwAGDcp9clf0CYRoh9iWrIa8F46ux0q92plQXjRgxaXW
vPCJXtR3Nt67dJznQsgTutV3CSRMoxkHs2xA518mRDhu2+7srqfYJUaEToJxar3EKZcf66zOtGL6
dyb3x6H5B0t+VCsHTXhrOI7tYz4YtC91i6Q6MnP0dVvIbBGrWqH+rJKafc+hPQxRd4NQ8ziA0qp+
zU3htQkRvkEgZKLOKAgsTgA1zPZBuy0EtoKyaUAFfGDVY93I5leKD4kdAc3bD0mOuHmy0kbrmsQh
ibSKKd9gXbgydrLfcEKr89wbyKPviNk1aXTqv4wYjKe/ymXw8tDSoK9bLtLAivqWhxs0jOrV623H
8vtB69E0d0lyQ2o1oGX7eO4tIBvu4v+YtvJh3vNkav/oFOH7uOqjkAewCTP0TCC6k7OgDJjrd5Yr
xPhsa2/MsmBjY5xuXbT/3LZNSugtlSZhsF/nW5X/b+o5mzgk3xs0LbWan9hww2XlbF066UqWtXzi
E5fYhZKea73rFqJBIFhc9gTJP/mjy4127BWbSYiEnLqN/BDed9yjXbBaCXUBmaMoRyMkdHU5rqfS
VsxfmSZZTeVBg8NHGMlur/5K3J3g133X9zu1bBtxclFx3eTZo2vpH89NMLsaI5TLVUaOyQew9iXR
GXMEUp/e4PElfLuGf7jD5NuGU/H5vfCONACtvKOnq9BGnTM7SlVpPF1b/Nz2LoA5Y4ePSfbRGWGF
cd/SLNwIBNypl0t+UQQ7sekWn6zqP0W0jIxJJGqNZHITdeRaC2jmyrG/5B4D7dgpOvaValra4sar
yHOcfGMx/o6hKeopCokItYwJmwaSri5dnF3oHD49XsbRvipdqKXptyufcuBZS9fAGfgdgPC63bu/
ziGuDJnuPqN8Oryu/Bo731K6fh8IRRGJEV3TyRgKEYn1tD2FLFvbNqMyYaBwzShNsobAcgJ2CeVh
F65zpKvQnFFpSw9AvW8ihli3oosjV0s3EAm3t0wsIshAhadtpq9C81mi9g7NouDQ4u1UFADQkHq/
II0z62aAkgwGOfoIksoohLXdzvZEfKrrdK6+UiAVfnuTRXrbuVPpUtvBryu85hjZn2Mr0nbIZlJN
llbbrLkDUhUht/WDEbN/6zFwn6i0Dkk7K+a0EPHbOy0wfTQbyES7+36xFPW0vFlffWVLUlGj4OVK
7DTXNJ6vvAXUwZBfzwDQhxdoxGQWpMi+Tt29KubXIrbeSv7L6ds9pMIKH2XXsj07+sEd/szA9MOW
ltHOn2CodenRXRtCk060gewzgOuEo4/S6wWcw/sjVUIb0NvRNCAmruyzTAU8g+EmxfUXvFCOiaat
gUZHfsaa0ygcKKLHEmMevvZs8xLDZW/QzZR+XX169LoUevd93CHO7PZCmduSUTXf+j1oxY6z3nqg
ozc2WsbH9npCwkcAN6hIGW4S6BiJRcSEJU68RzWJzfb8e0hD5zRh4eAwYtgAXgmbRpatwWH67OmB
AeAer5hezpsBGKco1bJrjbYO5rRKqG3unTSYBhDAWG8wMFwGTdGQPYqSIR5A08TOib1MW6TF5QIY
Q1vgOaJvJRlnPjSAY5K52l4x3o5cEJ72xG3KeIyYKMfzVlN/9NT78IWql2awvaKtF25XUJCBe8Zq
tQRx++sf4NCG2t8KS/NQ8e9Soz8/NWv4RTE95CMoEIQd6TrYWa53ESCH7ihhcW+owq7SBH7w/pmV
u2mxpuB3YF0/eyWR/N5zf3QHF6Yt9mtFO9xyyQVKqzgTxo/Dv97au3QIO9qxlL6Hd2+kIbXkW82T
/uVo04Hcs4CiWnEUMD3qTy0sv82Ae3W8cF+JcVOjpDBw8TVWERF8v4BbdjzRhxAZg1oH9sDhq0oL
XS/muGrMuA1gispjZrGZpFTgR9mKO784s05C+6zWDHkrfE39dafgVAlmlcFi8IUYcXeLwIC3UYGR
MRmVYfpK9sE+3AEbLKOitYD2n++2AKUrUVzEDFC0UcgZwfUv7jfxYFz12qCFs7d9r4/M8pcQc07V
dFa7/RnHOVnynY8S3iYBdhnJy/fXwI0ER8jo5yMaWFkX0kUsc70BH19Y7/roxrMS92G8AC8Sc8JJ
rLiKSc+EtR0Kq9w53g4pZ9oRuKnHOnvd+z3gk5ApqHJB1FUnAl8vxnhUlyGEjkVSJt1YZ+gzW/1m
yj3tSLG9RTIEPdmtQHx3DsjCDgH/xGxgkyXNE8+4c1wctXhVIogE6bDUxaftiolc76sdoM21lS7S
SkbsJqwq5pPNuyDZuSUzw48rmqaGv7zmHH/epV6695u5SZMLzFuKQU/BkgzanlAL4lynfY1stTYv
z3g8vfYJWg0fRAyrbAbrX+V2aOxt5qTVJ3SUCXih48TffqNhpqUXBoQ5maZ0IaVPnc+fxKG8U3h/
Y0SXdVhgNjLhjYh/I9smFP0tcn45wUYxRSkRTnczro/aG1Sm3O3cxX2inzeLIo/m8XOpwRj0dC5+
B/WxFG2HLRVkQF8v1fqDNjVULKNQ7tLb0vGWevBO4j7v3pK6IdViAs/ZfmKdIw8qXbFzeGXjzwJL
VILFs3TPBf35Jtpyt7wcWrkrZeQf4Xaq7GTG91IPDIklKOMt/vrsowdWpedseExx+UJVYOqgHPZO
3qqfMGkIZWzGcVYT61Bs7hmHVvG8CCZqrauGNJErqXzShKrEZhLB68j6ccMBiScO2wRKpX6kE7OW
is6mIE7D1He65ddgIRXsYLD00sdKPB4Ra183Ja3bcVQOxQ+BgMgwuYJ0QAe04L5J/9V9EustTUmC
k9arRCiUmDJkl7qHrgcJqYkHC6O+68l3thupbLq9vbLDGhfU0updEJyJsBoIW8rE6mK+QfcOnab4
WWJ+OsexkZPXyhfvjrmgIm1kuSurN9+/1BJkT5QN704RyGsGcDtz202SrGP3QztqQh1DllMJ9Pp1
b2aZQSnGrWBZGPUZrPZAgfxfTmEcejmJBL0m/bukhLWrelvIqFK6gEqqvbJRauTse9zxXcwG9sYm
DV7SVx6LOEs0LDU1mHdVgxmKMXrq5bNdITN8c92FAGqW4u8Q+YV60MbEtqP5AIeLJ6qoL5XQDze+
vQ9ZRLIOOEF+TS2RpULPY4FfLkZdAdHSPVM6a5Ku4U+KMVOL6Eg3NV8ge2cWWi3pv3kx++jmqw5r
r/y99iQ4jrPvq4QQDGv9sq1Ea5eobXj5YS0QlX0WCX9EdwH8QDrU4ABTqW24W+k1esXzj2eyRMPM
4svwc+ZHTKJ5W9E4zi+NoKu5kUWE5uIP8nWaKctfgr6MQeqinFFoZjnSCpmK5wwQkYm7pe19HSoF
FBzS6+bed5upCdw+PmYyNWXX3D3WvwZKds6Pdth6Rrby+7R/zt6Rd5YcBU8I72k1IGMPhoLwfPIc
l6Znufbv5A/65sfCxikF0/wFRzuNtninmiKRy39lqEugnd/e/NxOrkbDLTJg0Ca999ggc58KYT2O
UOattf4ploGEn+tmw/nwYp62A5JKQcKNLdbMsiEIp3cpG9Its68tFknxJ4th5waS3f5Qw89OKETh
0Mb6GiSnGdDyMgMuwxawyjWuzIofliVCq2HwoGMwkR6TK5FttCakKPjCoykAefmh0v2AjlpG4Lfj
ltYHCNGhtlkmrFOlZje0+B2v+J2qaOC8snozpmDL5k5/5WXiI2vHzc7fYhQO9m2bXSC2ih6UGxKO
1wtkhOH/7ZToPrde80r6J7fY+4HoDUEJ9JLWjUjQkG5M4vejK/2kSJdrNLrl1IYbU5mBE7ImzEFb
5OJsE+tvLdkyn/okwy6zlLWc4MrFGl7t5bny6wjJTs99z/IrP10MvwifAzOmwVkgkHZgbE+c0biz
UXx3kyvbCuAHQsPvzr7dOg5LL/IZCkvSvfcmWH99pQ3V5pEKP4o5gWyeFFpgxhFwbDdNKkSOg+Yz
KIwJtR040qC/vxyu+LtkgQsHNRYvctxFejlHEK67pNdP9OQ0HugF+xrpDu6yLpWkeXrFrv7ElWqL
22uJsP95yKNlDazMrETkZZJtK5HDUVYNs1UEfqskoyCB3qM9+PZcTFXzZ6XIbian53XC/xFwWQjj
S0E2WCNs1VVBhPMM5ca5SjtxdpMhfwJOwYyTk5UjD5L814AWq/RkZrnPPxe1/YBv2Qex7U8JizsC
jBra0WREmwZb2Mn9+Qk3HdXf3gimVbtlSTd6w+6d7jE3oayRB5lWmh0LVyTxt9rHczg6SW5Yxnmo
zkvWmAv/efdH0wewDfkWsqxPmOHClLVJbmW6Ur0I7u0GR5B4lSmYC5YwBonfXLaK27YJpJ2/1qPv
tmn7t8r+xn2ukunfem3vnMHpSGaCegqBPJv32rw5GofmzhtiDqXLCL24J+OfOrkCzdPyD/9NZG5o
2taDRIAMGWGwV9t8yZxa6fidNVdk5xzCG/V12op3LOqVV/TyLtERuUILkfKM0KRWKiRuhpyAvWOd
HGopEkcHGu2HZZEOF0dTesnvgM424/u1d9YK5CUWULip9z7Aor7Sf4BAMxpdU/pM85rupUNfmx1u
kKIk4FRp09v/DIoVNVW9IJB5seyBSgUVF+6NasBILKr3YyTNQlX+w4k11tY6cuRujmjFaEBY4zp4
Ub4ilkHLJDMQ5hhlm1ky7iBakgC3Tez7qIH6EeiVXw1WBBUF/UdFYYWnRPGGEud020lKnmdyzyfu
/vTJxGiGl/xFK3STwQ01kzxV9aixXCA/Fzka6grrTtfo2ax4wEC9SVli6kXEcv5PTh+fTh8d5l0i
37vTPah8X/I8QjjXnVx1TryRpQ8UYO/OxN7fMy9YD7HzAvlEE0q7aVJYoCkrksu/rKwODC0ygTIC
3o88hYScxseuPY/qb7V3Rx/uIvry7adtNM2yHMDliIyU+AdqaygqpZ/mc58UIE0Nb6/dbMVeUoYk
GyxakCiPGCs0LiknTB/+vrr7/CLJ6tyNP+4gtp2vkH/uPUgHebjcBtUHRG7C9jCKEbxEitMxgvDs
tjmLfDbZYEgiFrat1xITFaJrMCmVNqqSKx93i8o0dE1yqlFsIRcPUYQruPnaKyA2JtxeJhFqWlR0
FJ8CnWDUXYsdVcmK4PC6mX/a3TdZk6cSrYkHyhLiopHHKSUi+yYY7vqCSkeOzj+6GSBnc1UQTLpk
as+m95XQS4Uaa5Hm+8gxkUOrlKA2vf8EjXegixadMoyiuT3AxWHDFMOEMuWANMiUV1YA4Cc2NdZY
t8qJQRzIIuzkZcw/hMYkAb4DXCnhNSZN807Y4Iq7wPbJwp43IbUeL5uZNBQINiEIIEGsKhOZz2ym
zcuDS6wEfQRYtcLyDAHtRnepAzVIa/cpDqer3DRpjbJpM8vA35eppnmx3alJytAdeHeE0WQf2Px9
w9wFctfJvLocvoL3b63zx04l/5yQZF7UoPlJXhVBYrmRK7wPpWdSEOqE9FxgTCR1xkd53IOnfWaY
hYPQhJ6fpjk0QYFPdTtchLj56JC+qNYNqwICn7cOHT4ejm3Q7eXn6qcjCEnPkvTbPnv+PrWpTQoy
iEPV/tPZgtorM7TLwExTh1TLouCU2nGP77AwsUCzLrT9kkwAf8Iy/jixo0QlqcVwjuISI8k+dq1E
t1o0bpf9dA+YBdQxBUt3vuU73+KRlSG4oKLoZC2jDbAcupC91Tb9yvTdbY0UPzMPiMa8ievr82mH
iZfUT9DLBri60mrz+SYZf9HizoNDiwlHpMUVmEhrfcRgeZZ1F4AVrGT4cAl7l2Rj/KXCp4i/OhVT
ovk8Z8tyKNUyfF54yScYP9qJUqgg/L0ZqrolEzTW8QtGp/CJ6zEuoJg9VrY3+hMj1l+1t6UyQ8Oj
x2MRwKA57RtTAFHuW4Da0NnKTBdZauK5l1aiwir/PjbxYuYx4xpYvnvuNyq3wbMXiIeKJkZLEuxn
sImItsPU8j3mETzQEYS5sQIDxOnkH6CJW3GtffMFiOsbxcsCvxYnwIKuY+5p/dlUTvgElM0dWaie
orev73D+q1Alb0yhGXdkEXrmxvCrWfPxX6v1gc3aRUQU7ZSe/6/O3mDv9a8A5nN0NWVWFrHm5MIJ
7q42TLaHoXDfmCqbv/Xg0v2oP4s1MD3iPKCO++ELzupXYJsU0ysRiGlyxtQr0aTgNnGgEo0TAdF4
Hpf5HeK1txiNuPkRNMqw2vHlgvKxg9kGIhh57bqAKwbzKU5xxYx+TWOvvwwQz/k8dos5/Qno7MGe
J9VIy57fZR4jLBWt0fVesGsISBMVyIBIjVmPWcpJkVHmfGsgRhlwN9gN9yfHZY6H+JXXsKPfu8lh
1k7JlI6a43iD400EvalbgURlwd3jcVBOYCTXRrBCiMFqFVaDLG82PE4H1I0hFWJWkoAKRC3uT0k3
zs6OrNlYexUcEqtPab7mfqVDSTGTpvYAZgikSR31TkKbI3EbFJ8L/CxIsdvdE5Jll4XXEtsvV0Cz
5e3A9phoGTJzKMwP0h7HV+8c/CvNMi09zC6xIDrfUW5T0A3RPNk587OQS0a38pd925AFq/bEwIYW
OKKj0i1RquQqjVP98XxyEzUnosDrlPGVPeuf4U9V5muOfbifXCbhhCdIDalqo3qtzz+nFoIH5QIA
KkoiAqua/Dn6yWf7KgYZbbXgiLtAqsviPPx4wPkVg0j5cJUvRgcD44brpOy7d9evwamjqSbGo5zb
n07woqbUrjbQnZ0O+p5j89tgEFk9yVrxl1NKYQfFGPEiHskG2xLVdpQKespGv3k0mNTrLdj/ozpH
/fRe/0myKkRkVLBHuGHgD0lGyi5SKetlF3mQS/RzXY7jAIzbjw9pOdS7UvdbjU6VTSklQhuZyXnR
5R95CpgwqxMBDeyQZxgdlrZpPfTe0uzAlp2NleF0fMpbEcOmDK4/6ekQ61MyRhZUvSsliSPnOrHN
+v5J4eWMd2hrSDorROvvWyXsx3VWngTH4VarPR/jRpL/RUV4g2DWkE00BZ1sKWvk3K90DoYun7ra
HXHI4dDGSN+56/5UGH2MuAvAPYMYj7Znl3BsjvtY4KzUKE8vcKWInnVx0bHOV8YdJYgf1NvYYlag
k9yeu9Olj3/2c7K/4I4Wkdg3T2euVbfuR9OQfkPtE0aGrJenZPiR/Ifr3dyxPTLG8VsZ7EDc19xH
wwYFNu9NuTVu7EMdUeon+c5P7S/RNEBX5vYRdvAVgYGlzWKuFLCdRiIthPqe0sDfUHFyuE4jjjcK
NJoie6W1PwxBbPdqhfhm/CCUlSoo1nNOxIUH0PpC8JLH/TMaujWmCObdNEK5DtA1RtH1S2/BLQky
gVM4lvKrdhj37sGi0VoeHdNicIqB9e14NmzD7mnfo9hRdIC9R53/YjDw4Rf3sy/OuCWVhc8+rdWX
Nm8KbafgEH75sg6+RfUXwRKe4GHKMMZf/HSbhun4K3gP8zxwZHpG/gSvvRNofNucH/ygeSaX9iL7
qQirYcCxy5bHlbYX4jhBYOldwu5FYxp8hHgJ7g5tZlItH40mFRLVfMB4+94ydtHYQ7jL88iPtu4+
bO2WnAyfnwfNN8o8lDX46HELTUPJ/G/wRn87k6OqLuOK2+kHLYC7PP4amzAxQGfusYmJH0lu+kpM
gTH8iMjsY5QyxmyLuFRk55yfxhksZZxTtIqEDZYZoR6GyiPOwS5VsupOIouq0xgPobWI6E12Iv+x
q/rxceE+fBskg8EVobLAZEKw/+crxKBsnjIGtGIm50QYn5cijAEAH7ixS4DOT5IXYCrQ1GCPHxZ0
eBPJ/31Vm/cLGT9KMTYgrV61qd2wz3KHs/OdDaT61Y4RinTQ2seJ3UdHnSkZJ7KfLJZSw9tuJPYG
OpalPswq/CmAuuEPexa0ARO07Iij8fEEvoeLO9ekfqG1qiJeMTGNFDrljw+zjAnnlBKXMkQ3VS7Z
ZP7UAHufFqNXu1qNYgh1C82nyOO7Qdmr9yAQWV1/TviUFMA45aXrv4su2OPVOC9OwQgDN70rja6t
V+T6/8e5etP6ZXPl/ioKO1DQlEqRszaINk7l1Q2C99EZEbi6xXudirySCf1p3g9IhstKrbZP6g9V
76R6erHt0AzYxeUrv5yRUJq/h60sP3Mz0DhIcL4VW4Y778cSQZpX/dM75unii0xsOgzMLjSAHykH
aLOToq+tar35bu2MkqcLVrDtE3ory4luNb4jG4f/q3V5R2hDVadi+6E4cCAXwKVz866w2rHAKtwh
GyBnYWiZ2ord4vsOgtefpspjhDRJrVpxmJODKdTHPa4NUovvPBY+/R36DCj7DAa/5mUBe5jtuYvb
Nt0lpmdZzV5dCPGqNTuVxfKG+VbGRQDTF9R5CskufCMEV1kvMlYtyeIheGSaXicvlPrKpuLpE73T
wF9LQfbcfkGxmgtyGuY45xpJSVjIaqFdAtUcItR8/W3OCX8ugQCcMiXR8sZpCZ39WQHjTz5QE1sY
OmTn/cNQQ0MIsbsmwP+iX1L4W3Pb13EZfbdoUD9Xh9ZKNdMHasz7NCrmGPzSd2fHUvsU858ve1fH
8BMOvizWAJD8b38SxI6UaHaY2dlNjVnhDXJ5ogzCFlKZfN3L4ZpLwIrZ74B7DBQ+2/y7bmNLirbQ
Fpoq7V6JAZuGFOCXnT2rhR+4ZjcKLxMOd+9GV7oI6AjaEZ6orUyKYFshLc616xkGkYlT6W/VfaWv
XMr71PgMjxOkRqJL2Yn/ZoodjYXRFkdH32VEBCoiSn9T91P2DXP86g1Kffa6moezJj7jnodsq0Eh
W1H3Q1fYKL07v8HjIupF/B5GOxYLkbDFBf+CQSTddfRWt3hXV4k9FSbeRIa6OFTvzMb5mimegbYa
uu5fiFa1c5Bm9g6Cnd7QKbDU0SG1pzuHi5eiFbWfxZIhC+dTZuvq0q1t9XSNit67J666uWblLX7Y
+ZXYelgrVpVwlDgdNQbjaAbORk+obIv3d6/5IB21C+SE8TltL02vp5SN0+DUjofJnPp+tiOUo+jV
No5gNT7jqPNFL4M+TpDojlLYIZSkHwvhlAPG2XG3QZQdk5yvIQmypd6NKT2v0Yut5zRqAa9TTyl8
KpVyMYDQ/SUjaCyv1Iy1MDXiByZZMJG6veqf5xseoZ36+zS2/2KuTe/9zc6o0kjA7HGoNA6WKgyA
/w5nk17A65ks950hvEqi4FzDlkaVQxPSsxdlTBefKyZyTx9vjV2clxHCm+iqJ5g4G+vCKQrS3FAM
bdsckc6PKhu8POR2KAUIxyGUL3xZ/QoEtWmd4hfyHHGwVy7V4ked9ELfym8vQnZv66Qb2rpCQc32
tspn2WCNlZjv49h8FaeQPz1ZgP8/ArPY2VLBeQHsgJ9I1XCaWarHaxb3cR5PORGwB7jM+1u3rLGW
SivBoEnUNDaoy1DKN+tb6u95h+H7cp58eKBDft3QxMfeuEI8qTSpojEeVdOgLGiT2i0I7vI49upB
WaNB23ySnYAqH03iJZcQXTSLIEesec4hR7obylx77C9NKMsBmfJObjHpFix0+BAWblZNxgvYwYBG
PacTE8mRo08Eo3al+ZkeYZ3n9qkeMAMMfk9B9Gbx/Mw6imsUwELNoO/bLEgTBzXZGPbPkHxglpPN
7zxGEA49guSOpSYAN5Y3121BIN+zhPv6U8SPpN4xpF6F5cypVKzgSMG/4oQNJYWR4pwGrv0kNuaK
tdba6nOaq50JJmO48li1r3j7DSqNLeIPe2BGqKbzGmGvg1EFq8VHDoKZAw2LJF1IEPXdcr/YjFJP
PWLwZIVOKVfb+p8sYBK4WiG72eK+HR3ndNr7l2rsihQn39YiSgI5FYN7cphBcMdMEiwbeyFDDnQY
dZxnCmNYT0HJ/s0iW1yFrkq4V9fcPTcQ8eY6aKlrJ0K+ksDsy5Ozcf2l0ZlRwP8halk+SKNkHBW2
X5VdPKxeZ4cG2p/jJEsVs1Kn8dFZ4MPd/retqoAcX6WrYyq+50nQ4mNJ17mA0tNq+0t3vJRNbqSO
CwmTZ+CQZ8JA0xgBbC3T0RIzR193RHjp2vUZSo/fjlGiHcfiQbrvSmfKuJ8F+PA/W2qk++S9M5fM
nK6YMFQ1DH4/zuRBLGf4GvtPD7wnAC/xs07MO2YXmaWJJc5Iw2Ixpgn5Ixb8BzgRmmZ0KAYin7fo
rtL4vsJfGD2QhouDflWnz4r5Wgw9NEGdHu5AdYDo5iCRdY+ZocZ3sOfTNJXxXkdwrgQzAql5elxW
ygcd9zZPl0b+6125NWkZruyMUaj6Rm8al4oXyCm5O1u7YXHxc87e+VVypj/H4xDG9G5YD3SbFbUB
9tjMOfHHFU3ZG7yNUO6YPbYSoq4Tlh+YQTPurbDq4zF88LtVoiQRA398DIvEAs7a4NJWRhQHwP9f
TQEjkm5UcXqwXAcFeTBK3iNBesrlfmvHQUJyRs+pNMmhsWvmMcDMwnUkCWxC+3WdFd2X6/V9LclV
OGPeBSGZmta25egdfr9ZNGe1DuN3zZyeATq3B16p9rjcUTu5Rp7s50FxyJl70QEP5BpN0MP6zeLK
DNO1COI1vdOcSKtaVHHCR3DyCy4F3xmVX32Y0/3EjQTsHWP/oUi4BQT1D4peOQWV5MN3flwdjFV/
Z4oFs1Dgg6E0O/S5EHNzUlaavRCaO3uzwFqaokCgVrjCLQT6BkGH9rzdCgm6kF9NaYBv9CUv8+Lw
IJywPVpDKvw+/IAc337U9morv14jPPRX7fu9T3Mr6jvNMLdhZuGSLZfrKb3BDwRCtQSF6azbj6mu
Yjllo/pfQI+BSySMp05vpjdCbP84uFTNfinO1i7GfnPggGjfIb+SnUdMhOSzxdvWFhfS+eI1TiwE
3/yQ1YtohlYS/m4y1BA2bJ3pzpudPQ89KDbbjurlx4N9L211lnZDX7Xr2inIEoDRh9a+sUhnLXBL
QWxXYCQ/aIxzBPFtolAWT+FuexIEyhJW+snXOCebwV7pHhe7Uf7CBf1WohnW5gyhlwbw+FC1ZjxP
S9rijMRuXwgbp4RCQ3oRK8B14LCX8qr40jycpMQbNyFTdi6acFvkqjJHGBluZbOttmvsQifJJUM2
DEWT6MJpzBWRl20UHuKrSEkN8eRotsAVk+qY0h7T8vTL7/Or+YqupF/uB84cfqlHP7I+DR01DEkE
J843EuEr91s2r5AcnOcaYxpFzbxXLZey2qNNL/wqXLI8YJbsUYyLVuXHTXIoXcZBSYIB3/TwznI6
waETDfXPznvkGFnN5UVfMrN4FVB9ghhixneTNyYwA/m2/3JJlGMY4N3IOhb5v/0K5IJqvdyYDOYn
qoZC3UMDo4sw86/vsxqEAMGLK4hlcb2dBCWhRIxzrVETKS+rHigH+v5zAlOf5mMBZlCdgbwnyTd2
kTp87y86X1u6S4jdjf+n9DuU/jh2AeeYQ/3MGg8XAEAWK/Ttiuwi1cztII6LneF6Umobg2tJLvYg
ZS2h3dMz7lE9xkburBy8u3wIzkuVvFB20vMFtW6pdDOWvHmbmmNsPHW1drxq28oemABZ3ZrvZ4UO
i65QtUDEzp0CHZVkZhZDEYepVRH3MKvvJNRHS21qx4p+gqpqacD5YoUsmLwe1AN/QsGrD0sV8Q+o
Mx6JnLhyTqx7ON2VqV8A1zKhBVEiNOOyOdt6UaxGZ/VCqmSRYuxHJCZ/re13HUVMl/Vq2oPjf82Q
FCefoQ5q65Ee1LIUgcz4jcZ/Xd9uRD5bTJrP5m4z2i/kK5qwCQzR/B+2jJf656oygOEb7vt5ikRC
/3vFOgZ1bVhTDVwPWzm9W8betWrxi6x/mlQruVotu7olpwTJA3yIIiWH1IK77LGsx2YIIc59ui4t
fOlSKqaFOVKTTEm5GFPoBRhUg+DPuJDQgpxfOTjAil62zl57+fSpB6KygPrtRJMK6rcc0DKD7OhQ
6D4UDQ+J3rcsYs14ZjzB36Zo8e0Xo82USMdcCbGFK9slQTMDft4y4j1emL26KNirVQBcteYNIASI
N+p2iYB3IRYUhZ+4JUG8iDNiOvZxXmIYr7NKrPvPpTT4JtkVfnsD6/KMCD1eqqFfjq1PedIu7yWa
OAi0WAACS1aLWwsw0V9WD+qtB55OQMQK6vcxrkB/zFmtDAB7hpaLBMo9r7qiOoO61PJ2EDzryv+o
UJuVnkw7jCqEHEIzgPSV4AWwRuRyYT/ZBCA4GZE1QTQsOwNpVS9Ch+PT7Gw2Wk8nsjNEmS1196nP
rVRmtlEi/nBpuPycGZu9X5C+bwc0qA1Q5dpmGiX8WbFL/4vaYo5+ecYMNAwIILcW2ogOLlE2oU91
naYbSn3GfRGGxlXdSRFXdSc+eCHjA4AV3bk29WMKX7bUjBEqgFVzeW0oK+8J6OkEj18//k/gEMzA
tNu4fsWe31CH2Msp+wh10p8GVJuQrgs+qRW4FOK31K0nBYJMqwCzsxkn7i9CTRIC2O5x7EozvL53
O7LOmmnDhxLu53K62YEzarrUAQkpuWEC9ILGNu6dSA010OaAQ9IFdAOPz3n1CJ2ggh/6fgM663zt
o//3c/tbEvxici5t8NryYHFUqpjPr0ehOKCASo4+yyKmnUHPf+T21CVZOg8OzUTQyKnyKs2JM822
i0Vsc71ArNRCqhX3JaOvg3f6w43MDDccZk3/x+rHFUATlTJB7wKyHnGbMZ3JqU4AeD16J864Qz0P
O8LocglD4NSIwjaFq5A3rIUWlRgIiW0TufJ0ypCX8TAOk2Tq2wn1qr2oKnTDdSAB3w8epubD3uIX
VeodXiP9l8Vr527WEay+oE8bPWTNAuw8gICXBvHVTN9J2dYgXeT2CocuZ25m4DGkmMOs/JfYlj9s
Z2PRchps5MzzMFz5iSY/XJvvwoV15lPQkJXh2Pu0bbUmKVsEb2m+TWLkcaYDxLvRpyNcZsnDHWJE
x/33ZDfdXQHpm5wdHUdMyVeNxqCiGrklwzPYZ2H9XRjOy8yKTz5AIt0v/x/bReLQkqTwdWy9OGRf
q99X7eD7FHAuqB0356m98wU48c2DIwEvm4C5o/MSiWx70k8CgVGPtZQoaUmmG8Ctv6QFnVar74+T
lFWDuDkWstfF/GtjW0c/cEwr2qGtA8chs/bUBDYy20/f7Nk+M3qm8L4W01jDXj8cjt8jaGFV/v7y
LZ8Xc6HEdyBmRL/fzLGkKGrf1Q0vPOaBIT2pXBhQhm9beAHPBmjsLOFe37RnA2mnuv49nWYH7nXb
nOof+w7i+mx6C4d/EJV2XkXTZWe3mbH08Fk3/UfNB+gug3Xvm+QJPiPdDKayiYwijs7UC/Marxr/
tUjvRL2zN4xP/TI1JBgUWKNhc3lN2JPwPg6Mf/BS9EEt9EDk6J5pMCT3b6jFSLW0AFZ7IuEOyA5l
HkxuYaJZ5S7RDNo5z1f/WhOOZ+1mFzdrT4dD4hJ2Hn7XnkcUVJ3zG/HJFVGoYhJhYfdZTkr4C4/T
s020B/I2SasLqEZOaiss3sESI/1WZxP1aD6VuVCFS17XcSQnzhNXCiJ1222fNPVE3OYm543kEWID
BEI5u6NrmeAxnZWxDJZ0kMN3uEDQxCBKinrx5l4XlSvhMgbkQmSfp5evZ9F5Soh2LYMS4kByQuWb
d1NbEc/E12CVWoN/qH3aNAyzoQWjqW21DKALdZlJom0y3Np5EQOKuS700cdabw/nYPY7CZac4Mk/
HetShbUB6/gupQFSUVVyjvTmt98g46AlMeOxmFRDfWntVjPBFeDQSm40nzk/pZ950ZExVCuViosk
tcQjziRzJ0GCudw25G6541SRu/pCRpW8s9kz/RuERGkIyb82nmTH8jw9bw3FaV6hUuHvmcKD9kXh
1SeDmf5Ulkfb0BUtRhDA1VkKevr5tz0B4Rcsuzg1zV9E3m0LRR3CKxgscgJbIDNyfkW1MowKh67i
88p4e10hiFY/QhD+dhSo8ZD8tQ4n+8hTTIM7XVF8w6WPTatjTrBN5FkF7oeZFtfJbrCblg1Pl+RS
zLh0UF4k93qXiz1bJ0XBaGRqSXRLqY2kkmCvM31FCv51B0h4IP/OUla0lIltIIqEd1KpzYwtxCev
r/RR4NbDnvBxZTu6tvHiAgcYdLyUqK+SRxbpjWIx/NdmNwg1zgPzo6NHiBfF55b7xBAYnTdgH4yb
uieyZhC/STha6ghMzPWIj6hWmc9nhUaEZOvv+CAAj6Y+9bmGBB/Afi83HprGxZcr4nRtJ0R7sqUR
RjUOkO7Pdvx59T5DNUfaA49ekMhwFDfH7IUTMuY9fSCOoGQI5zQDbqwinpQFzZazggJp1LUH/tJz
3XYxb5jTBSd570sINx3EbmuSTr9aRfJpiPFy5xNFsXbRjaghTDhoky7vQwxFBaVs3EW8jTQjZYNf
6ohZ5CyTIiguHPv78iBky97TB8PCnc1EU7avBaf9+7aSn6R2QM1X1kXJtEOTWw5Sv0dQJ8kRPamW
Yl74HljExJq1ZwYNWtq3PKrLwPXobbb6dNliTnNivuDYiZgqKxrsdWNQn3rYlz4E1bRpyPiHNy92
MceWxRsOhrLQAmgcWLYWQ/dfGiUZLY8KTXHYcwr7x4yYuTcnnMlXWKtuHDB0euCYnlxZvSKOH/S6
2/PpKiOP0a766D/ND5Ynmavck/7ya/53ZX+WT2UqLGW1G7yaRT0Y4FvMWtLjgpz5aIGOtZK01CsH
mExJ9L5sbUxXd9CdRsoDiUifBjhgrTjy2e4I47DXCO7e9MjAos5qTBxDIwI8+IytPy7qH2q+C8eg
AnGkg+HrzjeXre5klzykYEcDcZ7s8oQjbwD6moB59rh/3i9AfarnVN/8u3bGC0RaBca5J/w2jDfS
YZMa4/21145XEmO41pF6vi9mFeDMh9e/ETGisMCERkzKCycZtirM1Dry0ZnygaFWDime3Vt9BXs0
D5Dvj7+zA2VbQ371JZ/AMBGu8HwFfApXhFaaTCRt6ttR+vh9UAIWDd9GYNkX+HfKLoWeSverHxWg
FblgFkpa/H0cNEKFVUcKIqic6EIfDB2Wyq6Z/SQE/1z/Y4L/CeG/g+WwnMXlLPs/m+8u4XT3dp64
EFS/ZGlB+Aa84qmn4SchKTmmEhiLnX4jI7LgOL0M/wQuJ7PkQv04h3uw+dN47xSGR0AqHt8dUjdL
XZytxocE3LUNfvIP7/fjqcERL39qdwr0NI9woJNswCuYr9MMXKeTya2sTKA+O8Ve9f+Lh6uY9iYT
+iDq3cy0T6gpR9Io2y88j+zfPmUku7exkJcz36r7JTL7IFOQ+pq8vt48BMZkTiVbXDkaSrnyzqRb
y8VkJ4kBUm85/nDlW/OgWxv6VtPH09xOh7C3ANCOkSj+8cnYgmrO14RmkIy8zX/f5G7VU9vli5Hk
xex4p0K/LPfrtuQIuw/+/zsNMT9FHVSGzUdwMcPe09RyjsjSFxSwe529kSvH7PEnSsE/Gds2P6Bw
S6eQP2n+rMmblX2oenkCrpNnz1TqbmK4El69CVvMA5o8KjD9AfjRy9JuDSkEGYJpubQHa9xLpJk8
MasDJhttC5X+OPEaSFymcrDrMbZ2xSWe8OznMpjBKqewaxnHVZHlKpjJEBYSg+zgIXu+4qh55UHT
cDQOeKjk83lQSpN9hSfcK4oNfGQ05iVQBTt53t4yyz1GwOyzOPn8pHxC+2yp4nxpBcLggX1J65FO
qX1ghunH+L3wUAdcJBP5Z2memrCkEz5oQslKOXHa6aZKbRDeqty8JCwGrFUO4LzJfQd3+9Up1UHv
aZtBbLoTfUvYKNmC60Cu3MfV/z54Hr5OMFx43Xow5DjS7ZDxmbnW9gxwkMPD2VAsFiG8D9c7IIiA
wPkuRixYiqOKeKZgjDuRcEa79a580lxX4O1M9Lktzqx4cBN6h7fs7x2s0bcpmq7b274pNN7PTA52
lr74ckVO3iBUTcCIZgDe0q5krFGfqsolpnMOQYvDMIUN1+KCbR8gI0MTOJXjxw/+91TvEtWJYPBy
jDTBzsJ/25VY+9Y3eXAUC7r1kLvJQCRaP9SezxpdnYgItFSqD89ZZ9I4SEYRzEqbyCNzawM1jxf9
/GCILqp+7v0vGHrQauec7WVVKSKsxmMtLgRgeluMT1V9pv6neyHzCVuzz2v0cV0+5xuwk9fzURnk
dY15jqcGe3yxUw5AvqWJWozdivLeayRRKm0fPI47Pzm9MMGglDpsYhE4PdUjhjm6wlGsG5A9+XCZ
gnclW0rGH6j2jnlLp6iA+MLtSCQv80lCi/KBfPYO1L6+uq1L1r+5uYsfd2SmaWnfj2nc522TedZZ
5uY2HBEYI8hl7A+U3La4zsxo5g6ALTTSN2umKQGqpd6S95FlZaqevZJ1OCSZUfMC8qV0tR+rxp7c
NjmnzslV3A26gJfK40fa7pYehfdoiQ4G8nmQtbm843PoPoE6ZqevSIjoTbtw1zGFWgorJ3c3jpfW
5VrtUkIM9Lv+QYLIafoG5Ds6lY7bncayFSzUe5v0OVyV6xhF3NiH7ut2ECqg0kzF1r4ED+LNcdni
uw886UKFqvbZkg2DGyMJqc+22y7k5Rj942p0e457e/U1xrQ86Bm+evxWq9OlC18dX0LlvwYMT3ZF
/kqnvVNnCClI+yNVS2O9mwNG9jAJwb4/UHt5g2c4EaqJLGOU1GZhHf63dKfPuiG27KMUzi8fm9Yh
DN/1/hCOXBZl8q+HdQXdAaOW48vNoDST8DC3Xf1fRX7TFP4cLLxV3xwO8wvM/UpOylkWyZVRi2w1
GhEfP61NqiS9GCWP3rKGiRzEx4DwPNjVUMmqZpRmmDcv3CjUNImCIueCfQOfIN7qyUVSrvYM77Kn
+4+fIi0wfeGN4B5DVTWxicgzPqvJx8F+JJ9nm02K2mYx7NG9xhB8hCRhXOSVDdTl8lfLtnVE8aSH
aMMIuGPqzhvJVB/Y3RWC6rj6SlOkYKEach76tNtvvhMRtcfVkiGcLVgviR4XKd8lpDcsHfyvISJ6
2nNzEJ7ahyiwdh4bZjtn9IMhADdXmEhS9QTYYARa8AN9S6R8sR2r3fjmNr7r8y10WEMe56P9qDqL
rGJQrfxKe94VXLN5PL83YsK19fyUEcVfquSNZ0AIFqXVtLcHDf7qad+yXbYVzGbjp8i8pRlxDKfH
w5IQWqJNdXrN7DEFusO4MX+He6wDJTjiARXBtkW/Ha7NSmLcIF0VBXLQZZlxx5ee1YVP+GyPSMLN
upR5Wn+QYazs+/elve2BukKNgxMLWUdITha0jLnPRPJo87V9vfhaPDMz6vj1oED+IrZv58TiIm4r
TxpkEffmzyTuK/tryZIe9pKWAHXnBY29Z6KPBJAQj7mASXa9R+U7YtD/7Hvx7hZJqqHi8niZ8Drc
ZMlbEbAl2sKqRz6k4MvkSiZ0fP8Y8JlOmsHVYEJKq8PrFm+D8aSKJRNCm7JlKifWa33pli/p+fZI
qVFFqFfpo6psRLQ7aCypQ8CIdtXGm05oIv5WE6p1r4Wqv+ytiGlrUweIprjfGwUX+zjGT3vA9euz
zmXi1lsX/veB8/v3lRPDj2+sKRPQkEc9aVHM8FqZLrS/Agyr72xKgED+Z6HY2WGKTYEpT/WBYyap
k7mxQOSN0v96vNk1lm7BiMKAu8QQKy7c1jBzGyxeOs7XLkqj4PnsjVEjnLR7xiRta+ZX/+LRRhlz
vfqRlhwubk+zvZvX2umLh4eiBAuEjCZZPtr5t75AqtgCRc4SG4Z7vHV13Z9EKoqCtW+HJ6FR/+vA
JpX4dI4crZaG8l1oBzSPAq1+6kyxoj9DgrBUp7aNc6OEq/0CbjqsjhZNUlQbK3xEPWvTid2W30bs
1qlwjtLG5EPxQpGJ6AiF4iqsRfKGa6k59s9KvFZbumfnKZG2VxGzIJ3AF24sFJ8zsnPFVqnUleK4
pne1axEc0AAGygrbU3lBS7gFfnE9726JjPPQMrGNi2BzH6egUtYsHK4jHRACVKWAJB096uvt2J3b
qzItbwOrNK9/4KP/G0dA2VZlD+PKAvlJCQ2k9VgijaDAAdkYKL4E54/WtH7lXyakqIRNRKKnuBaM
vZvXvyxyGx/dE/MUj/OSlUGdPUXHTlOFmftcPsiliQDac1PSUDZN6HYQmw+Hl7sDnYdM0SD9cdy1
c/C9NfZZgv/4amZNjEfxyL9gdNysO+lEAHDthGcBvvHJyLFNEgxuDgFQu3KMQOJMXNzJ+p85BBaB
vFUaA9MBdUl20mbjWQ2G2IQu+psdbQF1Z4kMp5oQHjBlDicVH9LGrrZ8gKqUksbSe3jX45VRWKb0
Aq/ibVNUZemh/dUqPD2XYk5LrBddzwpUTlY3MhPWLBbo2nDmHFNJbsGkYM32YxfzJiE1/W7h+O3I
UMDLHYTz+28Y/yKAY5Ny7Z50EXbbBBBPhDClAoJ46ziDDFbGyy9KIRxKmA3F9+bF8zfFbqN5oitJ
ie+kAgFjzMC+Pc9dwJDohPvHK1xxR+VJy3Aw0u80m7pp75r0M2FjuR6ipyDIrecmcgc/RFhu1nQu
Jt9Rt40DTZ1ed6IDhDOdZpU+2Xs0wC5UNwfmbgSmz3SEf8oKz7B0sd4a8gO6k76SUG8+odPT+zbS
Ssd/2/60gM7w+KzkrnvniCQNWpWHZ7rXcVoI/FAP0DN0k6MsijNiwZLb1t9xLFI4WiWe5wYuCvyY
K3+YLt/mHteIV8cXw0qfVseZz8skkpKJTMcSIy6PWd7UFaY2e4CDQhqNaOpGXz5X8vuzx5A4Mbro
T2dIDRC+bDunDh3HbdUEAEEFhhN2KQDsauJAwfpaoCm0OJt78xyIp5iI5RLSuNCZCHdXk8wUwHXO
rVC07vL5dV+m2OOFpwLNoNu/Cv6yFGpV8dlkTQoSa97pjuGRV7K1rnyjz6fGtU6fl4rUYqlXf/w0
EZOhJW0PW7aObTriY52OvvHkHIj9oTXdYyXTx/O4qy1uHQPbPJuCAsvkximLFb9dD57f7KxP+O7i
JbqsFCWcm52sGK7gymZTxt1lezcG2Ziuwm9N+MEnzzrpYQigy5vMB6PyHDsDsKBA/vgUnZlqGxJN
Y4k2K2RxAykh4aHusrkqE+dCRJ3/hI5BczehHtLeqCcI0mfEc1rVhZYgNrm+iP4cuPIfYOyGjfdf
xxEBF9uo2jwlZNR5oh51p29RZyGTK9XilypT3jW2TBAOC5WKoHbKRnAUJsMDifeMLG0bT4zqf88F
Jq95X6OH4OZFZKYkCJieRIw1jZnVH7KJvgsTeHip8gZtvUtVGtXUA1OyY/EWzSfprcz0uVRm9Id5
2SJpE/N7WfGIuahZBS/sBsVP8tdH0wkauv+uMDRpw3uHpIz7rqfeUKbkyy/scOTrSYTg0u7aM5q7
En7TP+ra6fcsVpmP82diX9ppM2UbwrzoWIgKYsHhqxahgdVmu84SbjkJha4wvdJSGKw3KIeDaE7N
bz5+etHlDyglWUxcarEUQZ5Yvb2ulBNrxHWcn9+3QC71whn1QkLL3hWji2Qd/9tjiE6Z5zT/c+MV
OPoKk7eQAeXfs4n0Vi8LKofdLH4QmJdBw0TdTP33N0h/c5ci8jdvi+PX/mhLnr8SqRUY7f1PGpRy
SUrExxIhDjnHH7ah8Pr3l/DQVJJzEoYM1MQ9CbADnuE8h12pxIBE3lRtBBSug1FjYFK2JVSFshJQ
Mt7KA2mIVUDWceFFpq3ec0s4ZfotnKNKOFfB1LIFoaeou6eA9lHb24EVq74l7AAqPB4ZibXCTjTB
phMd9E5dXgHgtXFOG4yaUZHSLOHOm2DAOXyhhuz5IlVnXkBsBA8viYfu2Q0i2bbPiMEMJnE0FMlW
I6IOdoAaExNYLIV0p00dZLrhGCawgW16gxh6KgtBpCsDYgmtC10I5XbRAtM5AM8WK+9wlayVZVca
ttYrAZfz2B5uLocPEi0yXAaYXRa5kNv5fN4CNhW8sEQ3e3Ui1dSQfgGKV6swlLMQid9cZiQdjubB
95C4BHTpZT9ystUDn9p+lN1pnNBvsg93sJlt1hDag27y7uyxKu0eONUXOtxX/HBHcL62kMSLx6Yy
eW7NBOxDK/bA4k4b79naf0yHwQSCwUZDY3fl9xHOfRbnm7oCIoZm0gfZX1taxAE872zQorbrimdR
24ofeV7vyOH7X4nQHIRyKiIbP4RDe+QemOfJ2d9+1a8a+zBYeQx8tWF+tzZ5qgdN8HvTMw95b+xl
RokeRn5EoNYkusaRMxvXTvg8/65ZAyxe2xpl6v7XKTO9LKYwMNq7NIfnOASqGDR5t/pbvJM6Hzms
fAI/TQC2pSm/ZusvcZnBytQibZOG/X7t34CaxL3Pyy1tgB5Bs+OKGdg2H/0+dP1Hkd4fP7P9urck
6yF5LRsAvTa8KnVn1TqOu/CtJ3jVMYhaQn9wyZO2lVuPn3Lni6D/JO7CUj4vYM+yFeePfRnNe0sV
vU4rozzo5E/8iNqo3FsZ7OLzENts/uEorMlgQ2QNi8jhVbMwFYaw0nk2PXIAe3ZiaTDQSfMxA9xJ
MdkGQ2LYMQdDaBAiBx8l/mGaaOK5ny60v1XkDKerP5aYdLtD5c+N/QgOtPYpH+tv5MsFOClqPYM6
KnkJWRiyRGaflcUn9zD2Y+ArdIdSmK8JiWaKi8VRB+IXZhrdK2L1jRK9ycT8XJaitpWqWI7MefIQ
eGy1ATm4SnUVDhDNUMthmla4VUhA/ki0QCiDRzbw74HDJxfY1HeGBlUJDwAoUXcujUigpobKH0cM
CV00XkNI1rYq1WU3mZG/j7jpAuQhTYPwwnJ8V4DOIte5jv86OoMgiYvXf2vgh7ekwqQyKM6GddN0
+HbntGkAFpsiKjlnrMAAc8iH5RJwyomiWfK4PeJtqwvoozy00i4WVHZxYqgUKLkM+vZGCQ+aQEUb
4woQEbJOV+3S7jHiyY3Vf4qi5tZjmlT3iRZNhLPwUUIj+1+AQBzhYiUyk6aicCXG38hEyjUCGEgv
4/7v//2VOJZ3L8ypMi0NwiiSlnnmCy2+lzffUiw+uiCV1wqLNdiNmrCtFv6rYl64TRE59ZoKo0kx
n+jOMr60XFWxnpBDrtbSv/x3hDfduUpZy42VBsoBKtrbdvQLC7dF5jVHdTEXMvt++bSs8PGsaMKF
2VMMzzBTEiNJQk7f8gbBqTSqm7IlqzbU+mTA4/eJ5K/1/kl9uCyXBKR2LzdiOXComHK57JwPlARg
BPtslLxCv7dOkLwtqGupkbXhDxJp8gNCkth+ZdSQigknEco6AdR1+flnIglVaCBxTNwHY9e7UGUe
M3+xaeOfuSmpPNOjbDFvZQqzVaP4QR6A+elWOpVa43A11hu0nWgxdJBaNcMofr+Z4KldnsmU2rbh
p5iVQvRaQOyUMtnxV9xuqT8jfZZaJcJfaJZtmP92DTSozreikkGbfB/g8kjaLyV/tbJMhVwaBkyF
REAYdHaIdSuQbpJONtgOvrHX3fXhh4wsbnPRg2guyR6ZxmbLXqIdywv0jEZ5VbrgN9YyS8W+HUan
5sDBre6B1+Cqxx/Z9kShSnYkvH8p35qZx2/JcNOHzOpNw4IidMLNaChTu8prEZRkHqlZZ6YbJQYH
YS/vOJJeZm+Q2JTXd4ngVw3wrw0sUd5EAOEBmRVckljWX/52E9cllUqRz9lrn+0+TFwGByxgCTBp
+zh95AjEbU/8ER4TkTW+GVYAUc801+xAaiV38ntH0494rWASKozgZ/drQHL1LqaXtZ/2iodNGZZt
0v8fkO5AdZc2n8tCZ9WtrJnFmAllDNTOTBcEmcz1HAai5DMJ7hmymyH7AV53rhVOpMnWsziKMKlC
9Dvz7RstT35zpUQFRgLkYbfdzYdND9IKnHboAuiKIsO4EEjhgKZVV+gzFJyQdjkI5LU2OhDR0IRe
ntvn4JQOVXpd6xJxMLcIyE5Va3upgR0xggw3SmwlMeiZ3styGDbROO3bUWy+ZkCZll03QvTqtrC7
BTZcnT73UQ+m1RxNoobp8kwgVwcnAdUnAJkIXKbVHq3gDuGubzy3dBVl3o98OwoBqY6uTXY3wIAM
5sg+pgiISCprJRiIb/gMsvHiME6xFw/4q1lr0jOEqS+lgE06LBsKxVEVvpkoRmn4D82KghZQWcNd
laT45ypUczxkXh8VxOezqROFdh2cFNbLW5yM2V8nl6W/RvvOz+HJyxZVZyomLjUXl9X76E8lXx5y
qTZrMRNK0TwabyUs6rHqzqfdAeq87bmMlcUwgiTw99dhmEQMh8gjXMx8FxuCk+cT/OjgseAK0e3K
tn/PYPWIM6iMEI5J1A9Tje4v7IZrl6CmUBa4kzrUcxD0Va1G6s109TT+249D2YyBmkSyRjNCcEfo
tsNAYe426/vIECP+ZbUvGRmiIzWyH+mUFVtOIBUb7qjKGjPgJXXT2QlKMUh5oiKJJO99iymM/hDu
pzPXZtTBIlkdwWHfe99JRUXppahxfUkgRbKpbtz9p+Pm2RBIneDND3XB8ZfsAqimDZy+4YgqPrg6
lH/0qlbUcMJ8XN12dtFZAd/5day3nALMFi+wgijp0tViFa2Wyuv4dyVYMJ53tFdScfBpBAnH5Wci
23PQ9d6l35Dx8XOwfzbLTT8OADqRMJjGgF+Q908Lf97hFkgKrY2MllYrQxnnASZwX5HSrjtbDkIc
5u3oF14kVHUDJI0tpF3mEMNQgOFQx25FYu0y98JITCKv3f/TEM0ycN/GNDnZqiHEHz5WMLfMjBB3
z6yi8KKU/CBnenShDutqLv1KL5sBiUB2aJHvBpXAZIvi4Lg4VzonQLe3/Z28yXh6RnKzJ7sf51wA
Zx6vW8YpVBWN3DyUfDjUT0E11DB7ak6XHcbDX3GilGTNjy7Ha1aKErzEWBg2rWUWL/x0l5UQcGht
/Kk06APbIj9LKv+f/4t4F6Y+TmfVRJoCRhvKCuMBz6XOlde/Q50qvoK9sx5gVVgCgq/moUsQTpC8
vuoTQQZVfv/9KRiRCtspw26x25S2hZkxAPlneJjiBDrFoVwSAkTjoospOOHbxvLA6bC8v3TdMsXU
pAc8jUHK4CgylMJ0WNdFXkPnovNdz1BA04p3A2Fu5szhjOCMcRmEqOxt3uKbhNGHaWN/mglR/7gF
Bia1vnpMog/8AaNeWo/7a7ZTjiyhUhYuYNsjYfYkwJuv61Li50C4jkik2IIXDaHRmbZDb7oICKRz
UZvJImwA/cz7MDqTGVC6lN++ezKiEslGjQNyRuM9XINE/g0b82hVMX9HZLcxKJcNKkbe/gvepHve
aLlmKoXx5C/rYv7FbIzHdktO4aZWgzU2oxEMrTdJsWWEe/M2hhUUwlHHjQ7peWYhN7YcJU4ihE8k
jlCBDW9H/AHDy2bw7Y+2rPpxRDnnPo2sTpT5A1d7ERPSb+CMOz0IiBH5IH5oePqdk+Em2SgceQDw
7gqFO0I57MbYQHS00fBHCwpVMmhPq4Jcpyg0szXr+LS+KeSvQE6prBc2cMBC5iA1BLpIoBcr1OCY
eChlAcSwzvDNC+HkVlRtb2RIWic5y8wqdqWvjIRfOZk3cZxhNDPAzF/eLwfJZmfi8le8/3hqzHou
FpKngVbElgF4XsmMY8THYSkTgApOyqB93vY+TdJtAprmWbTOJ0wYm5lt7nrbGPFbtlF5leB+ylRz
PFMRSZI1eviaLmnn7l7bazkj5njWOA1EHlBXCZQjCbw2PpiMGhJIYgHd4D+jkk2f1KYE5SX3u8UQ
JTO/by5Ac7enHj28kikK5AdWEBQKDZW/NbN5sf0XR13l59yAyanud2GZKi6mMaf1tSD1WifwMlKw
uUD7MnZEySzbT3vMXJd5oijuTn1OXum8dnjxNVpc3VCpV/7pbtA/c5IJAzmN7ygcH7ZvpwGnWlRq
sk7cRGEhRYDIBA+e5qZ6uqM15FAep3vQUw2TWexiYO8p1m9TGonM/N53BoQ9BL6wzaeZg0w7WT/I
6tBTMYPuodVi9rdEkARprDIDUR7tcLNa69w84JPnamqt5Pq7W4mWJRB3yD5MNadvQfolJRDM9PYZ
yXbb7tspAITbwFqc+pPHGtPvyopXaIgpq2uNzPKqNRR9LAb2hm0RBCtsY/Rjyr8hRT4GX4/ctGBc
qxf3blAAOzHykFr5LrsjZESmqmWYBwMqAI8P0WVPDu9IiJQmHfUIJ44XW3nHkV16q9sv5nF/it8t
Ds34hI6Iq2/JQVWEAAVa1GdM5yRUPieBnHqusP2kW9ajZNAYY8NUAsge6zCl7SWbVcOVwqzY3iIT
9rF3VfokJKyNeJbW3wBhKh958BzduuvPNf1mxHSXyX5Nxv14jTO9zXUzFHfrw8B4QPQ4UsBqMdNz
bdQ/BW8bG+q6b6reUoF3Qf/JTZx8CcGdF+3HF7kgaOHbLVLqcMYUxDRAqkH2+1jxGH97Hz9DAprc
3VKH45f2JRcHh0LabaaRyvfN9XaTINe1XEK+XTo4W6faC3Q/0RRilgxph4tUWxsHa0ushoSAhcip
/FHod1Gl/NZ+Dv82uFObM8OaSOgV/DO7KBGuVbDoAphtmWFTHhShaRP9Y5e35GkXCEF6BE53G2p+
7+VEt955eRVvlSWZpRRn3aJj8nAoBYHyEd73vu+BXpCrkGyTGi/ajauc/P8kvug4BeM4xxmuk097
e1GShgEi93zAB9qYP1k+KADUjXq8muwYCXVQC/hODzTOAvCeUGZKB0uya2cPrwe8nR6icjKC710x
mMQ4Vt1pFNsScwkcNfVb40J09QwkDN7/gX6gOxu+7piR5XLlJjCfpP+0zbv6MKfHzXUUYI1Up8mu
pN9qC/gFS0U2EMNuS+411UIBHtidqqA3PMuzcny0TsQFtk7Bi5UCbAblP4tVf/aU27lJn/LvDeaR
FZmnFNSRSmtNbBGBcAtS7gLTBcSC80fK+kOvqLxLRZlwUsITGjmN3RzGVTZe3Rruf+2xlCocqgA7
Mu5G+MBP1Z5Exiz/YVSfaGBKnkya2F9lkUvS4vTbQ18C3YF7yPRdol+grHbRqCo8qGhCw9upbOpf
hNfZgl0SXeaZ9dffRN6wyIbBbI1tIcSgCja0a9sK/EGh3FE7H6cKlba7p3fQbKOC6HHpBB3+F4+6
GmaJVgFcDYxjCGRL34rO/Gwkqlxhj1m3sIVaXpoVL3AwOXLkI5dyU57dREJI1212v2ZcIY3iyvwq
vHzFE0XJgct2uvVm06+Tx6H4yicyF6N07/hE2m9KaGKMLRjx3fvzooy792QBdsk1qaXp13eJtJd1
5ZHJ6aLTPrPrx2bLmSMEhHir93YI7umesl8GHjdxCT1qdWxvCGppOOeUj5DZ7lX+yl3i5sEir0bz
giyjJ/LUj0Eo5AVrUgEkgsGLwJ8S5N80VSC2CvZ5y6z5zsPt05MG6tYxE5jJ3Om+W1EdtSFzzuYG
dVbGy2NBbmfj6RTFWjNZS25R3ympjMk/OK51rC6iVx6aFj/Ow5sAg48MSh1fwcQaNkktPBr4ODD5
iuW78nux7NUX6hnE19FgHvgwh//aoet4jut7rFTTO8TmMj/C+dZ7Cv9nugwg7uaAmkYMz0sp5UJK
Vj8hiyHqH6GOASLvEvlFOUxTv0VaZeZs54aBnKER6h5NuPFJcEFvCM6vlRT+BDfbjiiT1tATrcK/
558vNR7LzHz5MDuNP8PVQ1AKRN7ib3mm3g4P0EU1OxNh3LblK5BU0sEVar2syTyEpRukqUBKyEeI
dY9EKmguKAi87BUf+m+BUCiNHOplBhqU0PrkoqHpgO/Yt3NEwFimnzGKnAUZS2wOEiWioxX4VOpi
YtueiycFRXbxvI9mrSo3dbocrLsN7z1ue3JCtfMvlwp5x5IaQ58zA1gvljBJNRLcxQpc0qMwK83m
uyIjoNCLFVX6YAGVkXi0mL8CIeKtTyzbcOSViV7oqiYGS0xQ2dzSi9r8NdDDY5mxVY9j8TIC3JqR
lce6r0N4vRMMSGvhgdGytg5x2MdUZWzjILkEhbYD7hsgKKe9p2mc3BJMi9rM3UfyKTl0vPs5s5nN
JyM90+H2vozl3PM2/FH4BNN9Z5eOyo0e8OTH7+lySFwZvcYDcZ1075X/NI7qTGhO0s4Msy85z0CI
h/AsbkMsrnhvBDZyxn0p2M8vw3R2esqfSuO2pBrwZhfg15eB9LE3Un83yA18j+B2DncPqoN8+Q39
a7jKp4YC/foOizw8X4STK4tUVTddW3v+W8QRYlUfCbh1dL4Us2o3lXAAYdCRzJCs4KLpjLkHfvhM
kwxahW9Tm2RNmoQ44LwNXlZUD+16Y+oGEwCdwC3vvuDWnCA7/tMFPyVYj4uXqs1slbGNcfcteSZE
UHwD2yIZbXEUtJOmH9pST+lsrbTfwMmn/OfZ7sINmTUrG2Sm5aRxSF1Re2VHlX1Uw/3pefubXcA4
JO4mm7DugBdducQWWRp3kTuKqytzwLlhdhpDMd6UDpidoRXun5RkQLLeG0nX/VgUOasn44Wyr4++
sMGeg0NiDCU24NN+wwL/uKkE5nw8HmiNHk7CDvfL6Jvr0LtMYJ7wRkI+vwThpx9erjCVUO2+1h/r
KkN8NQ3BmKzYMFuMEkVtDSnbtON749XDdRA1HLWTTmKPXf1Va1waAt1Ax8nMmtczweVotGyno0/a
EVJCIyDy+IuolxH4qzBT42bAwQGh50mCE4dyDegJUZAwPfrabT04K40y3Ql2ukzoOomg4FOKFmfI
UOQ4ULM0jTlD0rSfLcbD29LC3seCutYpKYlqszQegXxGJSsxjt+khpEpkHhECTAqgWkvrNzLNFzz
KbJSZWRr3/2SHww7d4DQi4JHBeNOk1wuisZZWAbtYoSpQlpUn6PuvED9Yprm7b6fQ/pLa79Dupg1
Zpc2l3V+Ql0hKdGk0RYNUUZQegR9sdwyBfZ9i0U2bz0QZBx4r3TJeAQBNBnFOUcu7h1P/aPGDWB8
FXPaRi8W1iNyeEsmD/9+mnwXOitdJJ8jE+VocHRCU+eoXvwydkLZ3rX/CMF05H/JPjwykFgiXtcC
tqFQXxWVvTptxJFD/5rl22JbLB8Q9pE5Pcx+wa+20+Yz/7S9kS7q3yrZ02Flpku47I7NZtwwbvH/
3HimjWLxWxy9M9FGEQhIC4sye3qPEeuLEXkXJgzHLegGIkyI6t9DcXegFkFFYqUjuvjcrBJJ35MH
MD7smQAxXW+Sj9NfgVWeSe4A5rWcUVhf6QS53mBGxBgwIW3D0n+leV/IeZKmc8JVg4fu4bq14hQ/
Ux02libuE9HQHTixt9b5gjqFDuLqRTtE2Hb2CjFWkFplgVqxGhTNjr9XOLQ6YlA3euFReceFroZE
ZKy9c25BT9vBIMm0y1KCXzcJ3NaUXAnAAkWIlX+UJA5IzWRE5xDfi/3mPUrXgGgbBtZtwZXLoJa2
1L1shHe66aGqlQkgsv+i1Zq16zolYe+S4UThMjYtCs36mUJ+LwWakKOPxQr2uIipbqum0EGE8C/O
isDJn6Pk2oNyM5L2WEOAFSi46mia1dKYd1y9H7dToimj7d/g5SoH4cjVuzBU3SWrYSLt1mYISG2c
F9d282b+LamG5iPpjZ5LuTfVblwNH/FuNCTthCrxOEH77u7jFhEUkREXkoXC8gLHWaRlKgL27jBl
xXHZxUvbEsoKCmZGuGYSdBiWgjDNrLGNMSesvFFh6niGuafGarCufgyeItNgjeTGF46szmfDJUz3
glEMClyWmR4VvugwV5sW8cgfjS9P/PLf387O6ONam6MX53xPu2N4x6J2umGFlff49RUaFWNOH+5Q
zmV3WdRVfpICteGCUtE5kJFnTl8SnrOPYV1YKvpTMMKEHumHiDJjyRoWZGQco9iEIYayKzpK2hlZ
nAD0PBNL2XU3BdzuFJu9MOURtAiUXKmwd5szJVaVFPPGECCCMDmKsm7SltlkCKAoV+wiN7tY0QSn
nd1CChsDlYTDLzXuuV/90rmNweCG7V1+E9lwA2042rxTdHMvFMjQ9lBGnAFxDgMNBhe0raRGBhHb
G/PiCYUFvLOr7NFhJiu7fMZsDChovoc4iMiJ0KJZFVtF3VDG4HgRXFHNMMUNhZRHNaFf3Lt/I8Bc
90j9rAy1CZmuSYJkbByUcgz0cpHWmyVJDkHB9T3ZCxx6k5UQ12vLh/Im3RR2Qczln9obLMUvicse
9s6EoSJbCu4x9Q3mAelCjY7228FcDguA/Gt4xCu9VDrvE7Ti12O1a5+GYJyI4dMcMuJl/IJq8kbB
kXDjPpGjsHaF/3oNoieCW7R/14xkyAI93BM67u8q3ctAV6vgDMRGJ9dJXF7NuM08Rvl69Wq9XRbe
R+3RO10wX9ei/8Rhl/KBkTB4yxUXM9VejWxcoZC6PGF4PRXUUTuEZQ6o4IhYCT9nHhSPN2aZ16cW
VFHzRQO9pdOyKEIKSuJHk1jxj1GGPotuToMBev1bro1TWvbwjUvPy2y5pSWFs+qYYC9tPHQkgek5
MWBnJ9RX+W6YCoGCyXuWsJTYymmXAfDf/Rf/nW0vXd3+phqIjR6NNG6Jo5JIAcyHjlVluNN7CNl4
ymwfkXjppbZpfo2eE9GVoVjKaNZt+wtmrHGKJCoGXmVXONkRcaMEUcqt8p0yg3nv05OsWgxAn4em
BT8nmBlgtX1LgeeC7agXlT8CEdNzCfKcBGrfkwLnGnTx+JZ+dqiiajUJ6JVauIdcsqpod4XS6FWF
FHiC4O4tWjAMLMBw/Swg/tXwN6a7AAm9KmEUCNBmnfr+4MiUaI7v3fbfgyWobZpTbnfXjJqvr8Wc
sKGVTU76SyQTh/fLhe8S9nuchFlI/0Czxb0UymEJXPFkDMjq1/hgGZaONYPpIe1rlrCfrHryt2nU
47yV9Hk6lQ/corzTrPcB9N707D778OH43ADKPUNztkBW9DtPwH61MeMkCGZlrXdVK1tpH0OnOSAA
MiUY2iOKx6xCnWe3MsQRRlP93xPmVLuoqOWAUsmGtjxLDbH2cqOy73eAysayTWBaZCS/KCo0nh3m
kHXmtlitvZ0uZAuhhKdwA399Z6j//bD5rnLuZmD1zSeuHjkJk8RfVauLVaWJWMPUS0h/VgTflXKh
uKJ2wY2e3YuPLE7bnrTc/8yRsb33Dt5QZVjRdyeBddpT2zvJb4B8/85UPqrbZC327vUBkpD+JwKe
aHn1Vr93JTTb3I0/fydeQRHqxhPB/FsXaARx/HoqnvpOeGDL8BOasGDGXltMkbMWz6o2r71evCQ7
TH9adVwU1aGRp6ThXpEyhp0BDKnc6QGSlYAe9XKkk2rpZLcfoOOHZzKo496Dt0g8C452ELF0CdP1
GYSiCFEpyiZs1jcB1LHmUuy9fuana0neBEf7ldYPk8lUWYbF2utAIFq8BpurvLXmVmeYH36Wc//N
aJtVC8E0N7m2RebIOe6/xK2ztrfg8J9dQ1+DB5MdTZNnRrujTu9SaTDwTLbaKQMfP+DNsZ+4vaZk
6ZFTMeg7/ef9SXZcBpsX1WZ0Z/KpMzR0WSQ6qkyeUiTrwBxjrPz9T46WyORPGvxaFz783G0yv9it
S+8WhMceyduIkl0e+/BJy/ddP8xrqqVxyiljeHBWo10Cea21dazOildtx/Ao2x5Bg1wbChALCmH0
ELuOKOPhHCqjrnhbtdSPrLE722YgjC3tuJYz1rF1dqAhY8GQWu7YB6qnNx/t7YUsdCYSXVeManEi
0qlSZ+xPGHO118VBm/qItranq0DIgLn0wm/OPLOM0q7R1urnN8Pi/S7O9JuVQbbqjZSwBRGNUuTz
nhbKVFQcYnIc3/lH2lYgeYRiXELjI9wCIyZweyPYrvAuETiN8+TVWGwGDnhJBYYZo++aiaHdm1yt
21RZqk5XISu3/aTtmx+dtnocRLe3ZyxnsnVccr0DVz5YFlEm/DkBQlLaiKQ3f4NL/VRqVevaMa2t
EH0Md1Q4byaOO5LakY9XmHvVbhvNwZSCeGcFRI5Qusdw72UOJpkP9kbIk0NlFL9uipbzi0T/FItl
08GokGcLkdGXg1nwu1mlS4NEVTbZsKDuHCLoS+P3DWPGDI2VlwSBgWuDd/RmTObR9g2PYg5iGd5C
Vc9/JkjnFuKzhsdavTY6DezgjLgtYxEOeIMF8K1K8ByVgw9RrUZWxNR8/hAHdYBKGnh7rW2ADmuI
wpPuEgjffZGqwNakvj+TBb2g+lzq+p7U2Wyy0LzmSTJDMkuyNLUob1P3SZEIXXwGi2xJHSu6LD23
bZ7R0gfkQalgFnnHXRKW9QqGMxiBWJ70UP9WXcmWNW70qqnAopBcdp0JOTCU36smVDrEWoxWrvsC
4GBplPc5ZIZ4ySsfF2lVVjod/sxHZpnbG0AdbGBlGPSF+SKY6+LHI2NU78ZQ//CgdQR5Cd6szHTR
QjRDWUxJQ7SyvSKTkRb5j6SruJWeFz6qBha0J69Posbywm1b/cN5sKSEGvSOxf1g4UuHWlz0Dl0U
Kcw7IKvBlEPm9ZmjUH0/QG87qiPqEvjr1UPxwDf854bjX6T3de6x+ZChhSJEdv0DitCQY8MGHIL2
ENzarsfG+e019/2BAV39wWgyr1qsQvqncTu7Ea+nIzxvlAgd2LFDlNA+O82zP5CuSTagvb2dha3B
bdebjpK3AIWQS7CYInPDNQKZC845wliY3RHKS/brYXZGCrY6FIZ8yyDKMbDQH/khD5u1gz2FGCws
h8pcX5WvTfz2rPYLBxz5rcZnh8JJUTq2R4wP2sYX3XOmtqEfDky/AkgXXuzdKSH6DL1kA2/U5A40
O7Mw9U2eDketmvkvUnivztCGVOJ4eyCyNKs4a5BXW0qb+Zqy2RC0kN83PhxjTKg1ixtxkPhfpoSf
yUZ/Ruhrk9L2lPtkreo2Q+tuf+uGL6l+/4ne9rAVKgF8X7UASrJrHdHsYxUzH/zRIo60mVTxf0jl
G76WvNtEtxDINFbQ+gd2s7L75JNT2ywIB76VzD5OQUUgrPQZJM7ViAzg1EAzfePsME1v9/EtVYyD
yfsxsX+K3oUagj95QBnG8lARXNPYPvHF3bXGxc4kk9Q712ba8cpzGYSGaLdmtns3vOuSkyZpEXHO
sxAIJoStkymdAafZ73II72lKGfvHGvdAYwlcVMWhivuQAKXWZPxpf+IwHKDTFK0MJ8rxJjn16qFj
RU5V+DNOZb/TP0JrQsvjDlalxioBzcfKhRVd7ctyaJyrz/+RK1A63dQ6bgUI66WCyc33WcxENqo6
p10p7vOxQsxA/iCipT4x3L6zsJMYawNVDr3Ln4hFVQKmhIgz9C3Szo/eVULa/h7LhtoPMIWMPKW4
gGmYAC3yVeJKfYKtafO5XqLgem6qYSZF9hLasSDTh7zWBAUV/EIwdCwU5IILtROI+atWry1GhTDa
DMwEInL323MQzsYghnWCaqcgTM06srHReBI5beJtKVw4/8RqVZkl4sejTFAJ60gAGRaiDKJqjsQo
V9mDpotXb8PkWzg6POp3xp+XsARYTQUELG0hZqQ6T3/PMaAyvxJ6BPiOoJbrK0+SwY8KIV7fNAYl
l7UvMytWZ/DXALcXjnDDinu1h/iTIbiVbG5dUe8wrKDi14ZfMqFjAxxk/iDoTRTy0o2L6IzdZWgb
S4ILfltHxzn8vRzFnNiPWcdyXjn/f7EZNhbp7FRWPaRcmLq5WHVF+ND+AS+njs8Nn0+Us7dw/c5o
DcvKlBQcmMSzdgQ7pTFSfvmfTYSbDVnwut78i0/ascvIe2ysIxECxjlrBJnlAOhbuzPXb7nXG0ft
xscwWeDjTgkkXHbp9mcAsV8xBp4zKq5I5ZjZQyVRvE+9h2MVroFyAhIW/T/IW5yoQNQ4UiBK5374
2RKWhB0o3+pxs/psuFsFR9FgyUAI2pEgF1EfRdyvIduca4UyXwkFtgMAPc0DTr7jRCc2jYOMvee8
JaP2Y1wk8OiwPwsBIF9WO99bUX7hRcBmAd2IWo20V9dMpL/Cm/SCTEEsLLYRVoz9VRstCt0fxxPV
+vm6V4PmiSGlyYyb0ju07XXeJN/quQ2kdVWlMfJJPRRmYNT8Luy5EoLdhHXHKP14pjpyOUSi+q4z
UILtCn3aVczCfLSdQnYbN77pGpWvsSX2jfNRBj5g7uKjrdf2I5CSQSWwIDW7M64MYFoyE2uafEbn
u5zMv1cP9F35Ii3i96HXiSvCfGC9QckPzQbTfOWSCLNgdBMo4ZChRygLAguL6KLv350VtVxoYa9L
mj/rXg9eH0w0ynAX3dfSNV0mJiAS1LlCZu+rlakeI0QBUBOToLPXG+op92eA1bJ1QP1qD+Qt5ljs
7aFkABPde0d2JkZL+Cj2ucPD8WGufjdY7aaCQPQmO3zgxDRMEULqTsP9lffdKRC5fmSB4P8I5v0a
vQMJbCiujwaYyfjxpyzJ7eLCMC1duc2Htdfn4HREYEtGyAf7oAv++FFREeonwekJy+I04jwRkWaz
YC/l3rmVfpQ22ySh+ZA4YjDntgKH7x1F9rH8rvjOqg5wyyA6CvftBFzABDk0HFmEiZG+sTayp6cU
C64EowI6d/eTRN1N+wfqLU7RmiP6CtFtkjf9gZiGG95g2FcikFwxpKIU98hLM974BBvIVxRbUTQm
KWsHm/4/V+fSgim+jL5xJnWSd9dMVfy04hk00NVIpnb9NYwBO63YJ5v9iCAzrNXpCZKQk9afBayP
QgQJBtoFIfMQia3gxW62OwazZf2yRumox4A+R1PYAjvPki2YvRaP76KaE14oiPZUPBES599FM1rg
rsTuGBHiqqy0avF9MUfhwwbEyYp22rZ6rX5wdZ2A39SXaVI4jt7jRVoekldn2GhAob0k8Jg//xGP
nrbQCsXCGKoTTQUA6UCuTgENc4phiZDwA9jWgMPC/53Mok9NBYeayv5HozURABmP8WYi1F9I+3Ek
aj1+QFxTkx+yaRdyJokYHutND6EGmOx5b4IfA8nztvz2aN3+r11JlSXALqcFsr2LfDQfTnqBmSnV
MnpwBLPMvWEJhNIY0iwL2nqnfo3//sdLrkSeSSBTF+6AtvhpYbeGUfsLDcytdym7g5jU5tu0ydNS
dpcHeXs1z2+9bcijgD7XQQe1fwWd6fpJ8GSfkkcfaBkQnIs4/Pp46X/ChwCplg2W+xEQA5D0EKl1
rMg/euGOhLtYSG/uORlwJ6HaU5oMiBrbBfPZG/6T6xO8wKiscx1h03KCOn8YJAFQ7eARjdtzUv67
ZltR3K+DO729UxQJoJvsi6/qxyxCAzCH2pBOpejiJT+QS1V0S3gu9Df6iNpJwzzCvCdSiZltY4VH
kO6VxE1+O3BabfQInIzGfSicZE3a9e2teTAg1zPyAN3SHXnL9ZWb/4O1Yy8CK4ijPyRg8DL5xB0z
RMMDd2uEiaROB0xiEekMgT4dT8JHtqvC+PfpYTGktp/Hs1mHeO4PJ3ZyQpc97TkyvFJP9nHN1ur1
m3ykAFMA0KK49gHVPNZez9ltH2UtbW6ImpFZGgqzrPPuS/ShNBmOL7U2wnFLhDijog8iWYIZVhem
BFQVfv5UYI+WNOYmH+cZKuQna0XwZF4zd2UkGp5wdKi19awKAa9C5g0d0vTFPPNQ1Xg+9OZxiNY7
Bram9apJmeop43opFxBQIi3MCaL8JVMFhio1JcB3lAExMZwzmN9o1dkD8GdXVdNog6ECgfNpZWaK
PfUhYDUjjhlpzysh4ZDj10xdwHryVsfeyQAOZgAYqMTa8ba4s6B+1zRu5YGhvkD7Y6bvTjAFDRKH
UBEU5G/9cFPE/9j2t2sVorbVzK+lgjtat2qdW3fSnEZTndbA+MQs6nMlX3wgMNJFyhBTU2W7QVKZ
+1aQU46UryYE1j+yyJKYFTv3gUwKYFmkGzqXqyhXj4Ttg8LXBXQy+rmpeSnr2nb6BvMbJFASYu4F
szpT2awp2BqCVoKlxYGmOCw6JImWD1/cLMXfBVfuPUFE3bRcUe5j15yYe8DDnY5RZ5VqbvcYplbK
yZrMfsTcJoY1mW84qXCmiVy6oo4JDi5MylKyv3lUQvNA62VnUM2PONZ3D+zrZZqp29zN05vg+3vd
A49mXtzDDXY+JbIpff8NVt8Dvwpme389GNzx0k2tO7fa9+KkNDrvwAgun0ejtK63us/DBS5dDIKh
1cT0WvuBdHP8m8eOgMra/6exKsv2cChYyb7vhYuXbfuItNfIU/oG3lzVHxm+7dcsOQSC5WsSqjyM
jhooa5Y1K0dbQlGosJthbRHwxIREsg5nllPcxL0CbX9r2TLMQerrCctQ+Fm5oArXww79/XTp95L+
3oZjATn2IYEF0P1PyHIf+bB6uHa8Y/pRAyzzIraTbp/pCtbnDI5vZSb4ho5qo+eTnhz9JhYrzmmu
7ySaAXuuLXyVySTTRR3u1MrogkOBQh0Yvz/IrsjxQfYbbcYNftchXIPS4nh9c1PA2ft4aP8aSCAe
iZvkPqo4eBvvcpQ7fGwES31eYR1cfWu/JE65nQLRG7uBolEryAkJQ22SUl1Pnq0M597UTdPVNILY
WR9jU8qmL9E8oaD6eTM9xYuFy+9wTnXWUBfanVlodlESc4eqTQPwUgilYD30XJCfjuWTru5TQuX0
jOlX3tNjAz6XKHghW9e9RaagdQyammOB2MtLgEmoS8W1DKVGLH9XVOycpBKpd6hhfHqbxRubnnqc
WkpmPjCI9RXFEKmNp0K8Z44Qg+UMAgSfsUhoixJG4LlDlFNBAn+t52C4+LAi9Yannz+S70npeBku
BaXNAI6ylrkE8pNA2n7hlkoCb0trojyfQGBaTHvdU5XxPquzx81L8rOL9UR2Hci/yCqatELh8BNS
G7BF78jZb85ZNl9Vtd/kwosDl/pZNDXFOZ2ANRC7WIoG9/7z92aIVt7oDTk16feIteB/cQ5feq5v
PUZZKdIEgPOp7xQ9kQ1wPUDH+wZRRVxblffK3PVNOZT04VcuoPnkpYfawL7TSjpK8YD9Mq64AFSR
lTP/I47Qxx8mm1dVYhMZCcmhpapsQ8GKUl4qJBYBiKV3mai5wXxqtd3JY6EBpC8aNKt8nbXltxzh
X5UJWeuhf8EdbsfoDPIb9Ex+LZ22peThGKTCALkVQdQSC0FrKbTTEOY8Fpboq0dpjOuxhF7nCYpM
pzFdOhsjuBWK2s+YQvBkz2cYG0i3miNUwtqzWEy8ARgpWFpYbpacnYHTkgAByDKOibqo4M6wSJRs
7sNFsdLmHVDFxK8d+O3eX2Apnc7+ift8Gy+YXCZjkQiza+ck1cONFJrPu8wq2nn8mGJaEJPeLXjK
CCDGOsVgIa13Inz0rzujFORJZp2sJ/lzmFj8EoUHp7k3yZIteIgAf1mBYjfQlxG++dvc8EDGqCh5
nQT+V92w1D6+1ZoRqNy/Q2A35jhx+0MNvyVLRy/sH96N06GsCSbxfmmOHmeQoaQHfjhjqmhqDzgg
cLKLtvpnMffxkFdYvpvqoGQDpykPa9CYrfBrQ9rVQVUk6scbCgcP83CL3fdNIkmud1mv4lWsPRSm
q4Y+E7y+pXnrDODp+B4e+Ou4Vy/0pt8WnpYtggJp9OX70ZcpOSko2rCrrIkv8zH0Anm8jZC3g3zQ
DrhDemvOXx923o3ZmQlfzGYH4vRlHvI1kR5RyUQTybkP6ec2BiE6iWRscDmQQqvlAcTIZxQ/f4QU
bqp8peTX/3+yYK6YJaT2lYDDnmToTLjSg9/gh7E2HRPa3msM8MH58/5m/gjST7Tl4Q90/aK5WO6W
cZyXnCbVr2xP5J0dwoT35r15PwcHZRNkJYwo84Rit5oWbwIPVDIo8lMuQaWIS8YeKfmI7dtDTtmg
GpEc9PJUQm3FJoaEjSZYSVqSRWsOMzbnl94QztDU7yiPBKex4PMDQP5ZYUSeZEnhIjXLe8P8mHzw
yqbqc9hhB0/a+4Jou1QnmQ/PDtO/md3p+P+BS6mLD4U6XqHV7UBFtz1MClT20/kywKPyZExt7xft
fkm89CACl97cUEl0HJTqkFmXu7aSFybti1Khr3trPiSMkuPblxlBWvtLtXl3GpLE0/mSZaBqcatz
IiKH3RIhrn8Y/SjbUsAY7MBkYZai+Lbrffz0VK4i7n7LIPOIEhOfAPrZj95Rlfi/uN1St+8ktMgb
Xxd/qjntB9C0e1dIHCQEafeCI4rdpbPci3b3lnFPqh1yqBx31nasiC4WuhD+UssqE7ia3EzWWgcc
wyLIwSONGBPuu081WzsoUefMA+Ki/SjqOgEo7n1DAxaAFSH1MWGzANGCdwMnLzy70X8DYcfn/tsW
Ylh5kBFeghZDM4hNH8MBlPiBpfvHz/TWLW8KkM3FN0Jl4sRW+VPZla4r5A5fxe87XxKo4bOQmSwp
XQyPjZdM00LrwOYB9tURT2BxlPf5ZYvo2miTibQXR6VdhR+K5Eo1Ri7OuXO9ksQRsUUQoYcoDUZZ
ir4vFNQzEU3CTqHj8IGb/eTASYYeZnTzgyrXuYxPilk7isTNpq7TeLylkDnooCJC3JrsYREnCsw7
Xox044WRQ+mQak9vZVJj4f8lOWBux/wLLd15jKu8yndOc7AfPCBSleL+FsHjf419cHEkxTC0377d
U5U1qqLacW4wHJHY3ujUJKUGY/maNneNSod01OLuokOf9LW4+5ogJb12jz29+il3JvcISFxl2gW/
0sXg0NWRPaWODV7Mwb0c2Lep9kwI2yzdjxGuL+Aaqs9Ec18yunsN5ikPZsbroXxNUHQQykPscK7/
kF8z2uUvIpu6p7V+j04maANIgEEHRLfeS8yJunuCBbiZiVL8S6xQxP/DnpYwOs+qLVoqKmdf1Thb
LdZV7q8IcLpFc8a46TXzpCsk4GqHX29HQTqetueHcw5mEgIz70yoL4wQCivPNPpvVn/EYCGOu+RR
J86Vnqd0e74gRMDqpgWIo+ylegmoEktgbfA+wPCgUoVDVdyKB2pca88BaiCM4CLSRi6HAAFj1MSO
e/IE4B09teyfwmGMsushwPyT0gK9t6tJj0aqPCnSGX7X8RR04PV8eLuPTUXxftoALqPdHaWfpEDP
tcFJP5QxgsixPts7IS/LJjNyHOGW6Jku6260KPWcg9PgZLmD808HDsR8ZeO7BRLJnbwmJE9h79ho
zsTrHNggLoYNksC2Owbi6b80eKZpjl9/JOSjz/NZorCYniB5OAp5hC1pugQzdP+wO8srYmiLShVw
WT84UoplOaTnrzKHPB0GCryRqj1eRiOLxvIxePslbm9xSItuOLlN3TIjuGx6AKYSOUr1EutEgUBX
5pMeK2y4N7VfewwQL6RQYkez5Lvv4PcCegPf+piL5hQBs7yv4KE8tgFu+HGzh+DhbMFpouVKKCoI
3NZcH6x0qY9YkLpbubK8NrSGTk8o0gEkNxXWVdyiruupAzWZtDSXO9sKRg8tvj4HRkUZp9k1/OjA
PBpJwhke2nVgq47e2ulkBFSYxUD1og9gnitOFmGoC6L8j7zpwxE06BqRVAa9Qcu5doYOB8afp0Ai
cVmf9JD0JZcqNRNWZr+ZwC/bj0+xokrRZElN1DHXaM3NigUbSGTb3wQEX9euYSFWDuFI8XJVjFGa
IyBNoyS71W4DUtOgWqnd/ZL3FgWlEs1oJ/AO9Fzd+UNxM3iMtHV7IrP473JuPCLD/0uOWCBcOqko
q8TlrriymGmnhp0RTsWTOVXGMB8KtZYlyXh0y85WoI9ZLOr1pRQseqgFrUWoEr3sTXobeLcoLcQc
LQXZP31DDpVmHyet+sJZ+Z88bq6yfxvyEkFibym/dYwVbXVgj+EoCv9FCVvnoj8Qi/YNuKNqAWh3
R7KKuWU6RJkno5yf0DG/eYAdoCebvtcYsV0LZIFtV+t1UlHs2yWkrxNOUzzMXJgoAUavJhAjxbMu
sbodoUBAsV9O72evqcKaeO3LGG8dVLBwgITsOV3QW9XtIjjDyUjV4UNgnrK+fJdSD04NmQgH5rm6
vdChPLbgy5JZIKBqBd9I0sA5T6GSX0YzjumVQw3aUufMo3jAi2SUh79wKpxbms20QQRNAmzBV7qq
CCKl+TXRFGTgUiBoXcQL0UcAcqAAlV/ALptmzhXTQBO+SzD3rihG9KPPoribdtqyA38zKlruxF0L
tv1N7KzACM0umojo7zzMvkPEN57j9a/1yIaQlg4oj5awkXHmMP7bRdMNp46IPsEu/paE405QvE3J
hd5qgfugR4p3xHVIB/Zy1jF4mr7ZRYWTUjLogPVZnHS6KyjVMMSLheUpVwmn13+PbR8ueDdlL4mN
RbqCdpuylCbqaScLUgbUTCnC7Mnxyna6EXMCR4VGwP8ecVP8MZQ//DR/14OXtCLZc8uAu6YHoEtY
k5SDmisdPe1CjXInr+c7meq1pfUOL/JCo/MF+H19mm/Nq7Yys5bdzjvb8Bt0Rkqnirgo8w8vXZq3
DwNf7gzUs/bdJnxdPBOjsQp1+SmX/BI2d1/E9PAgY5UlNXFWVBS241R0rvrMhXhDC35pMZ7UL9Od
KpNeCy8zdGttU48Vg6UB+/mrEvdBcUhVqfSq7+il8yb/5kcCiTDWmYWWSCNsDrUOZnzARUNLlvYd
SrkJ89J2aEWWdIHzdrSRePKGdDq8WGEH2oK0EG5uFzp+X7J7ffB8Mw9Oty5M73Keog8W2sSypGL3
blhQil0vZBQX4kwq1jmc++pK0wpoJ1ZasshRUzvFZdgEiIt+ghQkyDMixWcMcs+ZH55PGS+vSKx6
yaI+Pw5ZdbcryoG6INeQfOP9u3odGHYD3u/wgNBMR31arcoGpV+PXizNw0k20WYOVP7mNDSyBG5K
fHxZvcCf5abdy7huvVrHwW+y8JNL6CVzImuxXGBb1Z0dKFcNYRMZ76CIfJ7iRhZ7EmKO23HVwMz0
aDRjVnhnbaGZJPogkQx3cRlFuRAXCQwkX1nl5CrZ3JL8WQKiaiFYYe4Lg8Z1zmvjE+/ojTpEacmC
MbfWzDpJGpwTHgVMIvi6YMRm/eJ5cGZy8qesj/hCGP28M/uSklcXUrR1xI3dD6YA+dccku3U0mf7
3OdI4imo7nAPS4nvXVcZuy5ee3zJqs18fW22Xcjqa00+03dFO9hBdmBWTsGEaLJXdQIfcYDg0Bc6
aOVPvWVZYdqbr6xdfWo+McaugIMaEK10UVO8M9Ifd3jSCsw3O/RY2scvQWV1nLlMuFTxK+EKd+VI
h3D3z9kcjO4NV73fce3s6j8z5FY7RoZYujsqV84VwTyg1N19cfMevCZtajL9GjjHL36nJ2SJSDSK
7z9qeVrIQOA5Ofidln90r96A6MWpqbtRVMG7AmGE1cgr7L18MYGzzSkIEpKt6MtwyEk2lskYJ/RX
I3/p3S6ZAWi/yN0AdOoFOxYqZ97dQ8H7vsaegrusAVVtgSXY4JzwvLABWandhjp1+ViuDvxI70Js
FfgnmVp3lq9Y3s1WOcLFGaj8pzusvU+INgFyDBSNTF/rkN6vN679bnv7SXVAckB7j+Exi9WuloFz
4Yz1pFqbmiwbEVmZ+1xxGGMW3pZtosxKY9zsRLzGAjf07fyRlwWXO627gnkshAiAi+N/9yWYEPRV
SgWofB9xAigQOebJ8ctwZJROFdlbZZy7zShV+gUAyL4BMoixrYHI/i4bPzKeHcaWTNjsTfvK2H6M
AT14VJ8iRvOhDfCK5EQFBoOpxmqXXIz+h8ZXHqvOS/KC/1F08p9wBHscbUE4LjXpcsIrRkixJSQj
D5+MyTFEfIkbJhx53Lum1NPnPz8RmvZIZVXAYb0EqwJzPhr/soUtx1TGCELD7YoBY74vb6hv5Vy9
KIuI1Trfg4MQewQcemlYRgMCcBBTbFIE/Q+KbeDYA1lfwmptbfscjiQYkDPynfxDU+Nng9dLOqwR
Hzbc8DZmlNRlYz7fH8gJuIzQpPJynqjnIJm69m0RTzRW0YxQ2V0FuZHdU1aONas7ydVLq8vDi/ql
DEUBJ3pfpWbE9iNOoBMLEYTgkI8P1R/rrgoRprTGIznuzvd7ZLx6KGu3wcrs5NS/lkq+pzrG4dB/
JDUkCfDaxmkEzYHE6+UINo0g5nDcygp+FpBKDKhNgTZcexHbWEe4ad60DCmqZf0J6utg8/4mL/k/
RR/M6jiCl8JmX9YF0D1c8CPrJFlnnMOizbYoSyfhVobP2lzMxgkti9KWi3W8dF0oLjbMVOCK6mCC
+O9olgIJN15LJZ09m6VuEDXFlNoFEmnVwk/l58ziUO3RCieG5qSycXoZzG+ySACcdVlE/P/UD5N0
xKmsNj9QSTdzO630asbQHJRtOV/02hB7AkdrX1MTpsYJV+0GG0Sjc043Q332KVvFwZX8r6XptSvO
3YQG4I5D5N5CF0DBKcNHAITzDjialcgLTFnShG6aOGAd9EefH+/hdJc4wD8F7t31Dy0cqMytnPP0
MC7jy4hw5IlynfWd69CBODHjrg51l+xrabn51UqsC9kEl3RswLmI2te+NQjo50C3RZ4UtM5Tl146
HaLDCHypXUKdp5C5809GfB/qYSBhZkfBl9MXOz9kXVpJyHHgkQjkQL37XyAvrFKxZudeMOebEyDh
tB4b1lUYXmTEdpj1PazyIjIZ0uFSZ4IXSpG8Fpp5ubH3hW8/ZHA57jA4CLlmRAwgkM8JAdBDCvHr
HeEV634k9QCuZUg35nRMX9mkA5MeANKjIvyohC05ohHfD8IEAIJN0hoMAOY6OWO/wCOubxACMecW
btGfvx5xMbIghdlVPCDrfJh1C7/XM7pM9ssG/8DZvlnw8MIUa5NBRvJlPyn9bdSecJw8ZcHWPsxB
bekL/ePPjhl3YqOoSK3x/mhqEWKU4SIIGRYgUyAgtaLDqhOIF8vQut5UC2ji3pdNNTsQRulc5n0L
fCVr6F5ysem9UoQdSyQXoiHFokmrlVXwFa1YmKBXtisJj5BRAY7DqKwJkq/XuxBfyptW6ym7Ketf
emovllL8EmcayjNVGl0V1+0tyQ+02wMjUzYh9j0LNjuRV46V+pGYy3LAb/QMl0eiRx8l1W8otD+D
BkpoFq/eW2q2UwUL6/I+MyyNV2e5lE/Tfu9jY2wdDHgZJH+4uGH0KKCZEUyZZRctkP/rTz7dtroi
+obGGZ9QDSTfeoLK72d2EqaHDHYVJ2yfC50cW5YoWL04go3hkHba0Bvc+24czd3G6+40cH4HxjPD
JPx1jScGEBwmYsn507wwyTkjNFPLT1acIyV4byzxzzPz2ms0io+CPEX0Uczgc7URw6Pfz1mZXXI/
S7AHruKKND0ch1ZT3DyeKXFv0yqYFeKUL+JJGia+xLJilUE5M3W53fdiI9gFG43GUiZtasw9xS0u
JLQcWh9eOpHv1mGnraPQpnYuRJKNFZDDH+/MfIUgeBPkmRmIkblle4B5xLTohiOFIFd+vq7/+RX8
M+5mDloR+RWMOQTTWg6iXoDMzMw/g9PUjfKLsTLnoNBO30tchQV0sixKlTdc0RZcS9BJ/eb/JrCH
uatpx9q5JZ6ZqsYCUyn5IwuT0V3ySTjBEsB/REWf3cjkahBmLRJD50Is5uggYYvxASIIN2tmIOD3
Ra5TVcIGguxqwuuM9RaqIBMaSGusjLGxsloF3MNemTIkSURp+NPaI4MFr41utWgMgVVyIDrgSMTy
W00rNA41SL4mvuGMMNwmoI0+OoyNhBvSPfzSPACjVIHIfTZirr4Lb1VUDqatmF9eVvKwmj4SzOqk
9cUDCuAqb9mSZ4auqZK52eR2FqBAiBtrGjS9gYvZsI+iV+qDswLN8/DGBVC5Php6214LuO4XmjRs
V6zXAPqyaNWtdfE6qsDUhkzFxIGLI3vKewYKUVyxlBeI5Q08z+Uw566WCDn3Nqj7H8a+E9XqmXN6
LRZUkHY4bIpXFFDjvJXAJvD/zv1Nzlrjt133TPfUcHaWFL31LpS2edFnAYWQ4fFC3jj2KHXJ4y64
DRmOVtTygV5vBSLMiExMhzGrjAaFYYpc1gQXM+JwtXfGep1SqYt3QJbmZY91VWwC5hFJhsLyOpiP
DXwemNkz3Sgi1JkhWIJ79+ZUkLxzlzElt4tuYxiF++GbbzTmc12BjNwy2HDcZGoal4kEGuWdh/Qh
1Tmb6codT9c8Ub3+7RA3jDx1QHbvUneThxq8JWJXjyF6sYwgcULeVecErssaC+XpVfgDOe3ch7F8
MEMYL/NjpOmVutPzNlxmsudeAWoX0Xhqoig/X3+407JWdqJAQkemJdSgSHj96edLdc/HoWWqEWuq
nlNWhDX7yW1KNdD68MZU2xR63FGrCir0fhViEabzUAUCVVMQYzC2T6Ge+VwRfEaqWvC5RR/AA3OG
ZhTJzH3on7b9I3dWykvRAyWZCkF71+guDFCho91rVNQEBMGSfhdu3c4FCaUnzfA+vdCLCTSmQUum
t0RbhlbR66sYRjKrRP+8Noc8Qcc2LyfL0KFmyvF5dqDpNksE2C0X91GWfqqvtfXJT4A4gjpZgcFT
bAxPyTlQVnQ89Yw8jMWGjaEBS0pJc+eMZctbyQQfEOL0+WzfSJolzfpsnRr34kjL/wZ1pdSLqNY8
U4pri1PpaDK6xO2TCGQYUJQd4pVgEb+tunP2jUcGKg/v7njwAXYUvOz3sMjQ9K+j3VG1TxS8NwFh
cQis2tBfOzPfHbD41yY80yhAAJ/lNgVFtEf13MDYJ70vMhw3H97gE2usNDKsed+RrD3c6G84/a+I
9vTkKdEVxCXcV/GGUTkHggLTanL8+diO0JBxBFz24GkmGmqSbSXEogN6sEEBOTiHmZA3dzWIg0dm
MIVTzjCKlOFLAZuMhqBLHzkT6yc5WFmi8slPM2zGl4clmxeIKlLHY9kZEXK3vTFcworGri70wKfk
MSvKnisWl/tUF5M9GYlB+31561QRR70cbtBf9Gl3BcHPUlCM698PVkUdOxf+zDGYNHvf4+ijSdc3
3E2RBG4QOUubN11wHpmkbAoQqUwuY/SkTc7buTv/jtONyx8yw/LXyvW+mjkwDjIDBbz/B4tnIw/1
eWIg8t5Yjdtvk+QiRCT8yU5GS2HUIXMGRanl4i28Y+TG9NSiW5vialkHtDdsHAeNiNmLGx7v3JoZ
+gqRWnGvpKygwaO//AVGxf23mbchgrWljaBQ0yTCpNUtJFeDurHDA73Ymj+cD467YZPGWVLoTKSV
9Y6OmsLn5pwH4WjBw3BiCwYK2oDLpI888RrIxBiQj1e7C1JCJLgaCfmSVrBQ/H3KTAJBseOySnQ8
vnpSNWReK5jJ/mSVxHEGlvG/MCeMyCU7NJj+CHULARXv1aptcPTVNK3LJLJkRoA4wBfrvjpciwbk
xToswE5oIVFAv3eStAWbnVftqOs85FY9vehsjqjzwspx3l7O4KiEVo28fE6PVPXRcSmz58QDwgfl
Qsaai++4+kbinxEbEFzNHMOxMZF0I0ICh7k6jxdY2P5TCdlCrFicLD4Vkr274xsTnDaXRPj5kHs5
Xf5ixL793eS973xkQ15c4aJYRkxEnvGFhXy79tB1JAAzF7gxv/3Yd+Y/St+guniGwhKMgtCAnN82
1P4ZP6m6a5SPDJGTfPy/mAck0gStU0ENkRReppJ41rA/+nte3rZrUTdM6rdr5RL+AXztdmnMzTMx
XBvn0gngWiVkhRMQdZtw7byE/b5++1Af9x+OpoQ4GGJfgQ0Nc570Ex9AWpzAIGyag1YNw/ru5RM8
KTI/UWDb+9Gvs+mWJbefufU0qIVYrd1iCPhvJTqzpU2U9wKtbsbyWpD/0JBmSJidGuuOo0cs+ItW
7n5ZujJm+t1v6VmAMADvhBSdtXf4exilC3RL5s/7PPrbaLHE004fPMr9yQ8Ne/EOvPYgl2Y5ftuK
zIL3f+XM3iyJJCSl9vZnOliIAvCbDK2LFrwnXvE6dL1o75wd+t5fRfL0whbn6NIeP4r2gaeUdIQo
R4LZvvU7QmvTVZmX2NBvd2t0Z3TWV+9UBjGigllArPWDJ0sqNzuYI2djPCW6nH41WBjUrfWHgN2/
ouH3ZY5S1iFQSMx9rFMfd7PuThX6IiaFSJ+Rx8uRDDcEZHAtgfz7ku2f0wGuDex2ujhMoQmDE+Aw
473TB9C2zIBbodklQ+m0WrnM06JWn5FETRrb7fFCF9xgy9FRqzB+Jsd1W6xyIzg3aFMXwynCPEub
eo6/VPcf3c/Ahw2FOVNyLRkE72MfTwlOT8pGP+s8ASMETzXYu6YCxAmEm8bnX4w4J6UuFR+HIVFE
eIR20cHQeh1NkFyCA6mFnXeVIU1+OGkQk6SCjD0PyzDFkWGxrcUa8ZRm4wyGWZtAQmQKozr129QQ
SQk0ynDsPyleHXtqSw2Jp6xwUtOoFcX34K/TVxgTbwUbTb2wE8cYMVeGSwrgLBVXGRppWEJMtljo
W3g1okw5kiHJaErujP+H/aXmZZa18MTPfGWNBQW75Xy23NbigtX3RFgpYDADJYIxv+IWUrPB1qqH
n/4RHo2x92cRjOO8EeKxLjWq9uN8R7k3fsYzVRg5KpVAogmcOuIeoN2USADwLbfoV+GedtqGk+wB
2UwkHhNBnXPmUB1l6nUIZoC9WnyrTjAp8TfWz4EBvmcqMqssvg8milJWuu41OUNRpBHH1KpnmPpG
ZWRQx3knxzjhcrnI8JYDibI8JvDk7CUgr5CnlBLlMGeMllABwfKrGHuYkcKdHkRNjIefnR2Hb6dc
dCJ4Y6EPbo3GI2cyfiyWioF+Qyctnr5FLuGMZ2aHIIVs2QfT3Ex+QXXsBh1JMdmqGY19NaapNVub
694wqZ3QQJxoENUSeWGdnfxVz+3GZmuHZib14TPjykqBmwL3Wpem3bhYKcfeqgjNM5tRsmNF0Te4
cUiF78mnu0U6qbbSE+41KEA511shUaeptDBhud4A6HIzoo/RnwgM+uC/4ciuG54tM9XALUeSbZkU
ElxDIYZ7d79pw8Cse5iTDxy/iJL4MzcCmYI1Lyqk6pRANhpztnKzKCrL5Kss7N9UfewULbujO3wr
yDUYEW+FsamFf1H3sctRJEhj1vpeYqHvBeSKlk34fMBtRyzQ6Zl9lSMwFFuLWbUmogBtzCMxdIJR
kvQmWmu0/mAf6qRMErWi6+Lvh0HKAMYcXCE0ETR3HxPOL9n3IuxEdsVNEJUwAr4OSramneT2lZP0
4ydIUIjw1sTRIQOS+3ATlcrcoq0yuYVRVsI7s3NQyqmlN7mXyVgAZyb6y69SsSSH+yLZ4nxkeulH
A4sd6JEQ2RugX+bwbe+wGp+OPGn37rVATlPV6XlfHXqOrDMvVND90r0Wt1WGXeR+YtZAw5cfxwQZ
aDrwsLeh0cvL1pzlHse6M64nqsjzqhHEZfJfihIYOnfJ9190bxuwDQbdHqgA3Q4pcW/Fj0285Zky
OwFHUdEudXJ6Xo8JDpfC7y26X1YqcdgVGghcy+DVflpE/JFdug2dOml+10jlf6qpb8zoPZAFuqet
zCbjMSZAkd4Fhte2i3BIxtyo66KuSo0GoEObT30voam6rseKAhJQaUBtJmhSyVa8eKgaI9MaGqCC
KStUGIkqq7O6/Aq2FfJuy2p6PUGpda0U0yK9TWrHfEFqbnG3rdyx+gY30PAiUmHZrcvT5YbKMMC0
ojAoZFYpq1bySxCJPFJwU9ARzcBrdG6ROMjmrUZsP3L5wiUunBbbmID5ELkjcYDHIGdJOMe62LPK
z4DDsmLDeBk5b5e+W/8OhCp7Kqr0xrBvt9MfQKDbcYIzXd6ZMOuLZwW0oYJ2t1Cnm6QpgVRPnVnX
1CGbSxmmBaIeRtbvPNwaNal/3dAuXGVpgRiEXU1B/XJ35+wuB8shTyHJkYp3ZGJg2WtnIynsqj3K
rY4+yXG1d6a6/ekyQ7jvAPpLxi0V5CNHCKh5eGBkWLmQaeF3k8vSI+4hSZii93zIr/+0X4DySQ7p
F6IHR5KqQeND+es2HCp6w7OrkrYcoHeZ/WrZf2KuUAf9443pC7DBc3Pfzvu1u+OK079YILNuzjwe
Do08rfGOvhP6QDc0UZtZngaJ6CoL7QFvCyAuJANw57JmgWpM/0qDuWbK4pM/zxN01IyAGiRqPPpe
eL16vB+rT2/skIwf5ILPD6xi5Pe0Yfx1UwP4XVcqFbN3dW7Hf1NW5EoKmPuqSXAPLaPVW3c2qUrB
jUST/8Z9l6/RqcdPjJV6tnhN5jW9ey6GOapuvNNCRM5zbXxrproowJjpVueeWSXRf56X5kHIx/rM
Dx7FyuAByVgRBUW6JQQI2brvh4Kak/1iMFGglyErwcgmBsbKrC3A95s9v5qxwcq03ktulaMB2hil
bJY+4mwMCXqIgbiGPpDzymb5QBYlmK1kKiVeZCoc1Zcfkd+ZfaZd4I1544wyMzPcqnb9Ukls1Nvo
1BVvUl7hB9V10Gq5pI9iM7HmxRjIWpB05PKp+PTV2/MgbnvP7IqwmK2lEO223S5WokfXhCKVIMzh
cvY2+WC2xcHRXAqRmXjJk5owY6jSxJvpQ5RyRRzdS2tq+G+n54q0bC4oHxz+gMxuXNnD9VCCeKxw
+N41q06CgjS4BoTUVsnzGBa3mcdvnyI+bJU8sqd6tlcC/y2djqWTcvn9rVAByTXZiL/2C9+2okog
H1gManj6myTCcLt18tjyfbwsB2HFKMBzq639ucpic8LPSZyiZ2zeVCtsTwnSXiyvvMpIgnMqHW0P
JWkUjXTnps4Rg5mxUETYJAKPvnrtv1G9pfWCUYpuXWo7JEoDARXk4RpI0hQ8l3rlyFRwVxrw4ArF
pT9U6icAwos5Qu/uvNqLX1Ouy7o5EinqwiPPyJcwql2kwd4hULtU+QJA00dni+kR5c5/1igiD+1K
sPll50uiIhH6egROwEpiABerRI8LvIlMVNSkdcG46jjv/NMwUFrR6u0wfRqIVPBZ+4yejR/2a9pN
aLdYkAzw/+bpb/ysAtMEutDmbnXFaXZFzX8CDz2T2IzVzOHmBF2X3QB+9goh9ABighpS5H+ALkDN
3NTEPpaHcK2ULZWt1mXokShasxr5z0k5eqMj+mW8td0Y6rQUtlZ/D5IwON2Cc5Q91vmDgNjwjSxk
fhuZjEAcdpcpDmC6Ja9r4wBTO5tAJY8MIlnXFInK6Reg1Sic62b6JdMO9w9d+9hRI80ZkuV+CD6n
nLHu6/uhYDw08vrPKjimmkz2HcEuLArrzbkn+82wNpHjgs+M1K6CgmjPtKO1HxpRXLPPqnEZfpUL
0PSdLgXfoFRbFKFUZmDE64lcJkLNHINh1C3h1bVgsSQTcOYKcVKuR+q1PRcoeZkC7MwPdbu2j5La
uwjfRpcn/1GaY68ijgRx65VskBhAzxeUXbyRYkc+GZE3aBvXYSr0e/CkiTlh8lKnLVuqeBZbO1EX
WR863+7JkWYIPI8JU0YBkp6CBYqJii8++PYWes18Il16mGfbtzvDlOfZ2wrxJ9KUXQBqJilxaYXM
0+cmMZ/FgryhRZs4ngkQL1Eq92e0Jha3Jc21pXLyLDu1qNRonAHbpU21tAEgSleukjBOE6e/iAEJ
hrukPnTtiVbOlrSsDpTGWnVhHEYsgVSEsjzK7QWaZHfN8XNAEu4UW+gHYIccvoz/lIeSbjoze53X
Sbs7u/AGllIIdS3SSp/YmniM6tRbP7sUv6DvkBO0yHKitmrnWpNRaBF2ZRZpUIxLD5D5vb9eupiS
4iHyezY9f7xS9r4KEIUijGw+kFYZJjqkpotud+sArR5PRxx19TkcUo1GbwQKOVQTSa2evvHZQWlG
CojMc7D2tnJGzuv8lPr9ag3xGOwuItnwh94Dm1j3VK73e1FVdj/AFVM0S0+bBRN8BVaiuKtbIzON
k4L7IZ36RJxxpcwSP/rEbfFf9wB/bPl0rcA0mIZJulEqMRRXBUCjr/lBAQwGolKRztrwoRj7uedf
iMCxjPYODLjs/QiQSsYThf3SjqRM3oFCeeXcmVWkaHSX/dkMTQ1fKcUKJZh/GT92AGVA/BJ5IYNO
ZqCSenOJlElBWek8ZITP0ZGrU0DdrlFxw/h6SoK4tfLBfnBC9FMFNQhkTwf4JaYEpiNipg/kfUpw
Atgi3K+5IzBTA3BgLoen4+XOWU8PJp2rNBWhtDvPX6XzE1tiaeZEuVzclLA8nNxFOMVXwVtq8+Kd
L3gfakC4rdk7Mc4DArL2JMZ0X8JbS9Wydf3YNvGwZv9QOjMqRMp9LhEN3//hUcd10ZUnXZ/VdwUm
HcBJiaB+mTMFjt1GRKp90LmUG+v+hM2+2A7382rQQNT0I6YLd529S75pHsVRCqQLitOGE80dUNWl
8kGEXlxtXhxHT48tvO+q1KEataabCIu81WgfWh9IDO19CQhPiIE3/R3h2DIFTrG81Gps5b9ILJLN
yQ9f11VWg7rp/fAl3PQB8n8/1zCoBptvk02/CtOXgTPs8lupl7BRV+kIohkjJwbnjHL9ULghZbJ1
DcBo9FHAQTvO68294UxQjvUqptkNYGeIYGlrwgPIPZesvZ4nKU9WTKE+/8CgyhDIDQh3pLgkyJPr
M3owsmmyADt+p/HinMZgNed3jL23luqV9hLYSPafQW2TkDqi2QgnBNQFbCyboDNXrO6YA5h6GOOm
0uCpmQli/IqipvsKb4Wdvw0p9b6AkAb2cV5BzlYgnPtNYcknnya6Q14V3MSS2bCWIqWwrUKZgBJx
LiWVc7H9EiGodUIqbYQNOzfd7m0c94eGX6MxcXMCTtcpPCXMvbgQYHTspbAnssF66XYLbaWGSDeB
od21Aa0r+L5+ZyBcJjdsGFt0woqrIbMjW41JKHp9aUSvyNJSpG94QgE03LlFNDsG1TehoP4hMt/t
/St4MgmGwupjYeUCwZcIRJia1le94vcUQXK2y+InqFrERZXpfZ9lcgbEnfzl6JuSGYf6SQ2MwECb
JpI3W5U0CjePR0r6CUaPYF/oVNiVNnBe7TKEUqzvdXY2K4TzKmKkRDDgHGphY2ALiF09Mf9NavW/
PHxW8eUf/UX2wwgx6CkF4Id2+vZ2kM+BJOkdr3s8bXRsG3LZOtXxXC8pAuovanpw+hc0Tg32VXzd
ULEh6SM2EJ4iK58tsw61zsyRz6LHYxGwLpnCp43HihLu0rleKiDKTTjbf0KV5xpVxz6LOBbublQ2
YkBdtHzSuI2plaAceRwbyesZCU65tnlXpfdha0bsMD4zYuD3a4Aofd3reJpFVNanWPm2g1Dcd20Q
VYjGNBZ4lzl/EYfi2sO3VND5hsIJmGpxqBH1kgiVrYnrkDyiCFXpSM+58stDHxIEMtMSxrdo6keF
PRm3evbKdbP2ufYMrXfuD6XBXuaGj0SV9g+gaU5OZOPPZ4sg4+ZvS3Oyi3J+1wafMLkhM04whQNq
r+2E284O4p51rm1tazx6XrV7ekHbpj/EWPw+P9dr4We678+HBn447pWXBLhw+ZKHsJgyP+DHfF+K
UTuLP5wxNnz3duYrmn8pqcwqJcz0PfDs1Cp4BEZWWl6cyXvmNmwp2issrK0iqowQ1fSgTxrb+VSF
xcRdIKaalt8uXCTVyBXJv1+5jjrGkMWX7Ye4yg4gsbUmMzZW+YjAnfMePgBG4XThviHjm59reQ9u
lorV3Agei+YzCERebF3QGVH07D5oYJM4PDyXvurZfEkxiDPCeXIOW6YoMdcF3uZ3P4GukJDNW3aH
2CLCdaY10azwcrcPmdjBGVLK8uOSWglLY7PBRQRBiIy/rD1oakOzdvxDSAJ56mBmzLqlIR4Tis8e
Rd7l13+9to+lhcIGIfC4dHGZBgd965awp0UqLxDFEmJyeDNPiO0u4t9ScAdRg4kHIwyCPoZZdbjB
uCEBpmK1+4gth/LIlfZPS2qGpT81GgF7NL7XuwbBuaJMbOeF2m51M6e+VjccXXv0UJmd0wqLLabg
JnMu8VCceCcXSqqpIYt2vAIZkhd9MwWvOF3wFvmBBWqlHaj3kCrw12V0s2lSrsELYDdwOXQ/SDnE
nTtLqj4NffEtZLTmNA21yHBUFAlEBMGu271VzDAuvYySMbXnvvdQGoKiAQ+7hgkVoaECVnRp5/QM
3mxE6vfAkdc2qiCcoKZDNDP4U4hI36zPY6RlJHwNeFuj2EEDtJgL6Zb44s73ySna6uFvhnzH8Zn9
W/spZqDEomO4aRG84Xcnkd8fZS8XHVesJmLxUPNFVig6OB/A7ZfX3I+FUJwR/YZwFodnsCOHQbA4
w3LbttLC7RL70xhxNtAZz/lAiLyJyeLAAFi3UIfui2vfrUt8YcLmFAZi1WvHh6c6GO9UFGj868Em
apme2ykqUUID3FPRZOzfBzdhJnD0gS44YUs1a1x8eDzlfbcZ8RW7MTOAlUGVxyotaKgybRZJ3KFb
1gx9msK0mU00KBhSLuoqpePoUcbu4pNxshiWEosLkbXC8P6TpjcVak07baKtPUv0oxj4iQQBYla1
vrK/i1RYZkt1I0xxCxftTpAaXEfeD64T3czr0z8z2f5xV1m9soSq2XVZly0HHti0SLlApjJIfOQw
m+cgkwUWNof2aKTQ+0uCXmc3S8Cr2F1fjDIZY0lgLh3Fv3m4LVEF7rwjX2205YSgcddKOQgoi3jn
xBj+tzTsR9Xc2fXKF7S6Mu048qwYyPZsvXvlJwfDXJTTXE3z6S8vTSZgAdLU6sglIBXiE+AdK+kl
nOllC45oZP78xibFLU0XVEBE3JvbaaexwvagcMA03GVLescvapJ8gCt9TVBEDOhkFVDpWjkoKaUs
K3KouNWajkq7Gygfml5rHjbiEDah98Cbb0fnD6zIGP2kIt2LLU3dTx5gN3Nsnp7lEb5KfQncwQ66
Lxme9e3EVGIyBvKZJ1WOzeve+e4cePFBYCLk5W/Mo/wU/AENKpZJLL88qUa8G6i3tTecx2orgCcD
eUxsWkS19ENDUClLmq3AtnIwFF9Cy32+43M/wysXWOLWn/W4vYBebFFIr8GEOFBSnvViU099en8S
4t6eSa5D77BnvaJPG3sXXvui94FwaUIYzB1qRaeO6Lfa3LIPSWun5DOozBUiu3lt66h9n3tgbxEA
svExAySwdjjaa2+YJn/s2wKFJMBwZutAwtggOD/3sh4L5Qvmaw6BXuwfauN3dyY4UzFdJQQ2/lKx
qofwvJxlbVPL5zNCOTWbTeAEj1SF7Be+31MCOVX+UCWLLpSoERgrnFgznDLnqae4dWsfw5e59sZM
K8pirKCWFoVWbAnCTAmh5bT802JCcmYPaFxH7YkyJgQRUOpcUTyF3/9nCjTu/8rKfBqOaLWP4DQp
/53TI8+WCDrDZORJK1/wLHE6zKm1jsPAjgTra7oUrSC0KpsPSTT2fMATsRctu7s+4qdUm+aOYMxp
EnnjHWipF4Y5qqa5BNj4LZc4OTSTCPoAvA5S/sQ0cxPPcLejDgWY/y8QVAP/WaH5jAiJ8Q3zGSGI
vnk/ggqwAyil5fZpcJ6YNuTheNtSE+VKb7aacfeayWqKX+DBhg64fxgs7LUoI5BxGp3LTIg/Lzz7
Wt025IYPdHhO2Y9frioOJ8zZX138ruq+qdWciMcHmMFLC9Y8rJvO82CEHofh9wk1R8OMez6u7oNB
rbElMbBIUu5gsUCWxqqS2FZ510/OheeZdIUK8O4jea7IRkGZ8GEzeHQsUGy6YKu/knk8aryGgfdV
d5WXlPRH2N8TovmJyNjxumOKZFsbUGRhgsfY19M2r41mQVP93vyUFVNwM6aoLAtELek3z+V2dnTV
ySpQBVEU36ERzkMwvIN5VgXLxy0weVKQ9XBn7/4BPG95/BOfxQ1ykt3le/sjGRnpnLmcHZPRzxTj
pWKZ+32EwOrzTXSboNOxIxSDqvHjOLrM4QZuG0XlA4F6fv3dObA86tzJ0zqXFP7ldXVub7CYSRSU
ktcfP+seUewGqtipphuB33ybXfowycAg5THIgir0A/dSNSgSr/u8VUCw2MnvykwLl1+huVlkm6wT
N0V3Vja6XVQGNCaS7c0ZHpoNhbQtvf59ZSdLUiJ18m1BdlUpH60aqaVvm/opLhmueN5rHzpXOphO
XP1plXTH3qz2YrsxxX8IaZ+Q5jXTv0aIGBKOsjh9tk1kqUY+R/E+M+J+nBr2jfOXtiFw3ZYCZb2W
5TuN6F/3q0AqXktnmUXNNu7CeX1XCvZfi9eoBy3p9L3bbNcgGlMDYt72OSqEbhsAD4uS9FrwADFA
r2zk5brkFBtp8dkz5unskrF+DWyjpow/NIGxRjGvGh7JKYTmv0cmtDBa2YJAQOEN12qQ6VS4WIB4
DRS/YwVf+64GD9vuziEFoWt0fw8QHpOmmJfUfXodWakBnHovt3dUvsUp4hm+y4zs9VvZRh2YWVxj
J1A+EKMbflYR58pKEyk22YpVA/eBzu2pKkbe69kL+aFfxJNmuwZi6zCtMWeo+mUkxILknmLEIhKb
M8IW7r4GxkWVCX+lEQ6KtnjrTudpgDsPr8RZw68XvtzMGPf1mqbxlKIIQS2JHeHOWvRs2g1m7JxB
n8fdsEGplYCzKnrUDUu++1bdcgleSPx/Vd6AT9Rs7tQyldJBC1hKC1kdlO8D563bvHUU0Ex9UCfS
nV6Bpu4k7dfAlqRUR5oxOufINA/cfsYPY6sq6RdsuwiaG6Aa4vIoHXFZHTK5OJ8GJpuBlqqGUpcd
NHJxVDnJvVZRCRV9th30HH1ryFLjVeLtOa6LVpi1aH609qPrMuKmyVqGMxYzatjKC1eQTji3A96m
n/MnBBzq5NnLr0zoOkdnTyymHOiZdyB1giIskTikBah9ysV07aho5bjEI/Xqyb7zGcWvXaU+KN9d
5VSU6x5nPXO/QL/kDmfylmAE0ArPvXml0Ez66LbuCi8Mos5RlNmo/EKDCKUoaccJdUkx/xMD/bev
AZfP662VfSRZNb9064Xnh0rvkye9k+3wA8rSQYiKfRCc8K1kBRyd9Oj0N6x3cLHdq3WNDODzhtxj
ISqC071tY6HO0dQTW2YYP0H2ZX1nUiM0a1R2LryN2gnTf/3HTKTFW+xnVtyRqBhyUg2+rD+t3dh/
I9oxlxX5I9i7GqtMcEvIglyNGU99q5jHV2LRhp82mig3ALoscROQq8vR0/SQj/i3NBzsXgeIN7r2
yIZIaOZjdUOO8deR/g1aX4HeYjsZXszijtxrS7PyfoBbhA+buZ+pyMQXw1T/60zKltLLCNngsfJ/
E6CAYwHJKMuZiLpF6lgqlBEXnaM2r3XELPKIEVFOMUehwITdr3hx/3SN/N8Mkk8vd78QgKrC2p0P
qMwU1SyZbvNeGFj7icekyb354l1DmajsxrR1M3w1xN5gGgut/99wNVDkElD9ZvbgeuWfGOzTCURn
JOuvoqmwQnHWOEbnMvamz+fBkF+ovvjhVfEFRDGAEv+hFo6NahfbkIA6mmJQQ1BjqXBbI41LCw0D
T9NPF4KSxecK0vTj4mlDalwPv0NqOYoNIAZkpwCnuA5Ssi+WekaUZ63n8qaxBtccdoJYiz+G/u+r
+y4xzIgKJGhuTdU5rNuFTRtOzex/Ki7Ijoy073bUCxkhjAcXs3SPxJICubvpCuQDo3h1vMBxzyTY
zueViWRaTGqLZiRDjTISS9I+xwA3lDzgCjE/8Upx/hVTIBunYxSS7/yyqhPF46wyDz6Lovd/BeEb
5XEIz/HEQvZKCI0I4ovGVN3fdiBOLaHZ2V5aMsPvIYQ6OsUIQVgrdHV0WMG+5f+xXBdqhkAOf0Hy
D8qmHe+tZqgeGLl5UNDqjFbHkDlA2UCS7vwm+hQmDkQesgQFSvWh4iIY/USh9kqFOGBs8ErW/JQu
yj9XeSIudhywESjJc2uuglzDNsa6eog8xOUz5WLMqHAz+goVQF0i1o5CQqeI6mm759bGWdaGauO0
qnneCbIbZjt8vhDmvx+RuK/ec716wRTQWW6t8cJ0L111ijGmQbxQXY4nPzl7PWPzbbX4AfFRiqyJ
gt3cvT56nGsaPBgYT6kJhjgns0rVzm41bamj+RkJfkjLaVokgZ0j6WML2gnBtvTGO93CTriUBMXE
xMpxvAcPAKFLPhZTQhoFI6CkOr+qdAqjbOhKvWDG/BlkDcBUUAdNnbhAUUaO4D86V1BJrfvLrLMY
LEkNhBS55GIfryUtLNAtz8Hi06zGbDFPkng1D5DXwgt3Ug12SppQLz70Hzc4eWtvJf7fh/4e67sr
b7S/+vWkWGg4Sxsuzup2LmCgO6k8ehZXEIpioQCp9lr+Gl4gOPUF1uVN+IHkFoU6WzjO8IbRwcGk
625imUePJddRaeB5ufgKvjQ52fhv/wI3sbeOS1hzTGUBa/cDPsLgoh/iPz5JCw6j4yyFEnYXKkEf
Df60d4GfpIYSMqUna/HDuW3NPqhYGFqIchKnYYQJNCm3eo3FUCgmWDSyvN+WTrUDsZkjwZ8RPz4j
EoqpsP4VsU7whE64rQVcrXTP6+h1IelkprUyQI2Rwsn3e3XUQlExWVCP23pJQvhgExj6PaohWNa1
RELWr3eec1V919JrwAaVrplsxeCQ2M3WDvEV4LvGC9A5Q6BTPtZkjjdeDizyPX1HUJR68hisS/cm
+J//mX97CdQ1gohEmZL+l3raIzEoaHjYwPG28cg2Nnwd32LV1WlAp6LrN/GzjgyYmRytSyHmsUx4
PkDkOCBptVcy45aDoQq5KKO/uYx6iEwnIeQRwddqynjSqXiXWn4mnLhKv5Qb0JyLj975hOs8CV8O
LvKQa7zYLVm/Z7G3mYlt03DJAiz7hqnSZt/76B8/B+6Klc8mGkYGeuIaKi74SHy83aWFUCmGIvsH
bq5AgR1ACUWiPTO6PiOavXGOsyv+0KKWcmJnSHERLHzx//cH7ESzPtL47ucgtm2bibLdWSEKjsCw
vsgSz6mnh348S3tV8tMgwOUgAUWK5Ds3aBiq79ZduEAYna9bhHp+il+qeD2Un9ZFr/OOjMIePovd
nAR0zBnHzRgeivdxtaiUblMsF33w3lRa0GepnvcBNDWHS3g/GN41TaJXub/SyUJP58KcdgkBPxWg
gjZTZWA4FSPtkMe6rrz82WCB783kiYHfpp6jVXvf8AAQ+hdb4dAGxBHZp1USQlY9N8NGP7EGoKie
EVmKr04r/Cfx5EpYQIvSik2VS3/tRFyRu6crVDMez9YxyGEB4i9DGa5DLX2e6zfcs+xzTdC6B150
BhznUTPihJaHacE7onRECN3RTfXiLuUdTOisPRC/2fmHtrIsEtS4kgG8ozQx36XmnmwIhJa9xOA3
vJAe68sjnHZPxwZChuQ9e9GSrMr+jqK5qJiVjYxf++DjmeaRsFDnIvJYJFzVhS0I4FaszEzj1W+S
Kf8CDcxVGJm7iSrzGmgx4fL0+hLgdGKxz1T5q57pkNHU79yCHT+/XEq+o9KvEjTHPxVMJlv6Rls8
SdE7qRQFy4kI0bzBUMcdrz/5krPTBvx+gi5FM7avWFaNKH2rPh6BPjcf0IXC1ybfIfXEyp5syhTw
gB5LOLI6DNrueuw2lrHdIGL8l/JMIduFlibhu/QEKMNOneWTvJ17FmXKrujx9E4sEKybFGnajMnh
3toTCfL1NX398isa146xLuA5eyzujsvQFKZ2RNXb5ndv/ZPM/DUSouu9+obfAjt91JtkBMNABHIJ
tujyjkwFjBtAoSqyR3JoQTGl7hgylAnM8Cw+4SHO6Cks43KTuq5UMxXroCLNZ9IdtaU1uOwv6hs2
HGGbU3j8LgJog+bN3thOhBcePYfFDEEjm2+q0AwvB6jjh0IYfow1up38cGxIlmUhyFqMXZB3qooy
rcdt9laks9yIUD8Jpt/Zry1xZ06ON7oABqFgHZ6A9Vc1CmFXowci/kCusM4N/ESfCC9oCnr9241P
iovr0QAb7m/+I1J544fuanB6ecWsoqR9kxUu9uNBjH+ZRL8TJNaLM7yuESHBdL3CKfetzfW3qkSO
yQSCKNaDIqrZv88vpW5Sd+ijphn7gOl/cVDrPKzQG3aHfti/xbqpJE3W/+WvTZIZkm1/+3e74fBf
NYcCdtMd3VTfSsBZAPYDub491IdbpKh+uPcBJkkrXX/Eh3JHM/UGJzr7oIJ8TJdKa5qLdmn3PbVF
v6DfIZF6z703npSi6cA9QRaQB0cPSkVwexvO5vQuVFxlG9Ev6A9gegBtb4chPhjStaPo2gQXcyFS
++pMxB+21UlwUic+Us80EPqMnD6+9XOWH4u94bfpYqBgZ4ETDGJfpNUVo4nura97tNoRzl1Scguw
9JgTbQVEOvG1fWpsf0MTg4HvuR8AWH0C1usxdiZ19fEvlGCTZfTCxTZBZIxgjRxUwQDu01OWu0iN
0xa8Oa6dn54iZBFnlK4rdCu3n1RS6TA+2vrzc/e1zGfsVVGM0/xcgcocyms0J0gNerHWUt8R4e8s
LK9qnH6bbTHlI1/t+RLy4hPqeoulCqa/fyD4UNuaGaypx9NxLzj/aBt3KR9gmAwVh8ssW5ePoeZv
ZeiaBR8u3DZAyOFMCjUTT5oq3UI+GruOydmuWlZGHemDW6aa3Frr6KTliwagPQ4xbmWV56Y30rpp
I4rgS233Hbvcx2cY/jiBjEHqILefm2JxGDwAQoHvnUjBu83kmKMQxCy1sw1tEgli54i+MKtjkBzq
bgori4c0Aw4rGdIWAhBul3/50mQR7MQynpZ/sp2YRpOjWaVS+9S9WWB6a0rnAr47rLgqo6LmvEcy
SHvvCLadH+YeUp5024hqkZZA231aeS5/YPXJ0hYyq4Rt/qgwG0yTt96eUjdxDpH8oKWD9BUIOd5I
Hk2VCK+96VSOPhdX27q1bwJwfcRFLC7MB4t3tMan2nl6Tg0P6m0TlODYKCQyJSufi77vorOwMuzf
RmNx4BCBtbvJwRnXnJeCX68v3Q6NytGRbs6VdyLzBuvLi8KJCyKuxsT0fnGYC8bUSWZq09skULFa
hYV6HYpJOlliB5asp80B3Ig7WXWCiXwR+ETNBuBOLdAJyUimBJf2qB09hIUOsJA61SOdhgs5GOzZ
9ovyOVmDZ/qZOWxrIEPmXCr3y/gjM6djRsRdaTbriRESf9VgRD5bP+qVU0ZNjruli/BamKvuDK+x
GWCAT7z/hh6g47CWZTh9HkiCQEG6R1An5iIw1SD1NedC1DF8/Yl8aWIUtS6Q5r9CYTp2O23bnISN
M4KYEDiMGUimBmqVaEsvMpH6TAnug33AieE5fVQRkShVOPFKfOtSAVbPqPLj6cjsUSsliLyMf/N7
/vxnMGjMewAGEELCcytjiR2io5ev0HmZhWzk1+6pMCW2LH56xB6yYP4RJVktLlQT/GRP+KNUN9lT
BcDWwB7cK1I+CfQRJI8w65p4B0dKOCrXIlve7TjOp1ntEDHhO0lYdAZiTnVNqFotE1MHZ2k2e+cT
s3AhlW97t2AgVubRQBk5OqPpEoX95bbRRQomETbFvMOiW/qb1x1E9SlJfN6OUhtDE6R/MaFvzwka
f+daxk99mVcBCRkzgD5oZVuimhqWvDyakzGvf4lPfvuERWPT3b8pSYW/A2WfPFpvpflI2wKnIlLV
fzG+xRBBuMVXNSbxTqGWBW59CCZ4+qomhjG/JL1BfsB5nwPY5nX2bHsH0bHGHEW3qwvYWcNxxzua
vLyq+DwbKcqBT4Mrva6fxYCIM35EImb8yjobHxSdxxMHf9URsWsPaPyiGojYDmlDy0w7z6HSGrWM
RoDztRW/Rz1bTn2/x9A2y4/RbSYYGB5ibmFF8I1JwKLapTgASCJGTGQf6xvPePo9id1kMgOBFuH4
+muwDDRaN0g2Q56vtN/DxUUxNINC5P7atjt3n9wzDnw0q9SAUYEEJQ+FLfeCxidw/hjjUlZjRlhk
HK7J0eQKHhC8k7bRBw9MtzDVCBTmpGnNeNsM1eqnObd6ZQcCK4KX1kvUyVqczpDixSd+CvR2Hm/Z
Hc211QvsB5voxww+zXGe9W7yQlUu+C0q9z3wP5m2XaFFW6NudU/oqAJ1MX2yLQA1hOd3X60hH8KY
hk+C3SM8o8oJ5mizQMV45hTzdtrQdO0Ik7rckHADHwnq5w4RKUbw/9uWB9wEAdHIZrS6qZYR5pUm
cbks2M0w7iCBLOXWVUio3+rmQY3S3RzLoZ6mxwA8+lv3DGofRXAra2y0EfsS1MjUeJ2EGKRXvV/j
C3vcv98YQtXNUTD9s9YEaxfvFnxEqttajHMJnZPKcbhFO191IQ1rc0CshM68KB2w9SXsp6Go1+6R
7VfGnW3v1cE/Z28GUYxr5FeXgO4OgsbVAucnKciXuAy9sj+9C3/1v0fA4aqhuEeLw2m0eJIuggye
8u9fRuiMb0kz28N01E9RXvrWerWuTY6OdrefIBrE34hFsYKKlXu+96b0ufyZt4epAT8da8gIMQsh
R01VfDknUv3Fw/Tcsyo8+hBkKjksk9brf1TmA1QOkl21QJWSS8qyrhmr4se5vqD7ZRfR9Or1PKNa
+2GduzPR3g0WF4OrFbWLhnL6kcFgS+jE5tRYKutYOno9jYC8FcFeFZUuKK1gECjDAKImkqZsaTQW
0c/mi4yjyezQIQ9OewBcYci+H0UWs4NjU5zsj/1cOoEWQktmjTcbvGyc4c2EhQo4O8WGzhpEZr7Q
Y7/aVizpsrK9AmVQoqS8t7ESUZWbnGHihKxqRLeiTuvjRAhumHTyxNqPmSkWPmLSxYgDaogsjm4y
rAaEm8I7eLtEJgUmDZ80m/sISYY0yclMt6jIjqrCR17jP7E909qQEwM4TXJYrrv5Uy63bWM7TpKp
FvlxLmcn45g9A3aoKFm80NhcGkQGJRN+t0L6nyq4uKqXaw/slprcjsmXFTq8Adh/WsY0atn9fokb
TJ7LO2GH3sgc6MzBxG8KJUEA1LJhnZ2cPJdnX/XeCyB43G1URShjrU+bnMow9fRZBtQ1J8HBuZyH
LStmK7SwodtJ5prq32bqU8cFJI08iFjPtXvDSq3isoYncomIbBhhTOd8/HHxDCjl71b/S2A0J/gK
Eppw+GMoWIS9M/Rztl/a/t9BF/m9hfVEKtPGtKujJN/fYkeU6gZeu/VuxJRmsahf4+xgr7kPs/T9
A0acRqZYj5TyIklkFQTChQMb/bHfluy6uuV4xFTpxPZbSa0n3lxSAfHNFZBmtZiQN+AmK+b9p9Wt
Q2WocM1KgU8/wbI/SzcN0FFqk/u+jT3Vip/OgGQIJjvpmDvRuYaw94ylgSaRqf1HeoZckfHTTC4R
VanWO/qkOq2rzucOx63JQqFNBiKesGE2fD9hXmyoEsp2AHwDVxDKCDQXymoZFssvSMxXW7El0v95
0tZaXvAgzEQBuFsL+fMJYSjzZy52qNcGH3XwObeTegkyY5pvHMJ4jgy6Gz2qkvh6Y6ppzlVRBZgT
Tjz5L7Ou9w5st6OnPWZVslXkKjqirTEWdlxDfsIE3zsx0AS28wc4P6wDNyBGwRdlp1FK3sdO5vPe
apNYm7P2lu88t8Wj/Cq03tKMuaThmAaneArPZoofN+7phejXRwp1mv/81uYuoSmia52t35K19UVH
LVXN7mUWcgk5MxjEKz5tm9PmAn3L5gTUAXD2GpplNmZA75Fq9SezkDE23x8cuVjXHB4NzlP9eQjE
E1Wz6enjlxqIAUkUJKnEBCuxHpczY1jr26H5GfHf5J8rQz6QWmwfbiqGlnfrv85VU3PPLrrNgP4z
MUSbJoRCOQopwZ9eBWZbg37h2W/5UQi3Up7UP93U9iau/eK57G3Rje4Yv1Cd0EcxeTX9Hi6ciY5U
PKphKYhpa2qvBpWUIU+zOSt6G9Pbvtm9d86DJlIiBrUx8yYMO5TSP0vVD4nawubMHh4zkXoDSY3S
HOIOxxQzJwP+SYYC4tY00G18hgUOPOSJvMc5zdmRDsO8GEMKC1qq6DNs2cN3nI55/OkyVh1sWaw5
3Yd3+kxaWTk1BzC4FHXLYMpn82L84Uj+m+S5eFE3RKPD6BVJ6+BxsgxZMfFuroWqRGjo+Ovsw8Vi
oolsi3zVVlxgFlmtGssbh0wxFkLLdUeLwmylX8gi1Ks9/JTQkAtO5nbE7Qmg+dGrkVHnrAgQrB8Z
J2zs0k+JAyKoixOE2aNrkZ4GSpOE/TdaCYWl+IUMCyg9iEcwMNi77lYYLKQaWYYdnGhlg1578PA7
sJ8EgZE7pObUhXRaifIvNXtgOgce0fkcA3YAWxe2a6jipzrTCMiT1/CzyH+EdFkpWsW2YcY9W31g
ivOpBb4B9yHso0nA6po/JMjISaWIFCXIoVjC+R9qyG2aWkoe12wv6qZ8VPUbAntEzLR8uUEJ3H6x
dsV3rsvspdEPZ+mVIW9AC2h3+7rSk9nRMvIe3n8qPCeNVZvwue+hsWZuClnmSn1KzMrji/ZMcdz2
mfZSxwCTK/JoWw1fZZTu6RlDqJk6qibLXEuyq6OJaoxm7/B6itARoT1UkyDwe0c5pxC7NeqguV44
FQXf56Iky2hR2FtEIroAMZrYfVG+9X7bGvonc8/CXpn4UdXwdnY5O2RvusDqXZKnZF6T2aBl8/Al
2d8XzV5ZBnxvf1wvGY2JHcbNT/W8MtI40mud9IHicv2YsvG1f7/qlPIF3Ttez4Z0bAcOkVeIbjQ0
Zr0CMHd/OUMQNusmHYzUXVvuoKxkRlI/G93/sDn4H9CMm5wylIPVt/zzXLF5h0QTTC/2htMTVvTZ
VRVdfSYit/d52lXVRHBs0YS/JqGtKT//9lISbzwR0Oqc/y3/4xzQHTfi9vE/anKHjRiGNmfqYHEc
Hriu77GLEfGnyDTV6mRqRV7odBhn+QbKAVIlUt1pRZolSbakjagCVHS1VjYVVI12ezE/Y64WzQw/
eYO0T+zrpY5vfMBQrNPRLxX2tYG7VnFLKEhprU9WT57RP2i2g+VuHM4A+5ZSrlXSvazIWG7Pt8Gu
qgwft5DMe+jLSVojqrd9tlBtfmRy3tH+hIcuKdCDZg97FRJvHzr1Ziz7Yv5dEkVtw6Bxm6WoAE6D
qb5BYHjI4ycrHfkoDJpYME8RpSKBrpspMY7h7lcH0n4WGgr+yWO5nFp5VByfiKv/sVmUt3Ii2dgb
P6hjAY+vy+yG6xFOTyVtvDlkGbvleYFzmbKiGm91o+nSFxZ12LbKFUiwHJF6t4UpyNS/Jhw0j79c
uH2ox9GTQ63IwulHp1EztR/K/K9lVukNOvX1g0B/0nEcPPwH6ZW0uptM4MvOkcs6JpOCmfk8pyJk
p9tUEv98D+8RIsw75v50gowR5XlYWzNDKRM5/qm/UL0H/CeSBcsX2J/3tMWhpg0YXHFUQ7RzgOit
2UOXjznPlebM+K5Bg+LIQonbbp2SCT+ta4XnWjEzTTdzgSfbt9AX1cLFm/n7ZWHP09FtJ3JG3kgC
r2BAD3LrUj0+JqNCB0qjJYSojCrUNAdIzRNn0BRGAuENEL91UaTqilhRfrv4VlDpJgG6vJ8GmLUp
Hl/bQgD98NAgltZ6phCgz2UU0Dhf7j5Z5Vz3MSKH/CCLl4Tz/ko5oGrJCUKi6jS5Kf7z+xstD0LY
zWKe7Oj/fgLfC4SGEHc+WjUqc46/BpmheW4rvqVjPZqTD+ST0ptwcZlIoy9I5D7B2wXKPVOoEgAP
Ju0y45PYSTKJSCT0H1zQagyxd+RbmRSVW5A6NiS6RJ8PI0TKwFUXfZm4pQ7rPrjKzLp2u4mb0WBK
5kuK0Wc3FU5UxpKK7du2yZq4fhvnHWT8IDc8pNTlldne1Q8wXvBlkvxpo8m+S5vIyyfVoWGx0GM9
YKWPPVSEzfTJDqLoMDODSWnWCxEDYm9qc0rHoIIIMPLWyczC+vBe7lcSummlQu/UDfWj/T6goGSG
rJi6aP5j6GLO31zeKMakLFyBcAaV0Ct47fpUIXnNSVVw3mscaCUFhjGCZfgTPBZSHioQUQX1ia9+
J05eZiXMRnAX5BlPSJtetZeyT0eGt3i02Jd3jOb6qGtqyW1eYf+8BYVBYjw8cCV3nvgoiB72mtgE
l4L4r8Ky2HtfietmxdDbRA/1i96qt+okVEoetdm9EfHMNA0ldLyzl7AJM4jwtznFpVv5MwH4l+B5
E28AeL0g9TJ4SvVAG2gW6XPNMVe4j0b+bI39ziaPebeYTHgXxxoNnMcg9OQmmTT8V+uhIVMns0Iu
Thhp9dYRE4SmTcf3KYSbSvxMxN4x7ZMZ3YWGZ48c5XYMjy61F0AEgZnpxzXWksW1xZ399jxinzQC
bhO2fB3X6Vi+9B1mWz4F9eItJgPVp4TuagvYHpbxQpB6Hr+VHmYHYY5lxL6YzatAgp+OT2gwLTB3
1cmvvJb55Ou2ivWIhThfAfAsmQB40FZUBESsLqobftzYKZCwWzpUXG66KXsuzZMkiWi8PZkOeBHu
DRrGPuAJDygLMjuQapobemMUV5xw+KLKSvb6Y857EATT3qBdtzwVQAbF4hALBHo9ZVcSFLOcszcU
S/WzSTjT7PxDAsjLz6lDQDV+0uaconXLCcfhjVOko87J2VSixzUqrSNBQ0PZzbR2JgrZGtL0G7bk
ALrsnUFtwB+DRkS/cI1HDZHa6/RC6w7sRrWhZWm9e6GDLWv+SqvGnA6Hii1p/gwbZhotduO8dpMC
24oljlqzPYqLDrTT45wEaF4PQd42Tpa1h8O2PtMemom8OHiEc/qKBQEqTllf9cV/wv7a3mtKofyG
FkmMS+RHyTpfPGgoKw6z3wD6XhYGLco/s79UkpQkpEBELft/LIDxPe00D+ZhWmmeSu6VGg6NF/YT
PAYyUvXkF/zSa6OG/9eAbUH9yGjE2WIhZ3YnCzCub7a8aG/N7Wpt7BxKnOMRy0NaCB8oUJshrpt7
hDYDpnckyyN5svQ8Q3iSpiUzRa/iuYe7e8iVR5praWsgY/qLu7AJ18FZ1599WG0Urm9j5QPhe8Uf
AXXmPOeIolEzudSLu2s4hwToS92C0X6F7Q8dP35IPZuJldR0JSiuHn6diMo7/j2l3Pbx/sJGEo4i
TZPJbUZEHf5y1x8AJuVKA+nQ+CnamWe7yHUHBUsXY5MntX3sYJ/BAzlowiYmCT9Kryd2ftFxxeFP
gL4McfCxXRrZEtELPr4QpfTys+lTh9JGejywR2WueaDNAoZWMpPL2fItqD4R2MvKeQDovOs58Xr8
Tm/dOtPdF2LHLo6kanASdkM6A6nYgqvR23i7yd/ehthWd6vy8zcc9lCLfVmL3eE736o6QzgAh6n/
9MdfNjunZoli6Q1wqcCZZgRGIiZ4kXzkmPd5A0D94DYsa4DcMK+lf4pBx7a0wtVnydb8/OrBnN+Q
ojNBkbofEEjF17CD8qs75RopAt6HP7SCAYA/bCemFqDhuNxR/ywo59gIAfem0IMZlAua2yXKQX+s
OAMMF9UvBcAw1UhAn6uQjHCF875TXgAobGrqVO8YJh+vaJq6tvz7eOK08xwubgV9mzrF4zgLhTsY
naLs3I2L0Ha+uVeFPBHMXKelIkC6ZIwG4XmUW8qLoMX7391HSwAD4oXC/42Hvn/o8M7/A6Mjoof5
+oJDgXMy80nZohezAjd0i3/rcTiPQq1eIqR9812dOapM0uxsG6ijpbQgDrqaka/GGRel18SyDdvY
mpi/60B5t5f0VR9s5kksV2l9LOWR4iTTQlGaLMjx2Guf65TiFaHGmIGOKmPC3NFefnfStl2AlcGL
hO7yWp7WCznj8PxebxtTy2hx0XXrE48oEfNWmBGIM0R7rbdz6VqtjYbLlubWgWvt8ARn0NjzOH9d
K/NOreC27AarahMlifHD0Sv/QA8XpuJu668GmPr1/70NF/CUuCNG8mJPnZEAT5+rCwUqZGEMbDrt
YPh1zSvEs4WuVce9hjKwn6ZhNC/1cGcSsv3sONXjw9M1KgrQUWcc+JZ00BLsgQG3GIDHIGxkAXlK
9MYP8ky7PWTKzXX5MW8Ayn3TTI+ahykci/VCsFxnnt+MELGypyQvL6ZJTed9QGTs2QuIgDIwW4db
JFDUsoHO+4LWjN2k04tx0cikBcUy2CiTKQ5izEBRkvnM3VESqE84OB712VLTGBpLm7QmBvXQ9UtJ
DnkeWh/KdQfU3KgXwhGtypKs17af35tp9ej4KWU67Caqvab73vDxx1OL9yajsVgmCf7pbUxEyPju
CpgtbmjO6rlrzjdwd+7lN6I2Cp9cAqd1fauj6S4IfNkymBaia2ceaQxUBbHKcOqXaVCmgvSz/sMv
Q5rIxV2rmp1bSriXBEXKTaUiCCWBbMHZOdx45IggYrIbPaZfZUlL6NC8qfpSNtPCeTqDocv0W3Zi
u9vCmAAC7Ut7Kmgems+MYJ5vaM/08SwBvQokt24bnO822hBDEV30qnlRsPvIk9g/aU/l1kXNkLRd
nZBFVXg74x0dQxis16VYFJAbDl+7pZ/c7ktP9Vun4FkL14hTMINvw1fpGGiQ7QqPSRyqhfhb/gpd
XL044Mc6ttD22T32kGqlbtxeeT+wC0gwsnxRzb1OQPtPZH3acLVef1JDDYBDcxltkI11aeDL2oho
LmJYOSExqioyCxFqHNSnfxOTOGsv3IkaLUp0+xtgIySMvzWVlelX5MW7lltmEnbiz/slF6AZWN6k
avi74WSFSW3uRFLicxEvOuL/3BIhaz66PasD1HqVOOLgiiMSduHiC7KNFZuEBgsoe8Q/ccyEWm/6
0uIwTrLouOwOa6YSuywWx4sHf0ggmJ0wObGxPEZL2bMu07BkgIF0GcyHgQN25JW8+AltntL9ABCk
ShzMNtJzdtqvJTj9y6SBuf30HiZev1OuZkusm4KdYoXjJGEev4r0xnZKsLb+gVDddEqDRCJfUwUV
AkeTk4KYWXSYz07/qEXtgDWcqq1Z2b7vzXmBr4ow9KDEBzA3KlLHSR9XQ3+5+BiHeBNtdPj1f9hF
l/R4tDzwlhdnv+uXHY31wW7m7qmDRRj/lA9M/jY6svl2lHp9r3FbqE43JBHrNLxlwsGMhM5/8DBQ
eB0eO67ktDtwfeSlr/hFwc0lFI19hIF5rrfl5XZc9xeUU4GY5TVeiwdeqIuW6ma95pp7OSZ1LUu3
j9GhXLRkHnZc0jBcyg9kADLpzefQfGlV/gJh0pvyxgB+gLGS0Yi1nX07tI1N0ZXPW+X5zEf6xPFV
UWtBcSn3wpjFaFl6UnEXBjqgLa03KQRLTdf5vE2JsT2skyCn5XBuyo5yeFstY3PReVexo9jGvbrp
C02W0aibC3bBrfl7/aB/s0w0wMsC7PZlZ22Bq3md+sCd2LRJm5fXnaGKRBuI15IOqZ9/0L7fLLh0
sfDzrXiuinCroEL351+J3H7gWbuXsbIQL5/JDyoAx0lrLyogNJ+Na9DHeQ61rBJfEtScLXI+lDoN
FRFUupIj+DMIPi7bi+Ghi5RmhNauospwZ2qGXyat5HqzTNODTirbNc0apNT0fjp0zMMQOuvpXXqD
DaGWycoT7qrNtoKpHQk24nYErlvKZBv6r5nOUJuN2TOiXcNeuudfjnR43nBoyZUqfBXd3ZMlR5UA
HcQneCk3yBqpnv9tTDwQS2MF0nUTAeWSLneCVg5oBdopcR02nYVp32ez+NoL/C3/o/UGhUXaDCpA
krbdUW/XXppIzLqAkrnxCDD25RkcNQ440uR4gSzG1dzbkEyrphiiGMuHBNOhktWj9SqNz4SbSsJX
e3uwgx86v5SQIYbFex55m/F5ur/ec2kJUNj7SE7o/japU+8lFFOJe6PDZkV0Pm2wzOYmWS/oD+VN
3H+5+IAMFZALj9i7oWz+Yzui2Jv4raqRafaG3GI2AzlptrHr/9hojKTx9TLF1EYTtARGYv0JoY6y
vz/kwvWe2wP6Ho/89vynjxzOSZyNUIU+EdbFOh2FyUpWKwGHlmZP8kj1DcOPxLoqzv+tEdyEmrIO
wA8BIlViCYNYAQxb3OSwLJPXVxwqZCF4cKpB+c5P+9t9FnEdfmOOwzlWBmsPY35VlHVQJn6++eeR
7TAl3attsgVniBQ7vfWxq08PdY9p/X2uEOnhwgiLoXaurfauNbcFg7QW6ILupYL9dJ2MRpRKNbnv
PDlHU3ZcuzIbIqRpiR/dWjbsvu5IO5PAnLNId2wUT47CJ6eDOUTw6v7mSrxR9q/DpaTxvGGmn6v7
dL57ZapY/liGKu904iVy7paySpd15utvWvwbyYMW9SByd+vqz8bfIZLpHfW7uKJbaGTSUOgGSFhS
Z3fJlWXcgQraZhAfDex0ZOv5nlBjaAZFJuLFR/AG6yzUaKK+AKYZqINnC0Res1NxjvgPGa6RliL3
GAmw1fAsKSoGGu3OAyxjOy0J1IQXOzcTRSWtvek5/+PuA/pSfXhLDU/fWMSNLaGH/H4AGCmlq8cF
+iTUvlijUDoTWxP3zp8oXOGPDVnBniDb1fff8x0xYci+760npgiSv7zPAGfh9WTVubaFx70xkH2s
gQiOZ54YolPLtKlpSfo02oP0ndZIZ9SBIiWXCTvJOvTARSTNQ9+rTndHOuOpH1XGLvWaVLr0acCP
bROj+yFhjvbdV80h1E/LCFeLS4apw2NvxCsREhPOUj9zXrA3qsVwf8n0kt6drUJ2cat+5mtqOozW
/idMs3hzvkmgYUxsT/XXbHH9Ida5e7GISOLK4hN2G4W1cTdu8T/PiTOqThb3w/Q3rUB7/KCX/Slz
grP4LD1geVsinAZRRUYV+mtP/qw7qQZ/ExcWCYIg1IDLGKzAzk/sl+opQeenW/e/moEIOoUl0NcH
3Pc2/ickAHTEP1QJd8Mv4IRqZkLKGDHz1JCI5YUaUTHMRwgFryPg1VO6xdS/00XHj28JF8uKjrXk
QGgWERRywYg2c22AkUEEorIsG6TdZSN9iXvOrenZTIhOrWAWqRJFPlOlgidSffRJR21e2jHJbLyx
HT3lqJjeoSlZ5xKvdi2R2lwP5lU1WDhj36yp7adIHtpIOlCu5EaC8aMRBY8Kbbr9nqswAVzDYnrh
e1LAGOh3jbjcizOD/Mdkvu37O9mWxrba6E2bHDe8T22VA5tVjsgZ/1m9ZxqVf2lp9z1jyNLsqmK8
lR32KXGCgmHlfChpSvVokDZaF3ZA1OjcJOAdRrio+HnwJTnmAAbNldP6G/kjGi6zHSPvZvzdhTk9
jx6y1OCQrzLilhL8kiGAEofg4ZF83ciTDiHAxdov3zKW8RFzgHERMbuU8RuR59dw3ontyEcwFmCE
VOfVg3CeMnpCPJm1F3EC1ypC9GYrhimijfseuu6LJL3dzfneLOyfkTEc4otH0cUp6VeHmTvLHyQz
JI2R3ASZoWvPrnrnMC1in1bCCYc3MrHcWGABFZvdp8vrsdfBamCTlrf7IIimW2DaelsvFBebhBd6
KeW2KBwqutlHnK2vVSq1i9kpaZEKQQozm8LmmMaOPOdaAvhP1MxuVg007XP+NkX9n1O53FX81VPD
y1EJprtU30uV403/s6KcCEx5f9J6ApM7ZycRemBLrt2NhaUPfW3ZzgRues+XM2oUjT2BKI6xR9kW
ezde/+I7556HI9XMS/52g4bkVS048uvfWpVdnOBLezJrr8hOXPdpvpjTEFqivjIauhSqiMa+JqRj
4difXZKNc8uGIfhYeXm+8jVjrne/YhLuNITlSPBu1cFRNYNPJOx5fAzjx/bSdiql+nOvepxpjyXW
UwvPj+RaUkgKUESMdhmWZ0HRMEu0lNSd6fbhnohSEVC1gs6ZcGOxxccxJGwULIgHH7yV9P4A+mLA
m29PyvPLI0Q7t6KZumv9CPFz+425dGvZORa3Lfq82AdjAnGSVvUk3AVsPJXoapIg3iy+RFsf8MYq
xNKAr2TjnJlHN3xcj79snI1USxEN10M5CwamLC6rZB0JxdS3VypNPb8YoXBM1cFc3RL4aniel6Ro
gxS13NJxvI+CrWmKY9QqGkGj1C1AnxhbA8ugfxYLfSBV3FkaR3yBBAWotXIDU0V16JIhgeTMEckw
pGRHIsDCWL8nBV8fpUB3bPd6Mspcjr1En3wgqiUBqnZmXTbltCyWV2cumjrxpCUvgJi2nZ0wrs4W
xbOpzyELuvXRoikQb2+yksh0M2nJMqatueTUnsQjbNbfXZgtF09LiPPNy/QWpI8IKY/IG8qNOXuf
b/bozg/arzVhpVrnKswc8nUEQDDajaSZqzhIEPm47suzSkKTYIn0Jnm+7SBSIG9CncFxetWvuUFo
ceR9OxcEExGSGUAQMuIflfLyu/E+yWHNLLdaELuB3YY0uAtlZ5Glt00joQ9V7rDOHKt7eOAW1LFY
t7H3ieAXhwnFs/KXWOs8Jc0ImeIeyhvcoWcJ7nnwicTdEej3uVnO1nSYeUWghkBsWiXKB/rdWGUY
oCWMEyTGILxsx/t5ezZu/AZovJnt5uSB3zFXhoM31OC9U3i1C75x5qi65xobYbmEbWwL5/Zhqtxa
s2YF2a+LB8w8hwpTSmuArHjbBQzYlmD5SWbgwl7dlc1f1rv9DNurFKYRuq5kV4Z78H8Z+6Rl2UEf
kZHv91FVU57s0zjD9URzTXikwcS74ZmgR1fkd+5OLtncK3ggWXzVtf6ozvBbd3xUZsK04lZNkU2O
GGIPjq00LtGw5FVD98bfqJEG/BRozNzuD2420nlqmBAL876qE6PIRIENwhqO9L9OTnNA1PVorljb
glxxepxIj/0V7gupHBinV5EUYbOAMLAcEGRtMRKtZIz6RhGaCuXTv9i1mFh4azXWy+k4mCUkCgfk
ILDcl/2lWrXS4zjYGT38rqMbVax/8F4ETeNasM2+GuJcQ001JOsmMbRntYTdmT9w2DWZumZu48vG
5PlmsIyg7T6A+K1OkCP95Zwe/x3ImC+GKd2DuHhgymyCh+D2szqEBA87l6W+fhdZ2MHmScHAbJZv
i5MUr7XomZkNy+Sj35kBm9mSC+Vn7TMix4or3IXbynDoh/Gq9s2gkRT+2vMus/6pEmX9tfterjHq
paiEYCQIdur7y6QkkwnzQy8oJoqlTXxLqym+I35Y37Dkd2ZpGtH7trKtJZ7c2VXV9J3empaykcum
ZiGatkyBUaYa8sLjWACaArlCEDgW0duMchv4s+hiVGSikSv8letplOnmG/kC3z1SPvdF0thRr4y0
D2qAm6LXIaLaN+C1jCHDPPWJ2g7q8ySe62nEEEoUbnZj6qCEnrJ69nLgs1Va/eXiGFHkLpRaDwno
uab/sOWz8qnzVzkY0z2MUl0jm5yblU9t/pfmpCsxY6g6NxT/w5l0epBr78TPr8qOBYKLris9m4CM
/1jOgLP1+xXHCm6uynhPPPm9Be2UbSd1ggPAKrgXQgSOiI0UrW6s+Z1bhG+8ffdl9SOKR/CS3XzD
9S3uhP3yepbKgVWQfnQFauJzkCbdIjHjUl4qptXM7/zgK1o1AYoBIlxEFbl0Xxe8m8teLUSgRpZA
pT6B3hIWpQJfDvTgGo5DIIieHX2QenHYqCchQ5lNyo1Bi3WuxNWTitkb6s6KNo28Cr8VP1J4CMBY
nZZaojWO0n31OuuV6GdZ1mjBoN1vXly90t8jS3SiiKQbx+7sIP331MdHUzgfr+npFXe6uYjEZCzs
EvR63YHKoE/5udFYXDRDY+boabSbyMSGcTkZITjbpngIef3klzb+Fipkwp+x74Mb8Wn3jk/o6g0h
TRlnaq53zunzUhyXJhY/YfI7hNdp8eg0jKsRKdq508D+KOdcld9XqgZ0GRnizKIok6KyeF8YEoe4
rWQJRBEWChbmaOxDAR75w2WAX51ZYJwhzVpOyrvCXyijPNLPXf7xiqC/N0BOXct+Db+kOhFqvG7N
aJcSg86z5MjVGA6f7eRUr+MNzNaCVwQ9QpluTaczByZ/fBE2lmsEuKAzm2uBR8sfCfiskbBx3DG9
EF8yWXBOeu58aOWNSZVBIJxpkPOuWwW9brKHe8UkUfsJAIGvlIa9so5S0ipPs3MA7JMAaT1iXYY/
gcKVGGnglR7oYfSJ2A5+olnqeYl4b9QtzGDltOrvhSXJxFClfA1p4yShIHNx2y8Zk8oi8pBxsB2J
kLUlzKYOQpnSsmihtlAFjRuEh0tH7pxenCDsRTpnCaEUDJBiNHniY451RorAiV63G+wFIXdftHkZ
75eznaa2QkrolQjQV3tQtdtOUbG5FrhZ+DhSrp8LAbeuTX4/9LkJZZq4Qji+Z/9/K21ko9w77mQ0
sv32/Xd7GOwbrbxxwXIK1Mn+8OTn9zPVAcx7HdGdEX108ChVtveuYoU7SBvejDWOIEKF03KDX18q
qFPO66mPCKooL0VLScc2IfnBjpTpqtDNrYdXB4s12cS8oemQQUXFbhtyMmuEbbcAjqpUAk4GYRgI
NsWQZxPuLXg5yr2S7R2A8CQsFS7B/JQG8qnbAevRbPJ0UQeKriZYMip5lgctEnMblDtHWC8GpW4p
ktipLDPj+VDrbUzTUGTIXMmYxbeKyEhOLlX0zz6Jlnvtmy4mEZIDLB1k6lHjzgZmjsi0/LLOjCOm
bnuzg05YksE/6TOscCVgGqrbHlUQvxi56IsI7gOua5HrymjTvzYXoID9jGdD6R82Bx0c5jkQy8DA
lNKjLSo5Z8QggBwcBOwOGLbFA6OIpWru5XZyWT2i8T0WbLHej9FAAwbovgIlJIZpDZz7IpmLhX36
rMdwCSbn2hPgtyQTpWltENexrL4Q0zSjdIPk2o/V0DP1eqwTn6XfaQ6PC6soaxSNzRT0wsuULBZj
lJ2XKbcmY1cR2+oBti/J1yRBlhsWN///UF2Rjr4mf1SP9bUI9xtNSdhBax7fOSZYXN90nFh8UMey
l/8BBjcK0fN6S/f4Q8K7c082H9NLD3IhurnkbZm5HhOYaCtw9U2+82XPnQRxBCzXBRBRMSjmHvOU
xW3+SpTw3C5bDyXl+7duUBFcTk/o77PyZjsclGiLxl2AFyG1q7Gw6F3nDu89aPCaKRllUW8hQ7AC
tS/b63yoQPC1/2w4y3cl79fD5yU9qTRiqbtKW9cqmIuATRBI9PaednRW4RXO0VycTd8mwyfDl6XQ
pkw+HvrTSe4AVn5dwt8c/aU9+PgeNYLvaI59/AuAx6D59d7ekAFF5HvJeAwTBU7G/equB37wGcjS
1t9AUPRkIYAX7xgD/bzAXGAuW64/yqlk52TbkOImGIbizHafFrCb6GkHarPPh6GOJa6hflkxUZ99
gv1DOv90evfepg7qxRn6Ci1CytWthb+X6ZbkVcuuJ3sTBZQo14ALDmGODgOdW1Z0CB1CPborXtuT
Me85xTeg/2fLUg4lnNCaX6omnkIk++rKcZh/MnaAyJ8bfsCfS4db7G0kuWtH5Ixv7Mk+yMO/htKY
RL+dra9MSLAX8y7T3hnkkdp61QrzRvrMXJTvg6WDJlg6sWYZSFRjmFb6n9mDhdpM7Y5xMTLVFCY8
zwoBUGrdPCMllr595HdPvwORFbGfDF9c3ZqOVe1+5O7pwiSriDLyPHJ2HP3bBhWqBPZi9/Z17hRl
YagiYRBpDGySAss0zGpQb/G4+AMEWPaNKOVV+i3yxA2BOouDZABxpoW9DjTzy92Xld5nuurfgaIv
d09nYn9gQkAVEQXBSInAP++CF56GQTNws9Ki3Ey6AEsiNr0izF5qx9CwgAa+SLR5ZjYIshyZ+LsV
lICcUn39EEOdropHb5S8V5NMCThARzxnU1V4reXRCHMSUeqjPtRPf8/YD6VMjaQcYmpo/CGeSU6s
d8AeGioFC6fLNCVnWPnM9tFcLxjc2+iOzjjEkJbxAXTpoS1lWKes7MyVyvTnHxkLXF9891Svfnil
gWTX9x6AfuWRdVAfz0qeIGUcaxppA2FClz3Vq4x4EfMX2ACzwoWyZPKRTJ3rq8n9z3ag8g9gLrom
un10wpTqDDLn7c/gWfyTQuE9ux3VOs9Jo4CJOHxkd+a8bypoA36xLsFSz5pCVBV3s6uOX/kj+nR1
3cIOdx/fp0Sm2TsZtu5JhgKvdFzyDiTJpGndE4MhVOniGPiF1pYv+eGDuJePPuPuUKECvodis6Ek
IQUsYqkU92cinEzcl97kHK7l1AwfiaYIuv6L+RYzZg5klX66vKHi5WYUEDMOWU8P9HfkREQUa6Hf
ym9HMy0x232SYnWpWTQ7u0nQUe50cdueKAxkJHGlKgyhgLnPv1U3MLyXvxVRmV1sFvNh8HgpQ9kz
0Bk90cjPcIK1Wl/UxsWctbzO0VYphQZU+i8J3KqhkEXiMaiNTAkWK7GKXBjL+A3YzZBfvgJPkFVO
D/D4lE0brRPn6ZLTdGKj1WRwJugvxTYu501+WjYS+SiyY30obUXjN1EXqftI/FTUFy+FOKuZRtKM
xz1jpg8YSGM/mS8n1xGmZPTz33aMnwNy6VX4INfbD0hHRvCBkkpH6L3c7+9E7EqX5f4Dh84/Xecs
tU+nnvIL8sCAdQRkckIcsvbjzki5VsjREcJv9EL9om/V42hRK5bPR6jXyCZdFanyuplaLbltEXmZ
LcrpKqtld2O8HZSU1xk4IlOThFrG2S514THh811XfDsby/uRFpv63agLOBC2A0kKRR0iKclTI81n
aoHKwkyxypwqgWrP/LLrHYTLRVjfe9LuX7as7XfN+Oor7R7pq1XB8sS1IOKt941gRrn0xm/JLjgm
1RQUEYzGxXzHmcSXixPPGIXSkvifF08UzpdmzAtzAG1McZQbwhxl8yKjwPPfSOPTMvIeH5p8q1jt
i/Zu5SGDDshVdbNcDQoetsAbGEblykEH7y+fxyPkVTHfOOCw5syB7qJIDOdXmRQGyFoAnSKyFo+z
quEVM295jMnIH4NRZBvrezceQlhDnC9pHVRvT8HpyhdOqpPan1c84Wq6f14ioP2K9pGlwZh+HajP
kjH7TB1gPibTN7cuKnuEUbgbGn9UFwV/GFHXvOFsa/UHGJ0DGr6txWbLpvp5y6OQetElSKakhSZg
EC7MMfWfpP7d+/FipAGw2GNbDfPjYsmhKALcjmQWsXWLZoac6oM5sj2Z8YoJ6e9CjMLpjjoVbzhW
iGrUnnPkx0TSPBiYpengynSPlaxWdIZSBEL7MmZLKQO2c9zgr4z7K/Y1m/zn5qn8WnTkE/fDbrm0
PeF9kEYX5pUqn0Aur4Er8CpKGJWs1R3dYt8N7wz/oGrwZ3nMOk93GKrRG3ifxnZml+NBUs9rjjyU
PHe2JU/pGZXGvFfJmupe0jDUimKhKfjexXwCaJSuCY1OLaR10SovBbv5Pl9kC9Yk7XF2LhcAqfPg
ppWO4tKZaXXPiQHsEGyAb2F6mXrKSmurPcInfZaTUh4uFeUTFCQwKdtQRhBqVybb7tYi2h3rBIN0
rrlJVPjuCttmKF+ekEe6anT8WND08h3YN08pXGQfWWOi7Km7h/VoG3ROAMlyNgxZDLuLMdAb38TD
DR53RBa1+VYxwS7OdlnjrSQshyjhE1NcgijukutQ0/7nUqBYJTJM7kNk6yrNiN5uHiPVR31PNXro
Ug/Og0N92zrMjvx0udYK1n6NhbrzFdM32DKKaE93zlpSM+e36MyAoDk2cuxtC/51Oui3U3DG/jDL
pxaOaUSb5+SJ5VHTa0JTXj8xx9mEZJw38A9i5gRXlVYjML/UFmWuL6AWXfTG73odb3GPEo7L/jtu
oGnHk2kFC26tKk9w1p8ZR1FvefBrO5YbGgZTvLUv2dFsUMLMCjRdvVGLe5LzTXrPevOSXIuLxR0s
4Vfq6F+2NQxiy7QYMXmgrENID1oBRTrFjjCBuYsC/80aHtjULabVzsIVb5QIuL2zFYteWW89x2wZ
EM8kRYngZrcly4aTOVv7H7BQE062HePJVy3ubSRAEvLZkExvAQGOeYnHdXUX/Kfz2gLm2ohZ5GBN
DYTGev2ZYUmU2vknJd4TWZRGLI0EB2Q66XsnfOUlhj3bbvjWJuE81nHdMbwQ932yQcSMzFJ+UGf3
aZ+U/dAnksrX4n+iXGYTwDYCtPHDLQ4BIx/0qyHu6bzVyDqhv44D1oPIQKGpLScZkS60Q3MoTgFz
7TEj3aES0kuP1Hl+yMh520X4/xbrCa5KqeUFSBN8yCggR4MD219YuOTjC5pnFI/Yp8Lr9OKXY0qD
kKhI4hzI2v4CbeDvUPIBmptdPXeuUdF2ACrfrOC6OC+MrjufIkmgOAhBOpDke9CwHUljB1JtcL2G
PVfHyz8CdhNsktKvBdDvYwLNVHoFhar/EvibVbupcWElcUMBSXhSThuxbOwA+zavZ+aE6P45WpdD
Hawo5aKPckMUxq7X0jifE/pSr7SPuMDyQDnnbKlZQW+WHVUa3jS/XSObxj7BFNL+pXXIcXbZ08jz
tpHqw4LblV7+YnenYCBZrZZHHwRXeLcDGlP3dkD+i547qrqMKYl3yg/Xr/4cX36bPCKrteC9mczM
+/49ILDMhenmiSUQi76C1S+TCOzuTNYqLu+lCZmRWjFL+Wtp6J9dejHMWLPLPlXNlKkIzdi34uU0
rXSNQRt6gFD+GpvwFhEUtYrATtoHcizXtb7hPg9r+g3qyK1DiuADA34WncB6RWWQyOZaZsNfYP7J
BOBIOZnD8tkUL3mNRHL2VB5eVlKD5MC2bSpaZCrMHfIteybe5jiVai2/M/aUnN2TbaOvqcutpHXV
XWVXv3Aaj7ZT6uxwA0mkeg1DnRU5EjfBh/I4d4iBwGfkPL9ADfyOAqT15OYPrMDgtDseUI14kysx
tvq/Cl0AeEd2ZvjdKZqLFQwX4b+AUmfZ/iNaZT+pSeqg+eROvFZVrZA9ZNMgfffzf50tXLyMSzQr
/c9i7ph5VhN5NUD8o6RR4lrqr0207FMjB5qKzDyrT9ir1izUtPPJFOFgIgvzDAZ83J2cTOWZlxci
1XZmyfP/rT2twChXycfR3JulBnJt5IfSsdyuE6DbZdWiXXHbuLxoLrZr5daZxepD732CH9YtN6Yk
f+O6948ZIDJCnMxKlrA5+GNM+TsqNUQkF/ruIYsRsCzTJKcEWhg8rXyDPPqBmhPUXg2AYpiQdtOS
dCI9Wlj9UopLllCD2op29qIkOf5VtFpTD2CwQjNIkECrLUxw2ZKPjlFPhByqHFR4lERIi/F6R6C4
Gn9Cj68I2YqZ6MgcMFZcUxisen7NH6Sz5bXpfMgYug/TE9AocZ3UCPjH9NyD2uIvIaYhHlokWgj0
tjGHlJprnozcTJdbmQ37tpOsB4z59VQlQ9fHJF5j5s9CFk4b7HaOz5SpWBX4tK+5eu3yjrssTNIt
avOf7ibXEBK2uz74pUiBs057WKzg4gBQyOPOl8wl71Pqpv3of/HOdEixxCpcd7dXi4ZKyaFrgH99
idLnQ6/a6M28KGsSPfrqvi0gWfZ3wyqqEunWNgQCQnY2tqn5i/Nw/rIdQoHRsaExW3Z/7ox9AkFr
XYg6fcjoSRYtZYOpPZL0aypGYOKagBnWG54+AQ54lIyjEeYZJrrDAoPw5HuNJsfk1nhHBlPISs8U
7CO2Znh107EjZKzKwSOwOKU0FkzPQpmqBH9mp4hP37224VLvoWXT44jM6eFmmypvfKdIV63S7BLC
sB4QHy1X+SGW90OiSGoP8AlIYR0rg8xTmykybkQGtnY7xKADqoedymcJqvc6Esd1lOe7C/mD/I2d
1AFHR0+LLw93x/LrpqsAXBpVczP/6O2Y4IaLvD5rB7IquY7j4EkbWuJZt4nj1Wlffsi0KPP1CWLE
/TrCsHa0dw+LkgNW/3xOdntu1tm7F5vq1WYueKrqrGtdXCv1xFqUl3jGW4xFq+vnRvMjQ08oNSog
bQSfJG2E3yV/0XPOlhksVhNKog++GPH94IOfwO3a4yRW/GwpS7MwtU+7JM8KWvan5/hFUltpuJyQ
szp/8Cn3WPieyyaymij2pHj7nXtiFreyh6osANavPqsACsJf46sw/y3Fps1F53NKtkN4yl5i15Kw
xLIU45DycRjYHZwZlMM6aOhBLbvjCDWt+5BQRN7674zlEnEBBUW/4HiBlXsm5BErYOeNx509nfx4
Tje/GxaI6kcnN4o+4Ul3+6s7BNrBE1jRsB2hH6HYuW9NeUQdq+pQmFsZAa307/tUhOrYhLSM4tc1
0p3kq82Hysk7X3DNJM5qEaRyU2cvc0776tzgDoTvAtAwGZgzMRZ8m+4WnkzyuPdySdK6VOrivHRq
GzwrTz4JRThc/FMZyCxJF2tKS7SimFVwxcW4wZl2EJzcD7Md5KjjMM0UPErhCYN621Jv0HMsLTkY
/yhf+RWr3hlQVHDA6wsxLr9izX6rg0QJx3LViK0PkUPYI2G9hgnc8Z2IvhTxZLXchShuCx/nheu3
W8Y7vA+nVshf7oe3WPnAUhxXxgaS0WCkshmEtyWb6Z+y8bifktTN+K8meEo2rT+49EFRwJUkRkUX
07X0gnZa/DkV5rejJgl0HSw1mbYXJggqT4rc70la247vlKXKgzEI//fnzArWSc0gwZr0uYUO3jOy
g8PI62shFMbLfJXw98jVAC7ZL7dkAP79wojCFyUpDHcmk6KodUG9XgV4bmPePuVf0NM3DfRgiiO+
CyUp71GuuHgJcrv87nTvRLix0HQZhVALQ0gzW6Fcd8xeedUW9v2oq3tVEdG7ph8l+kcqZdjkW0da
JwcCFrZB2HH6Is/D5kcbGvaCThArD40gNmCmkRVPl5wJ64WDNiewiD1KzEcCz8wUzyfpj+s8v/DA
MXlrkIJNMPVa8MrIn79A1Aflai9O7IUT9gcCY3PgLp1Y06v3vvWPhUlNxGeKhRzys6rqDHyEQ0Hl
VxqH//r0gfkhm1QjCF0QtMeO+eM7HiF1lkNz2nipCGW3YEtXap0ngtieVl0ktnE5NuLL0lSYgqj8
wqUz5mpEDJKqvXLGrRAoj5NF6kHF2XXLq5+FGZAwaytPq7Aaib18owi62KcPJH6HdmhTNk5e4vZO
UEtleEMKhgQrCArNiQr7Z5JD0RcYDXs+Rd6psyilCDx3XjoJSLUgOHmDMG/zF/w9owkUCcnfSDoS
l5PON1jkeg7RFUKQN0VooS6S39gfl129tru49P6dzvozOyI9s44HfNOzcg3mLRK7JWf5Yqb+VKgl
v33EdQp+jF0QsEMt8sSFJzySFJ+q+XbW5IHqhykAuuAp65heB+Wy4wOBhKpd7k0W1hMqVF9A9DR3
YSep7QqSj8l/ftvSgE14jscvaPy3yL9LvIv39wsgTPO+3CPM/43rvCO18ofXxj/Qf68nvp3gXFvy
jIvzKBmcg2zdpI3IFAVA2H1IThoWVilRqWBdCFw0lJDmKDAecFsn+uJZGYPB1JyJw0jZ3FhekmHU
CZNTHAqnx98RROrP/ZoGKUGOrWIHk+EzZkQqsFQQdG2yIMAoHsF3V3Ee94bZgwyBFxRCME4timsE
gbNSlJds/p2gGzdtpaSQ0ePi7CMBtQqsCJobTX0jPjXpz4NfMJg//fsn4DWNOSWoaY4WRL7YPSHv
65v821ZLEk6AQxTNk8Iyout9AtZmBMysPJ+36lSkhGkT+jNiIclE5lc5rGdUZUgb1mRk4aMlpcS+
SX8pqPbguS1V+XHZpPWFXQQPYehq2a1I8LUbxZrbv4dfClFii+/17rQVJ+57G35URESuyfacSJ0N
la0NrjKhHM1r4JomcNYqN5Xr6sdvpmdyeROe0wxDzBW25I8j+hjtFQiHQAaVQgNEmcYgl6YdGPjU
Mpo8Bq2MKOjqVJDyyWEXZhxjuZyEYonPwp5oavQeB2Ozscd9d/o1od3QYhDxL33Zcmj7wcHOmEhM
hAf+SzevLPT4vxoS1iC0s5SzDqeCmCNxyo0xVEM71q9RsKMnV1F+qKd5TTSZP5umvBgO73quRRpY
HOQHjPL5mns/5c+li23IUcdyBsISFEJQsabcbRRHY1IY9T+d6IfG3oLHfqUlSZVgwIfJ2QtFGRyt
oQylZ+7WneHc584TyoFz8bR3lXofJS5QMMOa575W+absQMuEsZzEW6dDDEaKAdFya8WFiahtpUvC
Q0t6zYG3AmFK1vWiiBKVHv5M8/ebaJIk4WdFFLrsfFHMSzGjtdxmiCoEK7vXR5J+S3YXuCEDLh7t
0mRd/t7UjtAhgbRCZorjC136W8iVeFW8baSJLcWySp3Zr/IY1R7USXXVPnFcXiZbXLj5m9bYPXVd
0jUfo9s0959NeWycJe++1nTrMpeyXbpZDHURgXs6bLBPEmwqvp/g1PbblBDFc0xKFnMJQfrjvo1i
XNhnPPkkZf6O2H4TOVyv8bujqQtsjABCJOlVf/jctFX4bGsRpXW0Xy1gC/JZvX/fAytnLlJRhcb4
Zb/2zu7ZFSHHgqgU+1PUyXJSVw5FTZSucWwsiFRsrkq9OqNCL2JbU0VhORDdbedSfYEwhFH61zpG
aS2m6xllaR1x0XtymaFweMdygkehdaX2CGbKST1+6EdxJTW3/LmDnY5ZhtCFZ2K9FnhKX7yzfNmY
JDeNg6oGxb807CKU6ukdi3tVrNyAJpfO0Xx1u52yu64edLSzR0VEJJ1m1seILcySMSmmu8TDDZPe
sv3x8Z+6e7NdoRXLwiEk96ZTn0LAtDF36ItKJqV2UlZ2D/tv5AbmM0VFvNlzhtadpZFQLWvX04cI
jQeGfGPsGpXPbALeez5FznpW7IUFR+kJCUhHLBgVENx+7nP1HCDGfvUtVYotNt849eQ7KWnXbVHE
dbBzYbnzb8CsdbmiDEdZvYl7V/cVbQYtjQGIYgik2qC9atVa/39PjOpb3uB1M+VvOsNnv5DFsVBk
lwmCE2Fe2LtizuWxKv7s9x4uh/67xFmrddl4XBXZLNBCcccQSR0gPHM8FjXbu5wrqszZ13Lb11bj
12bJoefak4YK9OQNwLB0cW8NM6m1bCobw/gYK+FUNRutTkGXzxFpidpFG5GfWLboESCt0pPxHe6D
W0t6gWkBCPNhmLd3dSF6gJeRPgfgT8ULh9tDVpqrQD9z6xwfpXzFtqXem8cFZkZsLiWMfFhfcZX4
WXR6vQ3dOQmM52Mvrh96llAhUSfZ6nKyj/qoLdzdCM1+FW7Vk+j6uOOqRn1JRrHULT4dMpe8RQ6x
zz0IfMTBPOgMdCs09OF0SvX5JoGDOnaTgtFyTYX91gaampmiIoXzYwJyHN3yvMyQmq5BhIhxbeNU
UGKnxU8YxIcIu9/g1A7jjToZxpqXkyuS7wEUEtWCWAJg2bqJzxyxKOr49bD2Vh/TOx7pbsU5Zcvf
P8I2dxAurOszzZtlwj31e4WiHVAUCZKPVqpy/zgJtVBY5s6ocwc19zjWbNt/HanTly/+CxpS7/Dl
w60SRzqHVwyQy3D+LwlSAfKtIg8mHBMA+SfShYmN2kkprQPnl+4qVZLKRNCuEpQ44uCWOHKCgPpt
nXEBDzfNxzASodN7grbivJIQoqeY2N7nHKzzEJxvT0jnB/NaempmIkXCf+MargkM4uNgw9F0m0C+
Ad9Ap3x6+wZmfDHC6p3+E2SOGqYg3qI867KwoQ76vTOPh9E4FfVYDHZRz0b34yV3peGana9SAhv8
lWbEh9pyDaGm1s4vVsuXpEjxq1LDnQ3B2atHK22y7XfGCLVx7KOyKFY8QReitD6KEu9B0lZls0bh
VJRVQh+tf6iLAiwGq9fr6+EcZWxvjBb13Di7ycjtCAlF8WP6BXhhPZ1D9kuuqyYssEPMUxLShKf+
w3jEd92s1jqoX6hhWZOdDZo9vH3aZ4KGn9YAUIUDrSnP0wkXBxj0UabrF/xNH4Yx6/6w1KBC52az
huVno/VkfhBWTjqPVfCu5x/7AH667cetsosoOqSCloFrH9dbLDaQSCZUZloFephXJQcG/wV6vNiE
10XbRGz61y8hdgb7QGkboK1id169HVVC7UgIv62HXigG0Spt+FEVx+9Q+Ipnw7p7YBLfiKuaRpLe
76P2ttG4/l6j+i+G2fPaaH+wh85vn3TCAKI7LfL0ChUmpRniPiZdwF3TE4Dn8XyCE6OZzQkmL6wW
MDfxqIs+0MloYdAZZYTDfxUNnfo6PfJslSKYV+fJO88uM0D8VYrlaDsRm3sA4DBf3yoTVDTiXeKK
DOnGOekz094JW7OMOks3giiBcXVheMSFmUmw7bg2wtFbLipKrC1CTI8vdl24kol+oH5Xjkp5Szww
jXDl7ehk6u4QD+aLvCVS09ZKPDXMu59OQWH3kOcPJwnjlH8PJqG5/sxGb8TTErnh70DAZ24k7iSd
pDHciBGpJMfryL2TxVtYlHifBmr0m2B7gJ/IF3EfGuDk4Ie5jPFjloL4CJDd1ae2qMvq9gmgkbOg
yQNlQZ+o4dahlMs3zPSlyo2YbghIa7hibCRRUUEZVQJwENi6j7PX2X6oxcyli2ftvqofniyvmS7T
7BqAFyBmCVaBPxItUyGKCNtSHJEMSdoIMPZ+d9N7DDgE1wz64BIyD6abuqjPZdCh/sU2aSzX+1O0
uNk/P/XfP1Hw0+f0LZCFgBl2j5+zTefX58EFvUgYftvL0q8lTmIhSKAjhV44xjwoDz56yJx0KIXT
4DyF6CRfLzDX19WUUECf7bTNPQbn4tI5++PDvqgybrnlyWuyuEOCtvEBz4JVjtvbaMZqdHPCEfMz
jQ+Nw+Svpshhp2z69Yj33byktQkaUMW69JrZHb2IA+8+YfXrBOBVLa0IQ+kREXAB81AJK2Ux66II
dELh5nB8/SQYxvNChRI63Ui2X1gwewihsOsE+duB1trP39xdcolEao1jzAPz9wkg9BBwbjBiEkV6
DtmnIm0tW+Uk9XzEIVH8hxTOai4iPa3ku3EtqKjspt8EcmBex0im+35LbkSZvNJvfYhJg/Wntpbb
gH0Q3JyApAUOyfrG+RgkzWxHfeMAPaaXM8/46aWTXrNJ4ti2IFHeOxxjOhvVZZtD7vyHh94MhK8C
try6CnG8niyFZ/wLTiG9wSPxU9ViGLQcsTNe+xayTnA3B/qNn6ITZuJp/0pKZm5xCASE9jDWyoEN
nizIqW1ZPUSq9Kb3U8RDGxRb2vjzG0aWcxGjGB6/3NAMHy2toPWZEO/aVrr+fGQ6al6Cx8ZWiJqx
5PTgbe+7nsexAqkWpdTLlF5G2tl+cm+liO3Khh3q2YX2vITq4JTyxRoh2tC6X2odjh/VUkkl5isr
HuQ1rypYqb/HWx7qgfP4eYoVN0NB9GuHySKhSF5qFBxZ7PAXVWaglM8z4KJdqz2jIx336aox7YKr
BvKJg3x4iZIEoHh5gFOB1q6YDZtwEeaiHSC5TnsjqKPkx7NLaEYh5NdlU6RKILnO25ZmcGii69bZ
EOKGktml0eyYMaKfMEt56NPYQn7SXNCbHFcXZmfDonZLeHphDCCkg4SDxV9STUzIp/PugcxCswEn
Ot8y02Uato6VGWlKMG72LOyxSNsTjrskx/eS4dcs6bxMPGC3P2BzSBs7j6k6eklxhVLbpt8is4Ve
3DajOd8CzmxUdrM0Ai8T5uLDFk9471GnhAoux7kVwlwrpl3muE86rU2yMOnIujMvkUBn34fL2Y/O
vqkm/VnsopGqOAcT19uFheApjIJN01Puv8JWSlwP0pbtSb6d+aYdQDt+i+l+JGYA2syXR1MPVx8B
pL8HLoCAmK1A7/UewzoBUKZGFnJ/SDXYqCPD0BqK8fkEckJ25UY9HAPiCataUiG8sHZ73eI0CQhl
DlQRdJ77OL6oYqQbVkBNcGB6SLzUU7YKa8YpuJMyJLT56EyHbnxiGCrKIkbOeOkTDcC9Lb1FJA97
Tdzg9mdvec2p1mDSfFlVd3dEvtYod9nPWYoYG1f2KcMDSwVrprgH6EpEjOLyPN6F9O8CmqRw1cEQ
2l0L0JrEjOgx8iAii1UjRXOWciEGr+uO18qgrfm43QchKGeBYTdBAcjoTJsGAbM12NfYYAfZPbiL
MUQVE0Gm/eexGkK5UKqrXbXak/rufmHb3ZtHditZ89kF9QX49mZ0ikm48CsJkblXGBhg8Llk/oPw
g2OoEuCz/xVRxK8VO7cAL1X5mG1KQnqAVdmVWPMjfKUXy9uRJXNp5Wp9DXM5UwG+ikwNQ0Zjgjyy
ONrgCdwI04R3Hvf/G3Lm4yhvzxfWrSml9FKgiDcc0ATyxTX63sNtnMMjeN5rFJpsXy0bPcVennYA
HAlAh0zrlhYljahhBgZgACcA7evMjwcZfaX9TESI8E9oHpYfnA1vbtYoLGVeOp1/MD2qKG5EZTt0
lIxhH7oAe/zzvCsGpPYuDeIy79EKFEGUhY3yRwoOQgrjqohhqimevDqfVKb4nV3IYSYNUmuRXaTR
rrawibdW8ncLx9Jv1iSKK4VLNB2F7KIbX61aJFuDZkeAOOgKCGhk5/TgqmTBVcAmt654bPst7PZr
TFrGgRdHZ/mtaOTxDR7LvbRlMWsWGyp9oEfnLPveZBivu4UfRq2w3ul4qi+k5oD4O78YGrTT2Rsv
YNorPX2ME4c79X+l/UJs4joPmxdMl7tLxpeVEC4H6jxU6p23OKTwg4dtqhJZqPyWQXtgh32goz2I
i6hIashdJbu7OOY2z/fJ90M6+5xPGTveAFiEjSfp/Dg7xE0oKot8Yh8qzarUFiGyYJzgVyFynCtt
5MFTfjlga9M6vt6zEK4B2oD7dB3ySTbniTIO1uzYT+9lWIezQf+VIrFXeiIZD1h7ThMgwnDMU24u
xhaTT7zUKj9YWezzrO6BCi+Ym/ypdzVRi18c2hEVErP9lo2PLdldJy8m9smH19d6MfT/ENAhDrUS
f03qj+W0m6uqviCWcvj+vfntdDC43Cu4OQqUCgK9Pb3uaZ6ewgIv/6XJgL4DdIftv7+h+ZLfoEmK
p0Xwob5s9ElKVeSkSbxkzwY1J1yL/+VFTVqm8qm6VfeRD001Cp8BKuIen/nk3hLu20VM+TYllHfM
BfCm+ySuwr/zBhAv5/wCHZs8vMovlu34LyxOrg4Cu+Inqt70PoUKOOZ2bhfKU0fR9als0tVHinDp
aaQTDJHDaNoWwMC+AutVHdB+lcyO6FDde2kgql35YEkfw7sfv5Va8sKJfuAMd2qcjX93K2OlUBtX
a00sr886I045YI/eGtNkgflQ8Vgl4L01ajQ9Q4DiOJ9yALh+KITRHjejura7KcVrjEtnVdkxX4ya
GjYVgjoTmKCdwhyJSi7Qo20jn4oiSaxIEuvE8byBuqavv7P4sqvRv1IvqtTq77/Ntnz16Mz7MO5p
huVtvQG2ZvbAkYwtoSvQ0xnGOoJrEmS3oZ9gNYtPc4Xg21OdqV7sqfx9AztKB/+atRGoDToWJRs1
9CnOA2NYlORz6lWTj1tICSJvSBKebLMP6hoyzuo5x/b6pOokorLu1/HAhFIi0vv6px6I7gkqWRgv
vHwaTXAU8O+CCyEHCYxms+sjl6Yp3ouBuvcUDP0pcrcGcjlnZobb6nVFww8mvMT0qEIlstM1Vkgk
aEqOBlvSet1YAEnR4ixee484v1H85EHBRrtBJrFdNAKSspqAlSVQLoTMFblrw9oQKEuFK6nAeHgy
ujsg9MUz6V9j8Pu24CgEbQFZEnaguqyJxUgNhzEFU+Qos0d+cDq9YiFbpAg+76Qt6UBrR0DAlEK9
TH/ImiFbO6JzKtY9Vuy+MJn6mUeZchgM1viWWZ303L/MKYWe4j6zFO9Jwik2bjMFHs3FgdpT3axD
lVztYSkiwCTzfj6ylcGx4meAV9qNvHYH9PA1shvthDv8ojq+u0jhD1QmGtQCev0on+ZUspJonT95
+v5zGg7aU1V8acS+yFL8c9UH9ybKeFOlDzUH8MlKNHeQplhbP0/e1zOMskO8bgVvdlPPsZ+xI6Xq
hKephJjx6dg+E+5kIeFZbnQ6sECIxaY+0ACZ1GTpUdbviDCBc+bHgUtus+aymljIvS9HUhTqsvJ1
Yqsm+GT0cpLo+zb2rMHMadZ0rKqxfiN44E9RjWxOMYZpBD5Xp1iropyMwTdxvRX3KlEDLfLNF2pR
T1hTjTc8Yztz+7tzX0DTYWiepoPQPg95paPTf74768XMFgLdsLWs+4mCn245qtWOn38d5nJziGQG
iekiGvnAKdo+cmDvqxqdTCxaIQUqJibVFA4iBzzVoIhvFRciAWKOPe/fGhtIonyqZ/PKsE1+4H18
SIbiFk9Ocm7xon5n/8NWWCA6S1mONpl0cXd650CoFhj55pbSHI+OgHsiAKPM4N4n8KuqOQ8P7j9v
RaWLhPNrOUs5BjdWGmVsWWWANwhhDEgzdxAnTVW7aa2JBIgjMRDn8QcNl41zHtAi9k8t6aGMVu+0
nmf4dpAQ2QhV1Ira+lG1HtuCc7AJiobC4YOHeE8sRQxNItfRBk0r2UVlbxIxzB6xaMypDE4UHGx1
QB2I52cDf6WPJD1NRwCIS840ouVEjikQ4Q9HiEic6Z9i/kn6lKIfd3h+CUucz18dAQeCMiBZqSXY
PrtGxdYwvhMqDLMeBI3N4OtfTIv43I80dQei+gpqy8UmJ8GkZ9AUGxvPdafNamWzfEWYBh6FQco1
X1TCWSOKK7mMS8nGKZuMcSTagyQDyolYdu9OKxkPWmMqNFy75w5iPZofNee+UGgnPqIa50eUTx/R
6RkaSaiOLEMvLD0UgTd6iZu4MEiDNCa9XcYfsXLYJaIjZomEBqOpB3WFdlGNYdrY/G1Npf2bofLN
+sY23Ue8IHKAlDJ/gPJmceyvQ9f+ZGbFX/vj8R15JU4asks5nXmCOOo934x9iOx1vyKqTAcjcXqB
gciu9PG+X1+zpc4bPzIx+zmwZ7PEeEWP6WwjEQnUqJ9NAf4fy8wxwzlYhGDG78dj4xz/7wyChTOP
hYOmvbhU7eYDnddKbIk8TcgP4IiZ+Sg1nV97SD3KsN+tMDt9eEyOA/Uk3CmOAqBGgIKPcig2iMMy
wyYZoWM9tlMcLRO57pvNp8me19JweMFiMXrrzkzNZnU5HVcYOY2jkt92Csu72cDyRDXt8Rq4oQD1
6ufOZ5XiJrJz92DXdJqhA8ILc9pUALo0XUbehC9CC/7vBfPYtPTN7/9hSuBEdEtl6/szA0IOoMJM
zROFhtfH606CLyWVLhVZqv/0JnsMdKVDlvG7fD9ID6brL8H7SIOCvFSoXWh6CN3JAyPkt3iftW0T
tcGHqtaBQhG+El7KR31BeeXLd4uQrqv0D88TdnVMvUFACk56vdLtfWC/Zet2kluPyIO7u/iHae8t
oyIqnamOxkfDh8fSQX7b4vQYCx9QIyVROYeSL91Cjlo0uBKVra8FlLKK1zMWzRQWM7TFtrzRaNNH
U3dgpFSbBmCn49X+6uiJyDrIwCb2Eco/SJNGyXMc7fGYE9lcFK2DZnInKm6+RpEiLvxPJeXdwrtd
8agvnAgzM+E1k0+LcCNO/yPB/Me8bkcxVP6VyRK0kXNiD5zCI8C50URvlhZXM7n14LOa+gadfpIA
Y5V4OyS4RxdXT+FgAWsSxWOgunyO6uMhR8+L8qgG9Bl94Es3IV7Q5X9V5bpqUnDaqdAEheDHXBa3
cVwErh31gH6u3W1xvoCaujPlBftX+fEBUv+b92BeZkMWUz8Xslor4EJ81qDt3rFYWEkrv5evQI8o
Z4w69Lbpx5rkvgrQwMXM2DPtzYqTLVfrDrP02ERBm87b+q+TwPGOhyjB4dY8Zsem/iEQIVJ75CEY
ua9Szm/yL7Uge4Pw8tyP06NuA5daXgje1PtG1Rwk/2gfNBl2g4xQo+bF5eO4IigtSgdighZbYSsQ
tIMAUzw+99sAqwMKCSyRCHPfFygId88hn+g/RQqzmMKkdQ0gecqw+rxVXVhwvMCdzrFTnkkSy8hx
yfZwe2TcA29eIe/dwPJyUtt0WCtSsM2t5nTTmr128FE8HwcHD9pWVekKZtHLzBlsS8edFkCT1Xuk
tEMZ2LvksV3wnbpLFyZahYecvdDoVoVw8+IDPQXFEwlaxM2Eq6IZBHXOaas+ye2qhy2oixJ44R+D
66RACsL83Xj1eLCbaJBXNAHzqA49GCkRAUzJVJaW8/cIn8inZWnqWKiRicqjdWOficQVsfstVDw0
1usZDJBl6Za1mDPCmYS48z6rme72EWCxQaiuYZV/kPQEnjkj1wj4OUOgezILqrUMzZCLt1Xj+s8F
j/yBG6QIqRi+3gFcdjuiqCCpgugR6W7sFp4NJjYg2KfGPqF/Ee1/2jhJaKApHquHQMn+ivEWCSyT
YLaS0uR52b4JA0l1lQzLCMbb3VO9yEh2GWtHVBw4VQtIAU805OVQ98qGkh2FWYef6Sx9H1c2Fe1u
SwyDJY+N6+b05CIosDCSInMgvw8b5KBy+9kml/wEvvE47gAjyskAKunObQ318c2TcwinpVWVZmee
f7nQPEJGFrVskkPir8CmsMatX9E6lc9vcpqDi8Pm2CHUplQSeRLX76BZO8PIbQRqs9yJPuQLWgYI
BkUf2GSjRxubfylwLyuKdQm1K67RUm5UcJrdVTDycr2V+kn3MqbLwVWcBnpzH4C3XYBhFGo9ud05
hYODo9ecCbHGCUZBy/ebm9BODPfo4IRFb9gJ61amGFmVyHL0VFwmTW6a5TNqTEX9WZAbu9MBeoSW
8MJcAAfwUCHxTSQzgPHdRU0hzjztQbcmHh903DbuY1Z1r16S0fFKnbOKcgp6Hq0TNY491TlZ/QXK
ZyLkHV9D0AVTFn/F0h0HmjKDi/6Ep9+AHkL0nOOprMxzvzy0XhWBnB3CISdXkTCkSSr4ofudAEiV
QTd43Z2HwcjVNjS6+rTULWYRjjXQKTFmpVULFJudQPHPzi4mCFQeSTpO8DNCFa+OjzKphPdW6qzn
FvdBB9kd0JCmXOiFibRNMs8onoyhrupTmCTbMOZK/B0Ki8+rrOlXFEMp1OS4LnEc0Hmd6WvMNHfT
x6SOX2AfES95R4ErApk//kElZnF54qHc8S3zPuzQHhqFORkbrDEt0mqK/T/HPP5W7VyOo1h6/kGC
WIjxnx9ohSrtbz0jtqBOm9d+mkv1IoI57EgiWJXxWtYDSWeLBGUDlvNowVc2TyyB8OziHiXrDk83
QJk4OhdFh9+7IAaBvLFTwQ3JI55B8s/+mSVFA7wrcB4Dbs0KG8ylocpVp0JsEjbJme9j1gIzpjZ0
Sv3PQFiLpc7HlHM1dUxdT6Lm/1HfKCQwD5C4+/UKFym8igxXQ/tpk833RRwpcWZSDqG4Agcdfqqu
AJ6/DjDfVBjeWC40Ekfe5GMQvR0hxftUJnRlAZxG4iXuWFVofMJeKK8z1VvwvPZ1MTR7NbR6xMb9
ipoFn6T4mDkASIXZirQgI3z8EnDlOmb0N6TONqgcja44UH60AXcUMWP3CwKffz3G8D8rMQmJ2OfA
3weFzHr95eDnGQezAx9sSPRkf5VXbAKENjaauBsCwuWUXEDUW0tc6Xl16s7vYufP3P11pY9n0RB+
xfG3RL2YVLDucJBlGOur/j31z/xOPdnxJU0i5FN/y7RWm0tbUlJUwG4qHHz4BXTizl8SOFJ+J1Zv
LCXBaQI9sSddmj7WYyC2K9bKeLTsTIRnYqlZ3W6K3WMYz9I79iemjtxKMRorKuxVWyOQpKQS4Sac
GnszP9fAK4uhCBeK+Sd8M+gSngIKgYPXngiqhbFMcAgy9xPDPM5GD2RXYBGVey9VUFXUMIVhcmJN
rLiMoKQktMoPEj0LDmUAK/sGy8bk7efRAQryKrG7MySZqTWNRQMi5ZVVK9nGZC6+C2Q8E58O5KTP
QkrZXzg8gyUfrJyjl6YRIAumx4CMHV7uqs8TkJDC7545zeQXdN2aVg/Wo2E5pCFue6GEk+ew1Ptb
DiLwuKNcBAWbXA1+5ROn1dxGYgh8s+b75+8sYiIjGabww6KGRfeqqAz9vUqCho2Xdts8LO0zuYH6
wes7c1Q+HX0AIKOXo7+rI412wvvSExhjgG341xRciIID3lym4oCUowHAgrz9ZpsmTA+/mtv3pr/1
v6v+6YkyjcJoNQ/IGAVkcB/5TpQHELTDceqEnhCIkz/RgNddGOoTsF33hCKAMV7ZCUQRyigFvL6F
7YQRLXTkTCmEIinSW4urNqdP4s+aFrY6Un+76j0ZeFpIveywfeZdhABpshsOfOZL39PDs583npP2
zT9yInzu6TToKqTneUahz7FGcjkLrGsw3EQTvzch0gxLuAlJYW8SHkqVv5VyAtHgO6Qn6pqV0MCN
Gbhgsal9e1Zm7GcCKionLjr7RSFYXRFLE+x6d63dfqC8mQriW2W9ezBLVp5Mu9d8wmMRcdY/sVmY
VRpBiXjR+Bv996GtyZUC9cUta57h/o/HKX2feI6ODlwqU2+1iUm4g5YT4pppR8v3sz1aN8Tc7Ro8
VDu6LOeAGlDqQi0neRTF4CRT9dHCHFwRWrG8HBw5VqJYFf3GV7t0jN/N/Qk6qwH4Zlrq1fbpHYRm
Q3q3vGVpjGEXwP9Kqn6uYBf2l1mGR1wl5MI3Knxkq6a7M0aolBa6kXtEt/krZ5+7lDDWQle8Uo+F
CxpNBQArQQXDsuJCAnjD3KVXf3D4CtxXqogI8jXffMsAdGmVr8SKaUG/mXU0d3QPvJKES2gcxLaD
ZgnpC8Rp4qGDF9g+qNjyqjbnDLywCE0eS8oT74ABLL+mmfe8oef4N70IVaDdbKPh1W/mIGAW6FCD
scmmTHnuUo6hBs2hvhHN7talkeR3ThhVOMfv3T6FjIslyYIf/fQZYrZGxAN4UBV3h+brzmasZWtp
zhyVZIarEmO4cejzmlR+zcceRDBE79hG5m2GiSDnsF6+uHktK4ZyMfb8CYnREHcNXW9fyQyXw5xP
6mVgqPGPp1j670VS4hM6JhMrsxihmTHH4cE0H08uh5+IwQIStakR2m8PlexIfI1gMJgbuomE1OwF
KdJuDPNu/734gaFY0i3Z7XzU/O4vnxNj+9Bw3zUn2pNs4FdbY/yvjrU9xK/FY+HKWZUVhL5TlSc5
PzPpYtgWiroz0/ycnRCywDNCYA1e6F9x0jQOVUmoP5/afRvRVtgJy0XvtUEyPvBAiosMRympIHM0
i8rENzwgsb+fiboEElCT/pivyxuymw1e1mGXnXRsBwMWi/P4aBGNnzL6NS78E7f8QGvccmJ/ia0L
HSEFQs6txpW9cJTvrYVsqPSL+suyLlFNxvdjpjs7hGzekRhzFGtwYNuUNbh9t+3PBuc8Ig6E4v/f
/LLK43BLy662N1Kru/wi9D5gaxyXdlFP0Fye7JmzMxy0q9x7qQ8/zb6xErEDIXcvso9ejfdaJ7++
zdsMhM+kfYed/SYe5udaBHQYu2PH8loeSHmCIpo9yB3bD34Gg0aZB7fBExeXxrS6eE8pzXdt9EFf
NWYULEISD5lBF0EIkG5zJyDW2+6xN1z5mx2QlAXi6ytUzZMSO2RnMi5vrbxSXjrIc+W5LjapZ9h4
eXN1mRexXD710eDRusrFRu47sbOUeeT39cnHoPzsNUVPBdf9FtqMr1UHX3IB9fDyUd1C0s1BgEeX
CWXB2TTqkWkHkfFebustP+nmBLoAlWneoKi/9qNqow/apsSiSQWKDwhQtGZ92irBW1+TJw2aXA51
qQsj3sPj54cIKW/4DVL7h4cMad22+D4cYaWONyFCHEvzDm2koclU5qlPPifc0sqtOyON/ai2AArg
uJdbCr0YOK1E0g4/NrgPTbtLzxKEJf3e9efGIgNGatkHGJGaWBUT/WyutZvXK5iU/Of7oQ8XKbex
QbpjAqm9zqigDm0Jff6bVPR8EIR5Wf1meRmkkWqJC99rDyOK7S/p4uwSVctii845sboS3DjlAouB
7d312/ZYPgx00K1ma0GePOScVdTw/0zLt7/TzMo7jAt3+vbcXEySgjQCDrycUbRuhGxukMZsVhLL
NjN++jqMph1YkqFhox5tiHNnStXfN5KFd1f+Z0g7sv8PndvtTn7EICWoCj1QZUFei8bqzT/fT2FJ
YN0NFyIYkAFFk/liW2GOtz3/b2v7MGS6KX+MRECMfunkeB5eh1DgzOC5h4+jn8mNxDCExX7Z6eSx
NnqO3dsKo9CmEoyTIrXsryiG5zmD8Xm/n7Rp2vC7LS73UKMBfHk4Vc28izUDYPauuB9jaF77Xh6E
jrg4uOpKmOdr2mjd4t7kXzBFVPrYf652dXiiNBK3KZxl3fi/VZ6muYIEqkz2HM4YvTcaWvO3NSXH
4CbQ2iwQc7wXl5lJ4cSoQdirMH/S5xmi6L8Ob8jSvgt+G+EJx6m3w91wTpy1YB7lsUBS769sNASF
b6so0yYwO/xTEs4fwt4HJNem/unrJNu2+pNUu4+1s9N328H+ZZpIyOnxo/04AWrqt8BbaMc6YMk2
Ad6VFUXGnsKfFBdhP5is2WNg6Yqx9m3wtxa/mcPUjXsLY/fOz393y7xpNlqrP+jLGDHtqmxrQ5gv
4A/JjGIAT7QiRCBlNBHSTgF69Hj3k8rcT9jxkq1PAoRWokd1DQUMIZfB6yyBuyKcgjmhLgQvRHoT
kz7PwWSc5ek/xYuU6cdcvUTZou1LVzySNXTxP7sg42R4g4W3YaygNO7Wxd4DQ2+XjVfIvvlGZmgP
JgqFy5cO3bV0Vbb+o97Y3d1xpcZ1gXmJqWDbITIVeOAEpzVufRx4nsG7YBHkAfay/3uRlLC6vOdH
ngVoGTSuckpj5qrGRZ7ydVEOe/vlu2raiG22GwVEGCBS2XKWwdMRlBdTV9C4DFHREQ4OaFLbnOfk
GPCauq8ifOm/Nfx+iFHgMMsZ91/Ceasi2J9TTnXOGG6HnkapmMx9g+QsrgNcMwMRhtYb52rzZHxa
aG3i59JjYrjkzu6HnsLgeosTO0zJ2uMxRV0Q1oJLLVolykVI6qsA48SInIWbSeishbTvqpoPX3Ox
dgo85W6STlJchH/r5DaYmvKb0YIRKgkyeZ64dxP1eN0ViqLVyGedDDIe4a869SYCCckDGnmT4nM4
Fqg/vsRB8oZUwoWGGYybGDSmagzRECQB5mjWGj6TY5ql4pV91i7QenShM28e5J1e7Q417+2NaV9u
oF4/TCOphY2O1Zp4iftSfZ7IqD/M4ud1WsRnZUwhchcQY/Z+gQ13mKmuBKxCFbdQWrMeDhq7SGJ5
3TGTCzSYtjgN3n8BxER9ARuN8XiKVptqrvUxGLn51GfiQw7MGPvSa/Vd0LJa6DvVxGdKtLVZzYvu
dn7GhsoJ47x3y9C2YlVLMRl3/6UN7s9UFB9xsRYw85yjZJYxXEL7FyPi/BXavPUIaU6C2PLHvtMC
JoKZGY9hdGf7yrpe12+4kAkq8S+lxL/8Q/pZwfzo+UACajtEl6Z1vr0O190Edu/EauYjO4iDQW/z
UeYHSzvjP8qa/WsfVbY5alQQ1qMmtyMvAvXwUaFA6o4KL+p6KTPNhUQ8M6t/xI+rr+PLfIEgd5VO
ZgKzGuzFOl16OkaFC1SbFRwqIjxxJp+HL62l6CW93lAvanIfMiVaV6MJXW1W8oejc15vsTGhbRFm
2zj/quH8GVSzmG0UWKmByx8IHzCVSJ6GfUYCklVrQ6jXPjgNa5gJGd4/NhQn1lyJXS1zZbYt17DY
kZxbUnJ/EGrPUcoHsSOH9C/9xNY1vaufv8khBBjKRYueQnzSk4g8UFotmQeRnpdQda30Zo9bl8lZ
ZAAJaGf2QyiUqbrqQKiuJsTjsBWD3Iye4aM8aE1jqNok0z2SzNGAFfnAP0UNUkx/4mMhRbh9qysS
DDyaVqayuUFF/uxfx+OhQyIEyXdj2FLu8uQ9VJ5XMjrUTqPDhxpL11F8Ew4nR2hoysmC86t0YT/s
9hSFJL3z8OMT60bEDKUsi89hBAbhXf2yaJPfSqXAvB9phZGIt393NllDfA1x7Hk5K1c/FDq9z3bQ
TY//Nya1HElP8mtVEm0uEJLc1s8MRlu4Duqk6vUhhoHAeFC4nR29S85qAAmbhLo7IxtdyCXzAxR8
xC8UKFD46k8W49xAiMutgcmlOgMfD8EEgtEpxBSq7t+ASMsaGUK1U1p0hulwheR/6QxBpASKp6BH
ZjrKA1HLIjldgYmbfUwz44HlxkR3Gn4B04oeL0M/9t/KZiR0Odo12FbGiG1Xaz2X9f8s/Wba6OzM
2BssvHDyCVxTHTzejmVSSIOus6DFR2b5K9LKPdUGc+THesGMWeukjB/gZEM4A470/JlxxgXfkvQj
7EACpU8mzrN90DDKJwOdB+SpDgqnKadgGmwZ9vAohvbHqTwiP+Uxg27t7uPYeeBBmc0+N+cl00XX
oVOqYHocrf0dbASvqzhY11KJ61fDt5ym0qQcznRfjJa7Av4idxyMIUzS7M29+TlejtzUG/+23V67
DrfPvbXNrdDX8ThzsWsMmnxNzAgHtRO1tEYI3l+9o60v7lgPVSP93J54OKdd0Jq3RReqqGC+9tUB
iKPuEuJHHHz0ATt+A3NFflX5Jf2R751Yuj3nxYDBXjFMBmswo5n0skTgi1DWZyzStXb3WOsmkN+D
Oa6FbB6dK+gK/8/xbTFOF2w3fmhOn1fIS4yjQZZKvnrgmgWG2u8E2NYJQsT8J8jy0ehlInagyyxA
xsM84dGY/BivIDfEIv/mgzj3vhzyCKLSUB3gVTO7NZRD9cRFBa40QyWdInTLyuqItbDoDJSRVaFl
k6CDBdeZwDOdHYvc9/bXLJ0f4Dp5i9tsehSVvk2TPyz0cF2wSvFkCxRE2LcLf4dZ7mptIF8BoZGC
gGf+4wJTVuDgjvfxLsa6Vga1ob2VrxTQBaHWP/n93aiYnYnjNS8XtWqaHsqipzLnE3PNly1ODwOv
skO/+ddO2jARRWR36PPIwOnjOA7Bcu2g0Ny66esg1d0/bvWzgnOBCS/TJz1SzlYdG1SX1Y3knj72
pEOIskoixS9NaieRUNYvjpqO/GiMIJbFsxUQgFWvx0tzIcifD3IzLx+gFxsECQzprgt3NawfRI3p
WCL0ElGG68C8qqxVgF4R5XgAHtK1plGmfgkDEu1QMaXfxYb4hTusMNSCukUhGyEqGrvnrukGbNMe
IRGNO4OPznxEJW3zmCR7YF/YohlboEHHjCeKOOGpmxBcWfou0g+37D/D2W57906C5yjAXfGDyOpk
fvGZqNXTXw5aGza56lDukfrmsle8uf5tmjJuSmZgUPZil7ftZqjrFsAGcnawasbS+jenb4zFldbt
yJWpvvXIsHEa2t4HEyiKPs1+9mqApMcpJTl20gHvFMIJBsRgpmUq8RAKTaH96/tQzQri/rGKnl4f
sRvgpXm30A1hfAT4uQGzIJBziYCFpAxOVUIIjiOIleZdSb9DE+PtXJiljYctwzr8Qqg11wA4NfaU
S+LIfHoE2Y/566MrWeyT2R/y9ZEaOXpbimEg7DYJTz/eRpN/reNuPuFEnH4qPstESb56ujsPCSiv
feZtH93hQjEZY/srD06nUQELjvWgkv64Vk9yo1qbhsWi6sfIBOwYIhvFlC4KJvJ8PX5eMgL2rItZ
nzhGhH1CG/NxCbZCrrKWFWVTbL9UqpXZzwBHfLNT6OQMZeHMwgYm4RLJfFMoEmmdrFFDqB5CunY8
ly6zY9UB0bCMXcZdCxVQQWxLxsnIommaC5Rx8iloglRyCnZ5Y7OtDPcU/LpQ17k+UQrVXrv0+U/3
cv2UOsSryyC69czzPpCbnFOW4UwzqlgOZGJ/OD56iRpd3vcdtNFmU8dt0yKpcBunnuwrCFh2vIUl
1NAf0otq5GZzFNQhUnKhcRGxERCEmiH52opai0hP5UGbVT2TzP5kCgKMfJlupcNnflhhGVAnBleQ
iimLXSO7nyWjHc3qmg9Zgzwh8U3mdk+i+r8xtTIZNBi2QPxwV1SOunUACRH9w9VRey6zStZSGrc5
teEmLG8QxDat+EmThtR8oH2aw70sNsr13u8U/E5MiQ4kStUeYMXdMG6xWO2jSnvpv+v1s/UsgIaE
ZkNa66KyXVCyUdPRWf4DRQOW/PVRd3yrKbWHZdsdoXZ0SDnOA+I9vxiHKE/GcLpxhFKLJwRmXKhg
7PRhNJMXcQ5+E+KSgiKXBztEDOtT/9gN6C4DP2r+ElvIEP9LqvPanY/vX2e/ycZKwIqm6IYnKPl9
tUiiP2eqaXZpImBLBpjFzmfB4OqVc/12QRV8BpJWa9x47FSsqqoVZ4eSWJ4RAMFIKTcMc2fGHnLW
inJJakqpo4yQri0jo3Akis6azkkWCcP2B0JHO8RMIYTDvYbhk7HQLoTtag2tt8LqZh9Fn6MlakpA
tOBnoUUxXizsUJFvAClj2SUm9uU1bq9XffkFNBG2JqOWiUn99IhnYM7P7XEcMOieYm4K5nbyuflD
Rv6qvD7lunYKKLiGRG8hy/FMc1al6z6S5GJiBxmFbBkWjgmEk3FOiiG2pdmqM9zG3XIajDCqRYon
ad9KF9w+NcSy1i4emd3TCtvJNHt3O4jvtiMnS3R+QE93Uji/fw8dcVlw6j9a4KPsvkks1X0yGvDV
ScqOR2L/6qk+MiVLpnL6Qdmyx5w5ubd5B5ruoNe82rv/HD98dtm9FW9QDosLDVLuXtG+I7s6dKAq
v88oDWIwKJLvtMQPteGWFULDIvYt9FDtNkmf9Mzxi88kqtULU4DGJBkWZcYvuLL/o2bkgLNHncn2
vlo2HThRPcMdWcZBtAQJtSzlNFgUVzuCDpBx/fukVBrr6NrqSF4RlyXfRoMYgrtKdl983TZgCnyF
OFFJxDLcsJRoSZ9Ji76dAEAWylURQlXY+tx1m88lU+NitVrGvPhfAyn/XxRXFcA7BrCbCs/J6ECh
x8Qs8aNjPODuVwMaa4XsrLdoQy+N3WOW+GZ1K7TBkMc6k3iwU3Xle1vuM9hnifSnf8zI7oQuXHVA
+0MiruKyOR6y0/BhjDMOGuqh8ch2vzs65fnjgq4UUbxcmG7k1VQrMAzHbp1pUu0RGYnJBT0bVjkv
YzPtGAegbYyYMagD3K6BwjFemcwrBHJLeqv3vewo1sbWC1KpWAaxA0fFYU2abc54YHylT1Z/H39H
/GxTuXS54hwqIL6t/NGpNg45sMinakWOozsURYNSfWuBDA3rqijUMuqD4fXoglWfetCcNMAaTPTX
Gt/NM0xUoNlHdm+/fx9tejmmdhhfGd3ssXBzTdZksuV38GpBo6WfhkQJ5h3FLBvR2spaY1lRzowT
CcmDPA79A50M7ewnCW7MEt3Kirp8zVD4/oh2TjV+jGMxAvEOVZr6zjNVsliw5mZZBFXmOYAQNphP
CyAUIuusT2FurSc3H/pPwu2xvL1bO1TQMmC05prHqmqXefaDwYtogzG5CAxbnwI/xsPPb/urQHaM
MQBdoKYGDRCmohVWI2nlqQFtbMnpf8rFsBVYtDTBRgTYJFM+uv/Qzv12mz1yGR9PG/GeIO9F5QPX
dad5P83RpQUZFI5OgmvyKmaDITXBCmO6GKeufGqTJxwbIDSrQJVntnqaRXpeIQGYhmZ31Cm7LrLU
QSplOZeWcNl2TfQw8nMwyaGLa541oD70nVGr0ra/CvtMfQq8pjElr5qCBPdfcVahcA+CCe8dAzFw
gXL0taPTdeAzbThSByrTTN/9UQr9lKyZWDq+dGrddpoeG5OKyUEpP8qB0uylJ0h1u5MXHgE6i8fd
H8g8AaqOvr9hHfXvKasiNh109m8iYEd3buauDWZsYrnmBqkQmeAZVOiKS0PeGJcPp3xVfXCVY8Ut
y9/57KGPaIWsuJhBZKbP5C0nqT82LR/uXXVrQUdx/8Lt0G828HWsVdcp22oYAJo0bAUvNyO1ERB1
kHPyBy/71kVOWY2FBHyTPPhPUfFu+ZZUk1caIbjow615L4krPdkHnwhYmoE7i4N586fmvACQHLZZ
D3CpxdleGxD7xqXgSAOSeIVdd0lVciuE4vc/ajMYIbig4uugxQansS76dMa/V4GC423qWDvGfyo7
+oGecVtQmQ6RvjdTXvdKaN+YAgHboVBMR24oUBDOTaKLsBwH9K/GkrQoTOnbPXHkgLFlDMwptPoV
mVZDplBtS/8w43UeeYZUG9VvMPO3zlve3k9ZfTMA24cc/CDXcHCQVfqQr62Z5JVjSSh5TQeYgiQ2
xF/PEVNtirDGTmUk0nXCLZjoSmzAKgsAipIGWEEh5SSTCAOX6aaDeCvoVX90/SN4GBOTAShFpKo5
CiFPvFGYmvXVqNDFX8YLOx3V6eh3vId9+kA1VC9Fz6b0H7z4Vymj7VKbiShTm8dcKSqhDwgO2d+h
WbYQGePi4vC7foaouMvVTz5M6bhJaIgWrsDa27Kw2+3WwzKsftitSKSRFAfvZq6sp6jQYZdJ5Yks
PaoVwSjfwq5BjjMqrL0qIXWQVDgDbtZql7O1egrkLj9pRhAQ0eBwOM9BPxwjjnTwhHVHI0Fwvij3
kcjws/L2fxtmKdb1WfcawvtfYOm6znRCqyS2G/wakbe+Np0KtKOok7z4MqbJZmEm+aW2XPGMw1TP
Zo1gByL22CvqK5sH4RpFPD6GHA2+sVUZ1/ZNLqrg2CbPeewJ7gy1CM6ytNSN7DYyo4ePwx9W5lC/
jBQD6tigWbeQXSUkidTcv4CERxDmI37C2wJjX+sYZ2NfIsccaZJ90qHSkFfiJxfY5M5MsWUq0uJa
zEJKDNw5eIWet62QjLjNpW2qe/uJlhK23ZIUg5k/Z/t3ghjNw83l1lMypGXLgwPFM/7lup1LlY+B
HOGRvRNLbEm4fFZ05XcFBK890roffM2WkPl1M1XLNWjfccpvtxyKyKMsvgOqMi6SYstxb/aVMx8G
3w9ovRZQl/ci5AZM1IbULqz2L+IcVzRtLFXGJgMcX0vEiM5H3KC+w4sOCW2G2PQYQN+jL5428GBq
E6ARxS8Y47s+tnegPwSIG3Xu6bEEUxtZ2q4YOxGAfpZ79vt7Os0QOSww1e5+MiyvqJaUs1NQxPXh
RVKZ8PsBjw0AcBbhJ0GFs33pVHkk7JPCcUC15M2nuEaWIJhNQUZhZVY616x/5V1SShH8gaVyjc3e
JFkmym+Q7sOBhXIqCPQWBrdfDNqR4ojF1QWmUS5dGo073OmY5p0nn7zGTrMeACRVaQ58FRraexOr
yPydS8YhL0g7TxCTkXWFafkQRS1em6LEcwWKdkdb8fleLB8t+yAcZKflLQGSYZ8onmvwJLEJDGni
KN6kyYeHLmhXUh4uGmdml1uZdvHcK3RqY4wufMS/x3G6jVZPc3mK14Isp9YayAWL2nIx5zOf3wIb
v2abeoJ5lWx5Y4yjoFaWxILuJffDWjdR4BoKxKD6XZ+PzAmS47k01i/KhEcexN6eYWJggqZfFb7z
Ti1UD4xAANN6D8EA5pOLyVWMEWOZCUTN/odeekuVgpBaEPGsHo1rl/u8SYuPGFlFsf2pTo+qC8pY
vLkGdZk0CECAYupruGQQmEysi9yMKRmLfUisuDq8fBajgXxc1RYMdv0ulTxfTSqrZr+sZ6ScQpqD
YwkYIGT60TBLFlDRA/RqLq3idv7is4Y4RmQJcDnRcau5iiW3ATgqOYY2T1Bzr+LKb91ayqXZG5EM
sDqncS4AnXUt/9keYYHywTaZ5AYbu2VGLyXYP5XLRzF/kj2Hk8PmCNHCyvlLJlKmqGMUNiN6H0iO
/EDP2Z1SelHVatXKlwzIGXxN0s83GxPLrY0zyixTiOJnTX3KjtrHm/LB/yeabHReL2iiV1DlpjL2
WtptONN9ZSEzWhoIZkpcfboTH+J6IOrYt7U3rxU/HnCCbWUS382ZodW8nUOE14SKFIsa0geXJJX5
uRaqQrb6RFQX5AgBZvp3cD0tx9dEJg42/wrk0N2/j91BP2xMZL48Q3LCYHkDszv5ZHV6VYbMyaKG
wC9FgRKYk7R/QbHeCsGU2NHJqi6+jtDCTol4YxK3I53nssFipYVx4w45OQ326bI9IcpYxHkN8K5q
EWWCXj68hKGtbsjM43DdFCkAD0bCk9HGIOSWBlsXLHNRRnzxKMbwl6Nsnxus1o+lcDZyxSWg0UWb
XH7VUe61YyhNLFfu4b3cJJx2elBquIe9h8jcBsjSrRBn7znBdm6C9VpmgYavOX3SW3DYAxyZREBh
i1uWlhI5twPzcwBCEcaK+7GBzJE4mPNnZnhwj8y6nKvQyHnB4amOHRcmVZsUS/KgRbtkfar3H82s
Prl4g71oxzshTvmPFB427iR3t5Qr7rxq37gwBe4EFLQvzeeFfHhzhVTwjKVHC/VNWzDiIa4p0uFg
BdtNMS3o36AwnnhvNmQFszXEc90jpYrp5YqzR2+i6P2zK0lNJgjeZJgk2OilNak49GjC+bfpNt0j
G3YzSt9cESFfd2QmNnZAs68NPBHJ5x2AxWXSHGbksj7IrDOhaXNnuddwvvbaVV1KXpZZW9XnsDaE
bEU7SkL/ym4TqBb7RDZXJRVaPhaWpR4MzdXaHqG/aVTxtS4O4WJTrvJEU1dxL22TgSJ08AgRtV93
TVKJnfvl293MInQJTQ271724qQ2dD4Tm/n3jsDOMuGo4VbwjqlM11m9eOtLY9gT2rZ6LE+0ZtyzV
9zalaQj+OwRIoXAJTLM912VQx3+/QYCusEdKfx8KSId0zJFLONq+jx/C4g8Stj6RoJ2otCfVXK3v
b+XZFMDP2sNPl972so4ZHxrHU+9kUbYRsojdgFE4wLSAdWPalhhl8a0x4i2We47AjvLIq3c62h3D
GlZPeUPSh1hQncuX4nAXvZJQADANR8YdGOYsonhkBb+qXh2oOOXB/4W8iNafO1pOeUr9DlAQW21E
NlX0fbXT86m4RACVgQbp96UGj9uP9L/Z8/lszQGN9dFwN+g9PEJDLQvi1Q8lQPfitEQALdyHN43T
2uVEkKqbpxrsYa9lFAsX24vvTrR3tLG2rkvY68rz0GykF8x3rO2wtUhEOtirZp2MfhvWjIqmcng0
Lg3DP9GfbiYJMYJsNpNtZ8H9zFDb3S0eflZP/lrIlwrIGr2VAXq79Yb8xznVryEBXJfhirQXQM34
LVGnuTL1aKKeFPCZHS8CVWTLmGVl3whscoOZHIbthax2I8Hs5yeNyRT3KatScqGepbgNjQhOK5z9
upSXx7U36/sK2PLwkFnre+ss5jwUYF5hAY2UxsaHPUiucbaFWr3h9/5Z8k8Z33lROK5otgx5KBDJ
EZLIKix4coK7Q6AtJtDZdhMId+hw/WDCGDVdtwEHjCmNxPrgiJZMLRPdGT2bIVx6wk8/wcV5b1D8
m7vg9yeWhEoLGs7YIWH9R+fK3YETpQyarHkQbhVUcRIRwmQXDIM2S0Bn4keBaHUJmprtxBjZqwms
tn6iRxNoshQj45+rvmDQNT98XjZwJkuQ5I7MLYEV40PzqxzkBfVG4C/9gaIyM+sFOtaqRuIua7wo
Sywc86sLdPtdcgdRqzMDyjbmK/4Zw64QYCH9fvt4QZulnlKkyP+MqVqg/qtE7vBb9npe7AxJG1Z+
PYvpkkn6e286EEUowOC2F+mbYYaTx652u+fnGCdEIJi4eZxYUP9yKcaJR/90yPsIVPr8g5oOQ7Q+
mt/cpeObMP0Jjv6IXbvMCUJKv90/VfQKNGhiFOyNag7hA4sxar/C88IG7qnRckC3gaGcboHO666d
GtZYgx3YHUliXWhK/pozwAQRwP7pyiPqXTRwkRn+ogePysUrTGPOZ0jVpi1dvybhVXHPIFpI3KwA
SxDsr+NclKLZWDVGph6yflEj8KNMm3jNvVkQC3fBxZtzYI+fSBHWk0IVl4Js+Tgms1qeWw4dECn+
tRQ3wl6mZitdRetzHk8wm8xFPtM2agjjmllTg7GkdvNbeViD8mudaA6z9Xu3b3ZtcPTOBgjfaZ63
SCOshwYHvSKN1HJyuYUPef+UvrPE5cGDrMH8JX+kNIQ3L82TSiEcfD5MAGUoQ+GdNrdUnLchyRwd
rkSmnpieQM3MmbvMEdbNjTAG92PPzsmPw+S7PQxjSf5Pqp7XYQEKOLnFqxM2k1l34ZWSSNi8q2Ou
idSaU6ccqSl/8qFZMi6ULdzuxqLbPifOd3blA+Py4v8q3bTO7jEfFXgdE2DBL7DKyUT5oqyXzfhW
2s4Nz+uVwIR71HIz7GaBTSnxch6caOn2ftrgjqfeuvk8MaSbqd3QDngk+HvSQfPeCm61WDmwFtGs
rorI3yW89kCMgGt+iWaInWn90JDwyrmIRb2iGtDrwu1D6uvuztHWJ3jhQNYpZYVBBNNACNWSXwtd
BhMRLCbT5yRNcWtjYBj2wSe+P1kwCT2YyWxB4nxJ2LaXx7/zT2KxMl9J3mP+DSfWifRvH8c72oZV
U2wjfm5u8Jy2N2lDYg1nx2ENdkdTcG1thioeYu0kqJBTx8WACQW5LawLLpGE2KIKIZyZC5vfmWBE
YANLZVxRV7+Avp23K1Hham9RdIB/OFvdacRi+ra+q2+5eWR2qiEmXwN8aXAH5BIKZmaICO36ndew
LqAeCWLt+v15I0DjwuURZv/NZ6toY3G7ufzUQHTFxp/p0RzqmAMv5QfmOmqM7ex/ZE7eLkczatdv
gvSmqH/VbD9X3Pi5kH2Jhnn0aE9aJO6wGbDaC5CfsTstIWBtUsi+rMKZQ3K+K2Vb5SEpvCbcpcAW
yRu4OIeZS+gm8feVRMUzB3KykKEHOCT1+aqQSV5A/OVykIfUYAL5NYBfJ/14bnGgzG0pSF4Knouy
i3586b6hdYs+dfhwdcCA0oKz11Dl7ZaFXxYd/9BqNOUEsvfdubGU2/sF0ICXoBj2h8k7qxKgKyKO
yqwAybB27HJmasAItiXeVW6iwyzqu0NnEqStPsK6HXscegm/Yw1C+jt9Y0kNz7e5r7Xt5cNXQtGL
5aTQxhZlqsKcSnn2Cq33pDD+dnXcj2zGOJ6dBHrWhVu4uyVKv64EPeqSNoQtfuNzGQUAsrhf7umN
rACWyRDRuwyGdfatXMDEbuuO3ovHuWglCiVdKvGHfe3rspreft+AOXRNtJFEeM0B52ocdCEXewLG
OJUK6jyqhV5YoyMQcaFcQb+Gxnic9ieEjRjrX0e5AERCttF7xvLg9Ls/HrycByeBBgkU8D6qv6rt
cveufktN7BnRPUSzghZ5w5kRDhl8z87xYssW6TlrHmrSLjgUGeAo/fBVQLr7xD09wA8K8rA/dMGg
JTsj/0rqH7zuiju4pJbDRxppnhV57djNS78l+iB33Wen1A/o2lEjNI6Pf4Iprd9MGZ7LqAvDsivQ
wZAhE1nIT9F0EP5+U4nn60TOdOMInPez5HJNwL9hze/Eg2cGTJbWMQJQGuoblFl4B13K0qJQNImJ
ibuPei3abRmZ1Xj76cO8vbRpRl9cmWZGvCv0gC+838zzeJ5xip17m917+suux89YIbrNpaWPrxWC
uO4MIhcs/ezN5XfseTdV7pSPO3am73/frDN9EzdUE5pWHsmZyh5vGb23+Z5351m7ZCHmAoa02NWx
rg6Xt6Ipjw8J9r5tBcZwT6qMorthpYLQdkuTnVyiVJuavYoXJ/p8faBFjSQFy6ijLkhpvhnW9rLR
riEzFZGQJyK+TbC1sK55Z9PukvueERNR4Bd8cgv+8LtQrPOagFi78h5FKPAf5rhXdJ8c5YbKSA8Q
6GgokK/QJHj8i4m4++gNSWsteh/DyhPxZA+TVMXCe5ZIP3OFICVW3ucSg2/XuTs/hnfF71BfeXXR
8TexLBRDWZbPRxobFNV9EEMjBt0VMExtiEX4iODIeqWQx8ycf+MEEyi1YTnhDzsCCOUNIyv1yeKr
oe2EipwvqPusszEMjb/Uaic1kmG0BkH4Y0qghmShd2cGjmXLH4J4eg/i3vD5/TC4po198qlwTCf8
a0c77rsz/Gvd29r9FXlFdtCVol7/S3mqRxpVTCYM03Jo3LCeTOamJ+sEFgmdrIlnX7YBPxJiaeM3
sBVE92nRH70ZuGbx1J4AtEX0/ggrZ3hyWykFXsR6Dnn2ZRlnKpCq+54vkRM/x4qQsXPpsYivWSbC
ccvr4H2sd9p71WixGZaytxG2T9kqTFN2rG0VBwAM3vIH/3IL0EDf4GUyT49R5Xjr3fgNSqrI+RKL
YiiL04Xn+1gBX0/d3F4Io76pu6SBapepyU3elS6lzLDihRj28Sj4yA7yt6srcs2o3TGVRFSotumM
VVwnae0szBfDThYmt+Smbygioo7MWco0jTJDBEJaNY6rM7sOcGsyGlPV9UWV8KcC7QSi8kO0Ohvu
1F33EiOkT3lYmy1jFnIL373a1Huff3zinyI8p77MTMLC4uJ1DVshPPFUFA17cydIV3FtpwDwaQY8
9jN6YIUtTwn+8+eOSYJoU6icIJiTaXcEZnLHnM+8hVRLLKWWpK8VjA9yf6XOfdlRuOtt1osL2+NB
gBU2drJ1rUa3Pzz3kS9suw3SA4iPuIqT8FKNvKytySu43jfiNeKOLLau+T3fQVxZx50sA8J50cHE
KhZcu/iPM9tNjpe+q+t5DAprYRDI5iN48k0JRsd0LZqTM9pAmFl1Y2lnQIJc1vvq6upBIpCfrr0D
GhFhvrxNa9bxs0DXXDpFvYC0Fi0JefJ9T+7ds1MKf8i/zUSLFbrxSrQUyRLgibVFoeypeaBN5YZy
haAXyewqVMQkreJ7jZ5WTp5DAgH/wrlmxgle2EyAd3r+BsSRKnpsw+tK5dFIm2EJNkrVs6j42veZ
mxXPEVidNxL0YI+lLY6D32R422nQS4GgNUvAQM3w0+cYgBJJ4+akUafOXFOQX3tmBWbr6kMxN1T3
2Go5AD2U0OaxvjXI3/dZygWPvKYWqoGvTY2LzoY0u7H7SmHLeLrqZxhS0au5dPHWq4WTCa+E4Psi
oXlwLSTDFnW5Mo66irgN5PL9dTKCJCkp/lJRSxDo+HuVLHb+FvnEXPPJeAZrbo1N/n/6ZxNUjGci
HEGL9WMK9SvYAd2KToOLo0E9tgrAEeadBYRTcWnGMi7cZRD4UN/HN2WdInoyWvsafQbvazpG1rRH
iLMr0gmzKBtX1GMxse6Lkd4EbTY/suw93xtQaVLRmagIRLMWy/X7KMIX+9QZ913EX7tg0wEHc9Mg
PQ95uYa4UnHvmpa4ex3ES8op8fmBHoXrC/kyEAczQSiAtWQU7z7hRtlvm2kRJATUl3n8ydeiYaAc
ejwZhHEVe3btdJyVXxyWEVC6eOzF/LA4lmTsLcKCjzTLhSpc3eOkCamTv9dfUuhzWkRofF3wKICg
Ztuv41zYb+Pe7B+PTI6UNRmJrNH9NEpX6GYNUUFkGFu3zFgNdZ5mBVgZECpwpUjjxzP3I25tkc0N
GIowahYUm9fniHnOm4FEKPhYVwFGF2FmVlpoLFrfzzQ6bwoiHpMuI0XGTc4Eeoead++cRoTq1Upm
LP+oyIk3vLo6rI3TPsYQ2HYVOlwDJ6Ajg1Rwxsfb8A9e9DJhsi8iZmc4hevJ/T5XnHTg4crjPOSR
bAK8Va0mbqJ/CL+y70yyolvjwm11r3BOoDftgOOsrnQ1mcllWC5cAnr0M8iwSYf3Pqb2192cDCal
MuDR+9+B20ZdK1lyFfSMzS5RolffmIjg1nvML+rtILsxu+rtBA66Ct76Sd2aFD1whJ/oQjc/iAqV
L/2XX0PZ/JxL8cBY8x14YHSts99EJrKEQ8PKm0Jl3CsGS8c57hEegtzUyGz6TkhvKa0PaHXEjM0e
OWdxfxLUq6tOwoMRjClnj6+bEuXSP7a32Zsdvw9mdHMo/tJ7IkrlHAOJs+eMzoOnlYAsoPTktwYf
m+XMVq+cAp7KLbnaLdtQkUR3WlAyRC7JmWrt0H/C8Jxz0Ks66373dFZAjE6BApLo9Ldyve4+tSJj
RW+dFZgRcjdap4QyNeyVVAdHmt+MHa5z0gJHl02faV8sZEPlAQao0Tb+gH7AYymWUDUJWVaBysKJ
xjsdH8H/kjGTA6dIHVT6pUfP3CD6LDvpLSQlzTTy2If1PtiZ36e0iNEdeYwv7ewlafSChlWMLSMk
ynUzyg1RR/1o5RpHDP4WUMH0Z3EzGVpvsF5pVBdEzHnHBbPD6N2aupJ+QoandztdX/EdfT644qz/
8ZPh0MXxyVHOgIzmlqdTGc4L1RWQPWfe0g1d+d9dwizW2+llhiCFmkEabBCjurgm0GEC52G4LSY5
ZRJ+NV34Jn9TDxoV+mYeMImKXUZhWM1PWS6BDlYp0dACAsiXObMDPGohEEh18LaHEoW4eXM+Glp9
udORlxlZs3Ptl8gQkFDDfdHwG2sAC/qPBbm/NY84f4rvm7Y44O1FJfl75inrF0QrMBWLT5WeYVZP
R4O1AOiRyctkJ92qYcVzoHHqlLCu9kdfM1qTRiSaVii0TbTljwHZdJu4A6LYGH5cVjyhPtyFvcid
l4u0Z0eYzPaQ1a6dvf4ir4zo1guGq/naHQvQb72KLQEn5NOPvWtTQe2U6REwY4ty3Eqm7btmZAYc
QkYi35xWGHTO1cYcmQOys3Hy/jw+ajHmIOJBglKOZWxN4ejACYfCg9v4xNqez8XPerNUkiZ8nkKE
ZTTg8qmA7aCeHAHGQ6HpTWV+1fYxXdLT+m89wcclwbgN6oLil2uWLsPIlOL0qm1N+ZKkjYNaHxtc
Ng5f2is2Irqu7oE9K4ru8pQHNAa80TZ3y0ELm0GIclOWYJMCkUnR9iniCXAzdarXhIAZ+AqIlEJ6
l7VWn4PeXU/qzotJD0jXwpFA1rOWKnXjvwo1PrkeS0pPcuK1DRaUTmYoHX4n8FkJ7GnTdFyyA5rW
/NgqF4zUjFsm752DMMB5dHx/BZGjQ0pMinLJHuF/BgLJyH1bIUl4Qz1Mp1WU8hG5WqAHrZodJW8h
+yPmkS8HMFRGN1HtV+6j/LFPmofq9PvKwJwFe4TiSeqVq+z2eGFebXrhNrxyI0d7ujOWBmXKGP2T
sYe2d0VbWbn74DzWN2giJsA9QYmaXeCEfuDxe+G5VqD3wiYJlDPE0GN0GAqW0avjNvvQpOFmLDxq
83UzJ2Nwnz4oxvqKG5QFONnRTUNpx9T9SOgrE0JqqyAoue4QohaQEnc7L84z7Vq1hwdN+UBvhwyk
Y4KLefsFN5FFa41ONAa+RkVSZUgsoaFj4V5TPlEsTwkFcJ0TRitpkvgJsP0UwItKV9hGv5bYplbI
13Gqhgat7lM7dW++2rbOGXqgdxe/2f/By/xaGDkLezwh7DUUNqJaEs7QI708Cz1AO95gHaMYq9Vt
SyT+/xu582uPPl6uqFZ/8w+R2tDx1CKVNgjhcSmHBW9UwH/ZvCm/0v0Uye+U6EgC1DQjLW+Ehf3y
CnggXatkTCUeoGVyHdDsDHD7xFpfFGG8sWPPDCAyruoK7RTOjwYXJypjtYXD6922rEEXIzPfh2bo
/whuxygm2Uzal+sMxlY8MRvK5xtVZLquDgUBjHPYpuxllvZt9peOzvlzW6FTkk0kPfZXSR6pmBJ4
Ubf+cQ3O9z4cOnOikgmlcrFGMoC4zoQZbQzrSU8adxhWStCceSTdYKQ038EvRGgtrL0lGTRDI65W
WF1CntLx91sePHf3JxUtOCS2HTH+bpi1n664GwWCFkgZAGX2GkeyeqiFrh4YVHWtEhmj0PNmlu59
pP5koaLUFDksBcyl+1MS2rD1/WJ3OibOQNkUi2X/w9kR49sk/f4qsvuBnLF9z5BJB6c3iZ7A8Qe1
33vUYWyA7D98gJD0mAtAXyJiJwX2fDkqErAWO+Otla7GQRBYWVICjNNiFnZm+8Y9yFEVi2Ad4ayw
sPBPzv1UaMv4AHAM0tY1OJRipKwbZabhkxBgwMn2IZbX6la/zLQwWuSjoysKnq643jN0WwZgrpm2
xu4qPZayr48NcKip2Igxys2i+HOimxKZ6I9H/5Upnsbu/86ikN3XL9dP+e1FjjultWOjs2f2IMhn
tl+FZtI6HfDxNGuVswE++zHRucIV6J4nzTnt9CWbnkuCCefs+KrPbKESh4vf21S4/iHRlKP9Jc1a
o3AhpxeJiuOOrbvCA8+KC8/HMubm1pNk8WCkNdFA+knT9qOgTg1pO00dphM1+ZUcRZZbHU1f1TJN
s3BQg2T3DsbW0rNnOI0iccssHlUlpziNkZq02EbEahIoFox3ekPGi5ObHAE16OygbtmooTBlBj/l
EbjoXh3MoSYC0Euv1EFmoStM+y7KAjXgI/wAl9I2i7gmwBNz3W0qAZccTxLQzQwBeUBBdLuY1Evz
WVfR4HTLSb8+YwUO3pgP9H4G6IRYkeOPVxh36LRP3XEhHMzBOuVj5MeZdtCjt0928RF2UEEgSELm
rQTprbwoMRNuo18sDdBt9p5FfvpoFOXvk4Czs6BUwhmfc+6MjK1dRwSpFa37OrUTOjMUHHreM+Uy
L1AMH3VgLgBo3Sjs0NNw4TPKMXfER30UE8WT6ANgXKoi/JFWu5cthl76VqhUMm0xU53WVhRkEgFk
GP8lGsYZqqHfNWbSEkeiGGDmQqau0WKACFEYE5N87rFjPRwS25QDfHn9vF86ePIUOZo9PQRwew3m
d2k0J1r1C9i44DcpxcaalbagQtYhfg4Fi2oiaQ02j2QEpRvPpERI8ClkkDlIqw+rm/wmFz3kV7BF
cSZIH9+iYj3flZB6DInWdgABBkRYuvloP6aq1Noc+IRaIHu1jyJSaquH94qW2O39sfvskK5bHCaZ
vaurLtIaLB+xUIR3s4fK3P5EaYMlOF5TcmM0aknwG+AFQE2n5FJwZXIynLddFoxclq3jLdEX9HIu
6LIrGZblZGr36/SGdr3fI8mXDcdozbLMb53PTjTo/YKZWWK5rSHMvKLc53rNXAjzUthWPJyP8gFA
iMAWjd0MKnT53sbunGiHfnHgV4s2LUs25GuT8Xmz2LYhWff1zmoWhuLoE43dHYJrpSMUbsVVdA2s
UfIpgffDm16P+9pGjtrBdXzUsWDBIstbL0JC2EPTYg6t/F7WJ2YRGThX6uuWbxXos9Htf6lrEzNj
4cizzbXX/wt0n84vUL6CmBy7leGg8pld629wdnJ0gnmiBiaA1bt9ZvHt4lEB8yDt85nVpWbsN+eX
PDQQ1ylOQHrnjV4AB8R/8ENW2dRup4myevDCEWPNaWcUfjHgERocYzeFe8CX0SMIDrdawzMSQwHx
aNkP7R9hgQuod/hKbG8KNN4T+9gj/4zH8zkEq4hpW+dsQs2ZOFy1mrUcb2SoaUs2yvfEMcmvzfNV
moGIXOoVuaB2AuofNA62YgqP4OcTv+lkIrBw52CpQgirw1pffG1n5AAhkrkco8vbDh4ciG7EEtDc
ENTLIsNBptswXvw4GSMp3QxgxlGFrx9YuF31/ghoysodJRwJF1mp3TX/sBdSfNVbheA8ifbd1MaF
j03ff7sPYIPB45CRMqkIjZIKQUJe6Ca6n/pV1l2Xx/p1fY1C37cf029ADPA9Gd2me7VnqHy4zbl2
prVIqOPCm1q4n3XsnXEt5XYdr2OCyFiCSPPlDG4Dve6dPCV1lE+Z9jupLLVK8kRbs9RFXlVbG+SB
yfGQBarMlfUaZFw9aOoigjLKp33WxApNFEVHxWApnaWl6Sdye/2ConBw0WaiJvDMEmXLjaP29gQo
VkpSFfWTT7haoxZ+TrmvxiMhluCFwz2XHjVfFUVwl4UNyUoSuPFnJ5w1UVAwoNH0UxmV3UNRXIN0
cuEhq6FzY7KkVHsFldlK1/2eWXv66UtI4HdrQ6DwJ0bd5qZAQiMUBzGB51kyYJTHwQftabeIdrMu
O4xLmX1eSKSt+biZ5hJAV4b6aEHMT2iUs/IQfg4YXPK/LAjEL2yi2MmS6SQPb/sDlUDY678MTCUh
jIXc8hgtFARucc6zAlVBMlDqXcZrf8hKLODqGb8Fx1xFa+oLLrnS8WEx6S4xTR1QGn8DFSVbjLyr
dtDzC4fcC2MMSOCAbgfz5e5ggivRUtLVJSaepQd6nMFGMxQE6I6DxAOs/G5Uz0v4yO7SEDV0kp48
loSg4HehyHahQtPMmK2WXXi5s8xB5dUBVvG5szYkkqmjyVDyIxKHTl8qbFjRAEot3TAieB8RjSTl
BU1rBwQImDVZaY7nDugT40Dipu4+V/DfRxZj0vi9tc6OECNRNgiTcrB/banY/sbA6aPim8GD28Ir
J2uow5Xl2CBCZ7FZzY3FU43YYshP0L5Jc6OtQjGF3r17AusZdCzV/9poZ5rcane3xtf2EjItCv2t
zmvGVK9Wp31rc56koghegpAGS8dpuAVWCjMLcnz1iEE6rUgS1dV/OanxZfxkfs/YQgxr68mmtdgM
kgfvMm1fkgN8Hl3jHM92LuLajuxbkATgbnsHAaE5B+bL/JqR7gIah9iDc9M3M5V9OwEcWRpuspzg
PMdbhz69ykCivs/0IXm/l5ssYKKQ6mnU5KCkao2TilGv4kY4/OKZpWYbSvkdtaBs4a40c/nQf36z
fdl1brKi8R+3Nz4dFYq/3n3nzzqwrq8FplZ3aPUN706BNhM8zfAOAlH2RBY2l90oZrgmaNqapQ+a
aQOz93fLt+howzzb+Rb9CGbclL7RhnSEE28YbzEfvJ/dDh/kyxx/tK/Hd9N+v3B6U8QsuZcnz4ZY
CDnWvct/ZjSz5LDHn2t2fOazyabtYjmazUpuMV3c/CeMvabxqnISPSov8mFV8NgyMl/5wr92NEUH
tlVCpXZb0Vxx51LvtpDjyYaB2ADgKJFjADaP1ooV2DY6i19lJYXeLg/b+peLHTrZA76rDZXW4R4f
P3XAIV0lkL8rMyc+Pf/cuv5oyvd/1F+FL+e/di9pEwZWnUq7ha/IKFLZmgphC93V57zuMplDWurm
kI5YU8PpR/RP550wmWHOczmy/pqj5wAOigiDXzkVeF/LN+SHl3hwEpFJrvlfqVd8l4Bv//71MkMY
GZtaISGvinBfNORzNpEwWZGCG5hgIWb5WkxlzICXdDUCkO0a9OVSaoe8Fx3H/GQsMZdOPYLnwfw3
/9qu9Uj/WPvbSdSkwnzpJcGr4PcZ9kuPcLwUIDMU0dkSP3f8FPecg92OiNL5qDjjdeg81llK87R+
lls0dKbRCkERM0IKQsF3M7FMFwCEkkPs2Ns6fa6VoeJoKFM7/ZyYyZH6j/VAdV73vqER7K/xUBbZ
4TT1UMNWR79peRO2IIMFPGXI/WVqN8Ozp+59wXLpskTx9lcZ2gYMzet523S4Il2HI0LmsF9etgOs
HSLx3tWCCcRS4ZE5/3d+55TjaADN8BAWe3GXft6RzH+yIvkPLvcKtilups5Hq8epdU/3NaZ/Wt/R
3jbWOlLK5SslwjYhHEpjrPAF3rtc5VYGRMoT1/0U5xKXFU5cBMKQM2faM0HsoUS3AItRGKRwiXi7
DarTh21vuVbrmy1pO7zVm9dkYIlw6LboJx2TWwfX5kPIrgfFIhVlGi49sa1HfwA6OO9ooTtuhfv7
PRLCmoQpRtG4Fdlrlm7ZXwjJFIXm+HVewkvqWSH9x0kJf7hi2YodAfyfIfHhP/9DxItQfsZCyKBj
F452yJjOwMcTP3rzWiws/8DCvFNztMDRkx3uhVAc0WyM7YLQZEBx6Px/ExTxrMo0FbsNmQ4vkD8z
9AHMyuBCtlEotQX3YcqwSDvmRCqswCqSYkN5qSGTO6U3Wq+0i+nu3N4zJQDbxD29Y6e+30wAIecY
EXxG9iFaH5c8DZMTAfhxkz3LcWFtTZaCa+Fe3huZwpnq7J5cEojK2aWWgAKV7nzMPTkyOnBFNIrT
6zxxaFf91RmNsyWvCniTXFO9phRKJTkoyqPn6U5M9qz5uaCrImetQRxQ4lam129IyR4toVQEMwj5
1nxj1D+MKLW4QtVu5DARsY6Apx384QWhCvArInyjzcS3e+PDNBaHMcRNR8NBWDk+E2OIEks+MR28
vM9yVY5eMzwsnw+bbMtuwN1U5n5zgR0ZY7IguotrOf7eKEt02Llx0Eba6wcHkr4yHfDgKzQf09Ak
H/cuJjPZ0CRGZKj9JYtAv8JMGCamy2Ge0uYyZ6x8FQ8sa3Ig7VeDccdAIBlYMHq6ZoopHsgdW85D
nU6euI4i41svWdx6crWxT1SgE2XHtKjH3uPhgwL/jO8Wg0sPSyYvAzv5mjn+6Wz4xSm+3Kr3KzkF
3V9oMA9GnRLbA5Y/Ht0/ekw2Yqp8f4jbujmga2vu9akxPnOkd3HbJt5nuEm6dhAdy8PBwwlaaVrm
bEI8xBVwmorYiBEAob8gHMNRrbEC/IJxVHiDWY2Nw9aqHyrNPp/r4dmkkgMsGobPvqZ6e0N7m97S
H3famjN4Pfk3fenqjuGUPhB4gygTCiik20iQqRu5Zk6IzumSPfkixs8ZuJSsok2O7E+vW9Gehxs/
j7cOIjPA6J48gUvFCpsXlnFxXX2Sp8OA+w4uyANxtAMuY3W++vu2pmm18TTPnRXipahFhbQEJez6
+BXp4AVyWU36Sl+SN3woBXn/yhUeKjyaAtI2r9ymVYszNq4g5v+iaTiMjdBaKRcxIY1tiy2qktHx
s2QviB6iQlWzT8RBPzBQ2JoWXbleQJNELYoNb7RyyAzqbfddpXlCdhjaMG6kBsf0dFV2sUNfj8zh
ku+JHuHLCzXWrCexWFD061zejweq1mkAEVLfDd05b0p0r7nQ6Jx+HG5WfR0WskSEgT8WhTE53YGl
u/R/GNtFW3Kd9FmEfF7Tq2Avj/ptzmnSH7EXi42PjZ+dQq0Nd+fVm+ljSunckEUM/WebRaXEImcm
FszeEDh2iTC1AoR4qabS8UJkg9JxdtqOyAlrRuVXi3vxUmEBbZOonQ3vsHZMCWyF4ki/OXRxq3TL
6aV6Za/Yi3K77mRlLC24z8Jvo9GLVQ9jgJn5QxdBJzCX9ZFGD1wYPFKptob5ByP75a0v2K+9euD/
4U7P3y12n7ZULlkxkQ6c6pbieDBaZ1g2Y1+4HZkM4m37hQnYxV5JNpJFbXHD2e23uqxPc31r+fP7
kV7Hcvk9huLpNrKx4rB3Alc20Fd3zbGeYCyk6sAZboLfB0SrFkIMqtvlMNaKinqiIbgXyLttD0kG
DuLx4ELwHwiGYl0RIoNKRdGWKD58WW53dp+36Fk6R6Nc+hiqnyMUT8Hv2sGuYRZEAjmt9v+JqgqO
iKvtw30j9zuEXdcW1SYsXBdGAAllVc0YGXAQKx/ZH3gz97eGOrTDFjCJyf/yTllQ8vYMFl4LyB6T
9YtZAPr7nTuv9pugKb7Ybcqq7AGjPFNldrSA6f+OgsHx0QKtscLajcE4SHRg+vkXoWUeDSYM8R9V
aqGEZ+a9b9MDN6MZIK9nxNmaE+iVNhUqIPbHb/K4SBj/pA1uSseNCm9N9pYF2wPp49jvH6X941sn
oYeMrx8Ic7l6bAy38/siTtfQgMITWIo/kwfKW+fraUpMURMp/EMcIZ09re4j4Ol80C9w5n2A5pJL
+Ciu9d/9S/rp6HEbnJnjd1Fjx75cxIGqtV6g/zY6LCQl6lNL6miJ5mmvdXL6f/96Y+F8drU+4N7R
cnHfMvYaZ3+7XaM2JLquoDnhgpEddz1UWDVNZtmd3AhKOimfwhz+UfZdte4L20m8kspOggp2PAFv
QatVtxeNgQsLx59rc5/QDq3svedoTHx/mfx+umwe0DVY87P19OxCkjoSPr+omvn0C3E/DjMZqZ+/
dVSB9heXpmkzc5qIvFTiwfK1jLpTTaiq6ESA8GmR2JSa576rtGW7UnjJjkU7neZqNEtBkZH74ha2
zJoLYQYUvega/C85W4Z473d9RXj1ZKOWRbw7kb2o1LGGHKLlK0ygvH86KRN08UQkIW0GSccsD/xh
8ElF5lQdWKXwF7d1VadSjZZ4VdwZiCrNCVlp+3K+V0H+1d/xASFwFmPKGVwXTn6/jwv+64Rfo+N0
gAYZIyGmGz9iXxyBtdyzbsI/yvUdd/ufgm7OMYCUQQf2fASNkJeeUSe1IEQMAAqbi2K03IWXRfvl
wQR7DpBrGavCkaadfUb+vPhpr1XHMa0JoZXLZLcd4Ot46DZf1IVuV4A3w6GrHknkUXZp9CbukWlh
ngrop8M8M8VUjEhCLlEgfBYSiS+HZEXLEDKsO8m72whWxics22BgZatDTC2lEc2E1vQbXvUUzpFO
uDvWQfVUxjephqJKll1KWdqhnhta89rsAF4kMT4bhZWsDBZ0RgbHkkUN8RRuD4fTSNQTUx0TVveR
CMOhE+EwbgrRntdI8i1zKUu/PraiGFo7D9VkFUctxVz/3YNWGD0QyRRyFH0wKSsPLKhYXP8fS6IW
M0GF1HVY7NJmjW6fJ+VEfEpnIw0NweXUBxiHxin0lSWAvXspBh5xCZnq9Bwliw45SbgwPMOz6ESy
GMKjYWxsEV7Y0xOFlP2tYg2RnnWuCQ/lxO2TrMdfCsYltXetfwd47nNKvimNMYxsmXPTzbzcEiE1
slTKWi1Q2CfFrIQq/QFZ3Ml6n0U8jKw1wYffrWaoQbWDfp5IB7IUvJBpB9cUd3PVK1Q21KWdKgfr
ZiVaQrCFDaXwCP6UNO1nMomc6I3Tcc2phSJfmyvXFG66aIxz8W7V/vR6ETASLuzX2q3ZjwZuoO/y
4tuq2I//4ofXC3k1JkCmRW0w+o88OqDJSiYbBOrdhDmzuBldMClUa1AMiFgAyzFi8RUYJsM7jeWr
Xgew1a90O8jmWt1pPNzsJknqA0EG8KQXBL4uR7bq5EdpYYXAp/yoAQB+BUUlGe5vxmJOzLFLl/5e
PKAq8GeQDBZDgYlEvFAAO8E0+eOD/uQOynR6plM4nHAopbz5x+F3qpZK9LTGRvg9idUvusxwfl+n
wGVc9HIjVODQ+9Amo1g7S1JcMMWBiOda+PTEblHdF+aaWFp4KIlsZ08JbALrGjZf4A1+maHC/1jO
f8JCodk9ChkS91u7ZIEuceFpPTLSdO8VR7LDQvqz4/sN0zACREsCJ1FOw+7RcdLeblGY7ReMrLNe
i1ZpqHzRNCOFFW2mKZiWs1bOMfaxGv8EBTkuor15n9gSA2LYQZPGam7OyyZGiASJ3J1uRsKBrOsx
LO5NOZo+mLDJYxqiDCJiDjPBg7XQ6FdNFs0j/XZLuUAKT0KLirDfsphWZ6rg8RRxhULNJf8IpBku
i31CMjG8tBBc/Dipwab7ERcMKR93u24HrfYUP2ofC5cemr43Y8nut5ssnR+QX7Gw0FgkEQq/KBT1
Kx0B7UCc0dajKoI4BD10sALV6Xua26e3jSy2oOmVu7iyecPT//s/gDPmvlGhThu26CuoRuMrtzFi
gLpKSW70FjFBTy9tU7iGJalHwaklpV2G+jRNsfD0cDKO0FVApfzY4IltPdLSPTtzcRmFar7CPtXn
zZQUW9XjOJ+h0csQxCx1jq+c0bRTszJFB6Ck8KCNiocMgnZv9sDTq2509U+lUdPYU+3hOoVvLVqh
7/dGY1/bR9kE6Kj03Di7tM07FkypQ35ehpMNOZrNyUF7AhQocyVB+Ms3KOVXg9tTYK71zXwnDJ7h
q6DwlBAPllVEq+/RRLWltWbmhvow6se4nqib3VBl1PeB0bnyN9WKLwfGIb6TMtWJ4+6aYZbMg5+2
PVbMnHrkKIlilkZRRjEP+WrG0Tym7p7YxKtEQIRRXrD22s+ImgRVbRKff8CUVlrhrwJ+3eH+mQq8
Cdd52TVjeVNK5UCIncYKsSxtvZ3BBDnFXUXtSVJQDcQVVr7nfxbcG7U0yGps0eewOoHyJICK2+6E
DcEHbVdmyGtbfw9dVnur3hPlfmlSm67TDecZgPnB1GUqHc7b0n8FCE0WC1NwsYds1rm1WsMatZ2G
ed1r9Q0UOjPw2wKeevq9cyhgofRQXz/+6J9BZjwBDegoeiVpvwWMFvBtiTyE6SFa2vDassd8pZs5
hSLzHYS6GgKOpCI/8scw3hU8sHMWhUTnMzZ1E+WC7lYNRQLhxTrgc8EPSlmoDWTTRS7vqwN7Z+EC
tK24bG08eqxkg9UONMjgpxRyLsVTmQVhoNjheOGpqwRAqwlVNVcGByBJ6HKL1DDa7/N52kxtnyjb
EBA/M2VayH94Vdu+Z7zHPV/AQJcB7AbXH0zG54kDSYN1KTZ7w4+PyV9MyOrdih5PIctjWAr+/h7h
rFYwm3VTSjwEpNCr8/fCT4PQM9ZC7urQXHE7uL4pX1sJGLmaQ1vETQa0ubXiu/v2xysbglsyddux
nNcXWOU4VGyuVwy5iNiK0dBZtK8Ns7ilLaud2dUdMGnUhlNQkv5EtzDC4Kmm46VsoNnR6CZVZl1/
VrzMIsV2wVCDyDRbzh+tXovyrISRr3bVgM7oI/5k7SRoFtQkuTpgZGr5rkLJOE850xdvekDq0KM9
wsmmYMWN525imKb5ao2XM0NH0ZCt2a3pbaDYWye5xU/z/rXsVSVFZqWplNXaDhZbYqL4dQowVnaJ
0KVwNxUmFL6BIFPMuynqxWRsnVPWdO2o098NzHtsc/dK+d9MS5fowl4PvhjaTKXR2epWRCMtJ2cs
lS45OISygX6hA8XSEp1+FIjxdjq1OeiT/q/ifej9fH0PAjN8OCeht/ftKQx+H4Py0W+L5Gp2j/50
6HUehpLAaD2PNMZwx4F9kGpkr0HpYIj1skaJGSFbYV2HgW0WSYD0u0os4kRbLaVUIWHvKR/adjgc
HyBOfWSk0n/DxHlfR2GmHZ37BWC43s45V4r6PUYeu9Ac3IXPrOPWyBxmyE1+dSyHqSxcMiP+YeuH
0NhQhDQM6IFpqtcs9m8g1hMrRV8Rd4Y3hDS55oiiHeVVFGna/fTXRZIxMWMX0npstj6EQ2zIDoDO
d/zca8+agJgfZ/R0OePK2rvotoEHL4KrHsH/pKBEkhxiIc9GDnKVq9MLZ0XV4px+aLBBlBh1c+uB
5PVJxTTyQKZwzRyfIq3NNoBsOJCGm8jhCCHD29OPuyjKSt38desvyu/FPBexnoNWxT6XbQrzx299
XYPHQPWSwR4CDE6TfscpY/yYnElphNCZZDFvZ5OQxPBNrmIY1k2lfxkbOyPb4d9r9BeRKpoxFaqk
IHJUHS+QrotHPxOLtRH5L4j3rnlQ8DOzOI0HiWiKlBC/inMArboUPCUleuq+41gReOuvVKks/Y06
GUMkCHdsZHwiGyjllabcIgKXFxXAYQYB6EUQz1X8q8Z6NmNsQci36VcljS0tgLhot0qAgQpPTn1I
kCdPqWdWqOuFYt4Uk7sdhsnBQZEwDqyscvXqaEAtnFPCgVSPd2S0Fi0FCHkd4yYL2ImZVkHsm+Qz
PtMqIZHhdPQnRkYbZCIwSlP35q9qWoNd5lldgO8SAqvy4qKLAuE8/KF0F33tskqxdl8S8UqTMtp0
l7v3Rvg87gOu7VCGdHZ76GzLlCQabvctcJeq/fPPQD1XyeRLs1QHoAHaSI3BYYs6t5yjINtnStQS
4b7Er/0hL3yXen4DDFkgvBKBwf9hj+HHc8AZUL6Byq7ZMjvgb+GUZnPvtxZHPun6jerCyAuRlVtN
ffJcD6GbgdZqX2MJVKPN+qZ8nk3cv/clgreEDWKEVS7nRv8a8/xGVrG9fZV2T6W5BOjzdsHLropZ
u8/nWE8frhpB9S2uOlZyIDp1MoboKE1LGinAg1A7PDlwNMsv1fohdZQhlcp63e7fcIbNZzOtbKL4
lB9HUuJMMWLytUHUpeGVbIoJUoFGWs/n/qjRrpQhtoXBU5C0L4z/fhlUE/4YCYSCWcA1ue3p4Gr6
UtRs0z6E4AgDPL25SYjkJVbqPqZhoUEK82O/N8Fym75NtJjzgVI5V5JVSdNCUrm5UIgkOYF6C+20
b48t+uVx8llawZgNy4b7pqnVOebtRGbu5x44ICNUj89ctS1PHcwIHGS4QsNnIKIUbYraHUoCfLKj
DSJzl93Cw86Q1HDMpLHRLuvC954+GlJ6QZclOUMs0HfGxSszLni0iuSaNot3wYFpt9QFM9rG6Yw7
lTblqCQtZqa83u/b1P0uRpAqc8gELPHh7R2fxzoRejbklMvR4rACWWjiWUkbmTZYp3KP4foOQoqR
Dxv6o08TkDQ4pDG0tmMHbjoaOGrvNpBuqaMYQo8ru6HSrUyICnQQ+vNyIVAtbr4Sp81hMOHlwtjQ
4SI2tiGna+JtO36otp0HjV+xofuUoABzRGJJiQ0ks9lcwXYaDWdJWSu3eLRDzoYEx6LRyOqMZVhf
V708SR1iR4NWYp7tRqyv8XF4dCteP9XGX1CQT85fgFxmKUParjPbdXe0tkSIG6caDJYzx/7Mk5wm
AVpnnXkA7W/YoQZBT8eecthKpmUIItflENluLl/axwdbaO8V9o3ErQReqA3vA11qQGRNRrSTIP8v
XepVhmSzOUdPy9MxLWtI6epEkwNSBp9q9fjQfuFbhEnIYLxDIrydrxXz7j5sCvMVI6PDyDuiR+Mx
Kl+ZuMzEuj89ksXtxVx7/64rDLO9VSgva42KVFDfuzR/mqhLWJ766jhodzEcFUDB12c/cO1/j+sy
EddmsaWauG6yMh+Lm6KWM3feiNTdPXluxybRh4C6ckyA0Xst449SNVI91tam9o7FYoHI+gL8IRe0
97yeUtJv4eonxM+wexKqjxYhFNIuTPQP6iyvsuTidb2GXwOlOeFOIfQnKnnJQQ+FhPNwJHpxGq4r
A4O6f90WLNeQBrhz3n96GVgLZcP65wC2adHVu454W+9Vzg8HqzGd0FOQvNuyayvO3TiJL5ngCofI
SEH9uOFOUj1rHUXcTKIlnepalHqNfE7g7yXliBTW3W3pTHz2XYFmH8/IfoBpZhjSWhqXDOUULpGJ
+zYwP7YGjAlj/9Ma3G09a1t7uwM2214ksDxg30jDR730AofYdvLPM90pNsRXbI7ksKEIQN70mWZp
YgyOqsDl2vfvgTZCkB8n5lTtU5n7iP+qw3RXq+irTYPCydPhrIICXMCKyrBBM+S82TnfUFafxNu+
462KbiH1SP/iLHIvsAW3AGFLF6O/xeUxhIf5uiiJWmqfJz3qxu4cri0VgtQx/fzMrg7ZxJLqD/Er
VKHdYsZh5YYzhlY1IsWbPlrLo0EYowWWjKTlMvZTJWDcHPAoQici5ut+rTkYl7tAI0AnsWwBDgXv
oZSdvpoAUuZRYPMEan8RFQPxB9Rmsy/eRAZr0gZtEnNwskd6cPbBM48JOeRPu3IUq0pXBdj5wxXN
fTACxWN0NTbZuEPvNbeATZx+lrZfvYXG8jGK0IXcVjDJC60aLoUAo1wxn1wlq/MbCPeuZRAItygp
UNFMbO3yiXu8HtWQtV2u301RVXa8KytkpEmOfaSgstDkdw/b5+LDcOmwQ7g2B3V+PgcFBytbNQji
tpsy74wGTEexIDCsoYGOOY4LVt/2sB8vHtS0rCnFI2VFpKoKD0imm7Hb3HnvqBzK5N1mLr0HrnwG
vZDbSrQe0tZrruzFdsLexLimn25o6MXG3zvj8ab7CGjzo9SCnj2T9vwR6UhupLLQTTHIRHoWuwqL
jDNLxj19zyG+4/4D5IVz2rTIbdEP4dJDBCN9nG7lAjuVBkrf6mQTkG3ynG31qOTOMdbYbRjAd05r
q2mx1PYPBxW0onU/5vNIuKvBqTqY+2a4cs4QX2XSq/exiNiamDfoDktDC0QC4oiCdz0lcyeizc5z
n84ZWcNxFp96z6rlZHX2OP+1IEld9x3DBo2WWICbs3UeOy3YWbXTZMpw8AZ63KLTOZoBb4iCRyTe
v8HR7MZlFsQBil8ew3kLHskLyiHoGpltRPBMB5Tr4E7vsl7zX3NCyI8tCG33CuzDDiVJD3EHcBi9
mM3Lf7POH70T/nEwHkBXKB3QdeBU24OVLNCJkDqDY6fPcbMD4g9LCbA/8S3GOpQDbEWF4UUMVewF
8Sab7DUrNNRx9Ch4Fd/x0VaccOBa7f8ET1o4H9MT/Rq9ZmUpKQiftSRwAGPVbWa7+qttzhGQJidJ
UOgxeFv3iaqZf5CJZ3pPSYL6iqgQerDDxTlbC5ly2kMQCYuyWJRce2So5VYDHHNqy8/mWfy1erN/
RFocMsgg3htYLaQg4MujfFQMXeJQQ6E1c3LL67BxjWsibDcGfiCzws9gD6Cn33h15BiO1W1yuVVe
8n7fIn1cIHSCoJHOjFdoJ6lVYgQ1Wl4c4e4NSrzMm5YiEkvKzdA4KycIXUQSyOZ9Ud5Kr2XSTei8
b9u6WD6X0zgYYwXue50ldCATsOkP/tqD98zdi1jYBCrA9ECH+24NYJiKyeffyHps6Bvm9iUV77cq
ZebtAIBbocju1JQ4rg5ti4RIH1NhV1Zpcm3B6TuHnhAQ0bIbxDiMDY6RUvOZHrLCTR0j2Z38KIp4
7BYcbkb1EEwaeQNygIEAmq1IvoyQe+tdq12vDHJoOHG1VHY6yH1zfPYIMX1KbRExg63sQca1OzCI
f4DcsUlOJNFuGGMw7WEryZm9RNxpK51IBz+Q4LoMyX6dHGQ8tA9GLZf9yuiZjYDxckjFmz1RJfdU
tExG0cWmMkZsgw0B5vVYyLuDDV3eEGa/PxlkMsHhifobGoSQcMM9mZgwUqO00vBdJspW4j3FSqyl
jevdybs6Vmf545PVZ3rMPrgMxc6Tv1KTyfElw+/RcrLcNJshziThMX9MKgRF9/O1vwIfIoAIFKZX
gUsAukLErSFeYiPSwPB8HBcYaIVv/u0BjeHU8AaDWbyZPEIzVh3fcWNRAuhRxc1jp654GaCA1nQU
wj8Y4E3QhzM7o4UffwUWED5ZyPj0UCunBH0pIR/IDWIcxO51JSjb0n7/l2vN40pxeKgxD4Fiw17R
MtgN4+RLMAfzftGl7yVl0RRFcoYHQeiu0dCP8TBVJwjl6e3IhZC5KTiF8WutVhSf+mGsoz2JZaja
RjwfoiqzaGJaSIfgj//zl+Dws6b8E3ut44ZlRcnX0g59k7pMAuNgfR0vmiYBxK7P51LHCQ+kxPH6
6RP0PUI6eEjRJW8P70PZwR2s7ZrmwbV5pLDyFdniedYpmNKTuvcx91my7t+Y3fUp9GihgAe+JpX4
TkdgmLdspcCNIiTVAgvk2eC+1Y3TWms9mbJsNrCZw0fv1BF2tfc0F7GkM0RHV2mT35ioIcQbirV1
IOgb5YRQKOZDE47bSUEHgNNUImU6yuKMxcSLzGjh7Jkt7Vw7dwS/of5mvlXHlVOVrahcaRBtI6vD
3vkcOEE+HdWotti7Q7G5tJlNWvzdrpbcIXjZRO8Hc5WlnQrd1KFR0+BSkJtxXh20giaOM4TNMvkY
MXZ78TRnQO22eKPtf5IqFWEhuTsluuq1RlXOzfeMzNALVK9cg6+0UFsO+VRmL8MGsAxswP+ekN6M
gGEU9qcBC9etHewddJjOTD36NAP/tOpQ5Qw388cVg0HR6EnVP3youWI49rFV7J8GDEl3JXkvEc+b
+uiuM38Is5eqqZ1yRVyraTT9Te2gjGQBzLfvbIDeVlow0YZD2tplVamgsf/y5AjEAcSw+rdURp1a
TU3Igre1C+ACfz4XCiKf3hqtrgXJjJHVcsfQ5jfsSkzeCWQo00Yt3q9qmBOE1RorxSUCA+c2MxVI
rUhbQessz8rqdCNvkWJlHOp8Gellw59AKFOPyIRJRB9IXKOuZzCQu1+sdaF8Imk1IyyrihELBOuz
xNGUECFZVqPCSy10qoEscz0zI8RyLOPcMN3X3sDj+/v7ZrXM3i7fECtrBPiqeZJuaCk8KKuxJ7Od
zNMpuextSiViZJM2IlHNRgpbmfGQowxjvNlRjiHnglg5pjhp1kQrFj64EbfooJI3t7/3PQg2sUiF
WEhgd34lbvAegpsRXiVmxMiJ/tyn3WEWzCmdwtWZnvMmLBEj4G4yYLXjtXXKtTRoapONXHTJyQYC
NgPNGdPUpo7YHh1oRsKCrL3OfRZGlhdKoZyCk18faDVKTsW4XUuQa/i49qBdX4UrmR/zl7TJg2p/
GjrZyNWGJFvkbE3b9JmFmXM0lM35q/e1Ss1iHlwC/omh4pFIU7Z+WoaHDgvv2s2JZDlyezHa768W
gpbtMzgOA3fgtSPaPXprSHhLmh7ymQwRUBhv+Rp6ML7NlT9tGQv1SZ6E47GIh76dP0fUXH7qtZvq
3GoflWeD19VWZGFPAqgDmqvonU8ENRCTRORRdyxoAJ+R9mEd2S63MOSMMDcgvrZRCh+dkZxCJtsm
bLj+ictTgicRPM7xup6O4Vs4vxVgPn7HB6cVFKP1ZS8QoTit/qMIHGDJADVcaOSQTNu7uoeOqhIM
49yhwizaRBQbsG7lm33Wp2dfC5AXrkv/9xKGc1iem4hRyXbvhcwilzbBiONeUT5QJ+RvdPerhxNq
7QOEWOwF7tZKDLCcoadWsjd2V5XsHennEf8y395ZOF4y+KDTUyeqoV/siulgbsd5GibTMnAo8ZUC
ZhcEDBafpFGa5MqsDuNqYYwQLX6OarEH3ZcjTjPFlu4cmN2hSTX1J02UGzgKEfcy/dX8OlMMcko9
9xNbJive4jCWanWsIzJ1eB5WOBGR2SHd6x29iCebMp7vOXWNEqxsPSwGYyrGUr1QroCEeHarxPKD
K6WLK9K3rwHNPQZs4u+2FC1nRXzX0tqJfVaBcGaOgQ0a2IvsYtAvT7VgW/7UxhY/g2RZGamQWxWA
hXszcdCuefbIzpwY6LedPLeCla4TA22buXzC3nTgIdREwzBpkZLsufendIKmIc0ryETsermWHq8I
F6qiNRDXDyDRk++oB2rAJWU2TM9wIsVzIIk6/A9wGA9vbBsOvBcJt4T4fHyB3tm7kuXbBTGBdTun
5MNuVRRvQl6O7SpFBkYD9j7xvSqhTXW1yjZ/He4FOWKBVdUiLUAr7DsKFB11iLy16ZHD5OHNOB4Z
DcGa4WTKDQ5Rw0SNNqe/cpVrxViiKqN5ExesgF9dc32Tz9b6USsmq8r2g8IyasP4s/y5Z7RMqFYU
wy5XGBEuHVEW654P1SBMBBlEK/P+MbFZxsy4YT3D02jXXR4Jv3OPsH12fj4ngaIiCmfOsIbKsq79
SQdxxfCSUBdZ0u/sl1TXwxixx0zL++4HrpVpUSWAQ0VcVaPLYJXK1uUGDrA7r7ptkr1bSoERalJL
ZcqkZ3IDMGD0FIR28GaUWuPnW55j+2oy0LnhGZyQRzryIaxJgq/Rt2p9rpp1xWFbSQFbVWcdsH27
OZMap0RzGiKZmLWUKCThGM95XiKU0GbbImbScJPZcJ6pmESrLHseMQ23eGDYuomEvKSHodXBGxKH
XXicGWrOkPnDY07o3gLFYoOsdjTurE2c7T1Wrg/dwHmDR6Zxp+th1YC7o7PoEzcuRkE4MDaQ1ThE
+PZAyDg/xTe/y0FGHmmdE8ZZax5sE8EgD9Q8TCHJLI8qRaEkSvUNBNQkju2WNMiAjV2FnOtv0jLT
qvFCXWmp91AgHj+5LBmNqPTQI8Bllyc9CDQOFOUJ3MKf/lm4UqCU9Mp3+PB6GBGzEuA4ghgCQf0U
aACS8x0HKflEVNN1ZQs7hbk1FUKcTD+Olg4/iUFMyDG2lZ8H7SRGRDlc9r4U4ZonUzqox3rlxZJT
qGnwzHrrTEOFKa6iLcGl/+giDbCTSbv8obn5Wz3W6iNbPXO4Nig9iB5FqRg7Iu6GqVPdKdrwTq45
ZWqbPAmfNVN1jKd81PjfsnU5myGNAfz6r6rqt1nkl2gz9wEpT+2ShUe97rhz3KyF9svaYtezk6FC
hiexdpFEhZV8sZdueBkCb2Bz8o/sCNVHe4f7sNpf7wFjQTC5Oj+ny7raHEri8svZjAfpLGnLKVYq
O35cz3YfF7hCeX6Gcqb2nY0EW7gDU1m9wYIghcMOvQgrTLZMFhKN9VjmKcKOXwec9jS4gHiVJEb+
0T//XMNegFeLIKX1VlFdAn94169tlKsLxGa39QmdFA1VSSps75CutpgcOWlZ4dFFwnbMihYgfl73
unz+K+1SKq83+1jdG/NmDeJ+uUak45whIYe6YZGWhRCt6O6MNOeCg1aEf1BpPul2tR4m3sOZX32b
I8KaFVNsLL6HurnoTosqH5s8r7A0RN09Ig/8nP8InIVs3o7zM70dfv6Yb6PysO9Y9GqJWSjusZKD
ge/KGAqe+U575SvnFVVecUqTN4b2GdFdSn6rPrleHK1CecfRyvd0kM71/TuIfBJBk7dCLkLxtN0I
Sqw0jkskt8mGH8+aeea56jm7tzdF3NSBU0OCq92fmMBZJKCg3qAMZwRTpq2UmJFnx5DGibQ6VgCm
3XasB/ak64SbYsR7Kqix2fFjXWkbRg3TL2kyTIQV9tW5ZnN7ubD1N/8p5YUPZXSI0EAuDo7xpwTf
HevG1b1irjGf4WX4n5eWli+4ysWnmYhAdbf0LImzsWmXexsd0UH3rqH1pmMcDyvH5QFqFyAD0/JK
CpxfOaGCk9TtqJGP9U5x1VU/8wEk1Vz0pmvURbipSowr+CR1W6GcTuhAi99KohtETDpHEsECzTpW
sgmJZ0a4iT4EyLL6SIFkJCz4Bk1X37qsfTVMBVM7XpLI0zUdpNejV9Qa9rgXrEMwQ0jyiuEYq1W8
sqIB/GPJ8FAZTZ1VNm7ywprL6+WkzR1MMWfPfawvX/H3fj2GU7kj2RAe0zsTyAvT0pUOEkIDQLl3
JudERdl2zt5GLNpLseVdcczG3go98aRBfwUWSEtJiNFnIwqaQzR3H1GFQnBgAFrHljHOLa766y0u
dL9xoOUx2Tz3kQ26Pa1n0V2xZ3Ta305VECbj7Ju+s4vM8KyypxL8k8urnsibAngoSn4hV5FP1zW9
wkKUiDAvUiyhm2RSynhvWTwG2Eobt7PED2hB599oEUhHyxqFetsWfIgEmpjSiDxycholX3yfUI2w
vp6lSiJng9EZY5Uz6mgFe/BjIEFm+gew+8AXzmrHgk6ApqUBk6GLgaTeS+SSahYqlXBhUbQn/FF+
t9heGZPHGKVtgEwEsRIeBDc6yKb56SQr0gnEG8TUvMH1+ZGo26dj1KkfG1YjEqYkQzg2S/ixAhK+
oJSTEYYafv6ZsJRfONqslL8fOjPzu1Xo7q/OUJ+OqNVbgLNptCZSrwYB9a/jcdqVubkzqTcW35M5
J3jVw5CE3UUyg9w5CSqOEnFddC2NRYfFV+BCvuoBxKWfyZZLgDWgbxjutQ/kpVxczLBTIabCDdbr
mlllCP1UUnlTd9dMzK074hiNl5HB4coirlqL/Enl2dCE7UuY0k5ACspHXR0NfsHZzHOPTghpoAth
3tlUxa0q8a1P3vXk9Sdidw2xmCBCdqD2PQEwwgcnk9tcqMsUOIonlsoHLYNZObB9Lq2HOQ/Kltmq
VvIurftmf9ymXMAfzg6DO6P7EC1iSP3+fEgSyMOCG8mWPg9V8XMg2rRUxHnz2S4STZ0JpwXofkvd
cocTj4XAAl2PG5Yn/pZF8nXBzch0tfw+NSALvw7d9ZFSydiiH8L7KWzHjRj+Aon4FWLGfjJYo6vn
pl364qFGkWEsT1AAYJCZOiSijFNuKmeNtO/ckzFKa9Dks+yQFqA++tjpGIdi53b4PFI16qs8CT7s
/6whS9vmN53+Jdy7xwwullBVzvIo/tKg5UliQUs99MaLcs8wK7rqT6bCNO2p2qjrXStC2LneU01Q
wdxf/mdFUoPLY14V0ZXWe85CfXcpP94GyNeKdYglyIOncXplzTMRSS1V7LyK/E4JmQv8hKp/DIF4
lECX5rYMC2WHh9tPuw7XjR+Fmm/bAIsdCnd9zBYu8NEwa0CI1E4dfeTplgfUa9/1Du4oN/TM+ZGN
vI7GZh8H49Tc+x8DWsuv1X8WstQjvSjFuyCNw2HfXDyWRyguxM0OddMUYb/v5UcoLBn2zB1Y12Fq
Av0KRk8dqagjIl4v8p5NTiGxbC7aN/vTC3d2NlVXF+NfqhMd1EIzcSSe7X3L/7WJbkkUcXvedwae
hgqF1cKULfLx8UAelJzsTglj6nmu6l5LfL3vJToYp5mVIVV9NkYwZ74n+tG64AI7ZVJlTi2tSqZs
3EtJoGZvvUWnHJRbJujHe82oVoqtYvs+DEAmW4vR2AwvRKeb212P1q4bN298otc7h2rqFSNNYft1
4uViE4tE0hfjcPbKlD1qUVXMf8jUpYUzya5EAtuXT39NkutiJn5SusJXoNWV0rlJzQoKuCbsleU6
RYpaeUKdwEQgMTZ9vjyLBz5Z7qA/Bmjw0mDPbEwFF78DUPXciOL/eTpZFBihf4NolrxDxecUyS2I
qNNbOyThxoYz7j4K+/oG7qIrcgiIRoR2lpIO4fyg3CUuK9SsSSN5VeTOvbQ1w1X/GFeTUhGkrsrG
pIE+MUL5/jUirmLk/GJ3J90q3ja3WX79VSNGtuSds2q6Mj9CYXQhElcAp1OarIFPgeDybwF7M7sA
AdanpfNQXNFGtjxNxyzPhbxGNvV9LAOM+ylAz+sHMhd0MOJNk1uqUhPhSSR/h++xW1It9v1h59Lk
clS2ALCzLdilhBX6EDCFkIGCOfDOt8XY2qgxr+gSbM66fvdeT2CzFqOaaW3dRA/0dCpizUuBSoNj
0oO+4Yrmo4JL0mzlnz7xn6kMWQALhUjtEu5tORU3mcTKbUL8+YLC897GXERMbAOmLGgDJwhar9b+
WOOGsP3nju2KwpEg4DCrzcpGU+AtnmlLSwksbAkXE9JBVGpp/Yeg8d0qXleMvDSTRp692Kqtwfyy
Yn4jyxcV2UrNxyRPNV7UBppKmPnHQlPaYeu9bnjcskfbsxt3Sg/2lS29R5ewZJ0jCR3m/03MzZ2A
t7Dq+C9Nt+c5NBqR71LFY7u/i21iZOwxXaMubVTlWGVRg6Sxza3FVWZVWzvPZvbfM0VwO1lgoseo
cL9+Xc9fMOTxc66DmiJTBGp2fGxSCkDh77deBqmV3MYjb7eMdFOHHsMeuZfQ8E0YuEeijXXViFxy
YkCpuwPQ8zNhoKDO9sCg5gSbcUmMlVqmnTBpg/Zplj5FVUZZMwYXnmOaU6ERaIy/G3ShLXi2pLq3
6dFoTtYs5QAnjBeqSfdkxeovZkVWgxUyENoCSpZO8r+DLiyq5pEkRnOaDMeJQbfIyiedzddzY5m5
EQxfi8C1jQ2/wvpWag1ENQzeCQ6h0G2P5Db6b14e7q6fEBpjYbsoaHeIusmROqkYYcBF/8CP7HXi
1Iey6k6Bf2rWoCaG7xg0EKI0ipMlNP0wi2U7EoeGqeKpMsrv4cbFVMGVdNE/6kh+wqR9BvaUUTZx
FKJYPA18ADxyAIcpei1rI98s+rf+JlJAyfcVTDKeq67wm4zli7y9LX4+z9maMOFujMK/TOZRj5Pa
TjT8oAMhAP2fjfiGBXJIYIChONNMTU76vplb3pmjIoEoBTIa89Mcowz7C1SEIkg0WxcSU6Vkj/f3
3NRblL/GUwL0/VDwC5JJcO6pYYQlXe73tn23+xTD1RNj3GKtznpmeXMPRCTnOhTaioVsRIMQ3SwO
F5+/AldlM81ai7u/HIVKqskcy/v+22lMiw6t8gfu1Unyjrm/LldcHsMAJvJ6MTV70FnXe8yXWNJm
WkXj/1iiFNmlHfIyiHzSB8ARi4cD00xpaC2B3LcRj2Sovk7r3aDaXpbT/CyDVpqPAdbFVAUFCL4b
tW4Z0nvighA7JVbgCEsfzbhOWI6VRXi0ed8jc+JNsEDVT7KvqIFNl+OazlFSOaHIwBdrlB5EGS3X
mXruo3pLAix5aeAhu+xGo2jHmcp6MS0uQ61CN2z3FGUIBSnms7UONhirzPF0tH+8r8kD9e52ueEi
6vFcubna3rH5lla2vC8sd96222rTzWFtIDd6RJ6PONyXXlBs611aYDFThaOn8A+qbULbUoOP8KvX
W3yYMCHBRMot3y6e/l5de4gRHvipd8DEtqfx0LBIkNsqjFIW6wt9U1qcckH/xMqkLZxAYFQOGOE3
Nnv5kGu0yBrIKXZt5ZTF1H4Dw1jDK9eI0/j95kg4x2RGYiNCFkzxw6mUH/IpzveGrcZfG36PglXC
hIrkLuLu92FzyQzBgVuDtPohf4ilQf11niou8hvhvdINafEwRzaR/XzexsFyJhYH1gwQirnBAL2Z
W0BN3Oi/MSPWq1SRx3qrHHxhBvosrUVVy6ucj9WSepD2vDm6O+Au1sii/dUmMvGXYPUBdGn3+iH4
3vRabT7Yi2+rUSVWxAPU5eAXo6/gIb3VepWvnb2SAOrWBE7R7nEjJvqhiVnk8+/QyUPbzWXbI51p
XSijM044JfQhQQm9jvVhS+j5oArMcOvINSvbB4WBqe71UueYtAnylpfaLvHbZVTy3NRZsku2q/Vr
2HvY04/gix5Vek8mMgWSh0BJ6zzkFR9ZJNUWnLbBoqh3QhVJFKyV3+Y4XV1idt02PZvngEYOuHSL
WK3SYy9ROK3ok+Hp3bZCrUXGbgxPY72lG8pbTmwUi/Go9GkdFmBg3Vr4O4iwf/Gmk7qbCzLEJIoz
d4cKV8PqLDCk0bh4nUyEg13g9V/qN60jtJrVA5pmb4rSnCghoaYjWFJGBc38lFPuCnyhUIXdp0zo
jJgG1X5Z9rhK9uh+/2g4uLBZ6Ep3k4CZ7BAa+zjihG06BP61p2BEJ55l1lz/GIDQK4nHEka0mJ5Z
InWaH8oNYJgAaE8iHMwoqQpMEQFsiM+HCGEWQ60X4F8+0pX0qUw87EirAvhLWok6Mx6+3EETehG7
uc4dkkhBfViql8k81BrH79G31IX94sBp/vtBo8nyGEsVkMV2atUh9Z4wp/LNSvfu+T71OYcmQWwx
aUrnAKTdUNEm50ELBMkqhFm1jnbCpowj0MVX+qe5P9FpWYwHdGYCcLFv/zXK15YdvNuvV0Kmlm4I
RSwmYjBm4zs6gGZQHFvhkt7dg6sZV/derA+XBHZHD67knfRQDlQgKS7qbT66VnBBl70mxkwFciRM
2lxRX2nGsjjBCMT4DmXdI10WCc17ganLrOWGlS4Joy1+sNuWMTDlzUMxV+BHASHa7z8SfcF9W5zf
8nkHe2hLbtUdfiEjjMoLiMA3b3rwdRjiSYDpwj96kjcTnQNT2ydoVkbgLfv/X4z1hBszy3Nr5Vdx
voKB3gCavbrkdila6PzVgR//AapK0Iy0FIK/ivuLpQTHhtyc3C1XfYkwFn1+VO8FI56habDBs9v6
rVfSiyQPefyijReIMzYu1b8YUwBnUBndBh6yu1AKojZ+x8Y77yjJwDyRlH3K9YXrek+PxIBYJfJA
Zux1Xm1w3T313un7gGV1IGBA4gLJez0Sk0otEFISDVTp72BknxpVwbVyR+yEERmTBEX+jcfBE46n
IXmQEoLRLi5MCnisx8VdZ8Qbom4bSXQndGJ5p/A57t66f+GJYuvsu8FBGX4kVuhSQCiE3Emm+l+P
5d/hpEKzSCZcRdJlU/8yRFN7AdeTRTqtTFCRohXxUpvmowZGlcLQdqeMhZYG/mkliKE2xnsVVrQ/
Ax2VTetgk69SEt+sjLrKxr8ifsxTbsGKB/WQM7ZcQJgybpPZ28+0iERfOp/Lzh7/dtYdwPgCkYSc
qtxd6WRDEHGHEtq9CtI7dMqk9sYPp889O+sCJY+g2oc/cNBAz3tS8BYMHaGX0YIdegC0T5GaNYvO
arKvkOfN2FeAUhH+y6ZdYgrpSId8tTYaCf1u661OVGNlzXpIowdBFsYnZAVyBk5jRe1R0pWZfbZV
/+q+bDxtKP7oX8HTVZ2LfsKkbpPWV5GyLvXH75mP/odbAAHAhr+uIA7zgDv59VTLD0dgJfamEVFa
AR4Qa01PLvfCNb7k+kslynFhw1S//4gtAWmFOvn68LaEvqPOrIfsjiL7oZDI6U9M2ytwciX1Jfjr
ZmOY+FfiTn+lcCUGECtkSTExzeOhHJsHpjKaTtF9hO8kQfodj7wk29Yj60TD9lclHQSk8oZiQ9G0
2/2tIucnH+ACOP33GYIaNm1z2UlcYPRoa+VD6UGpkbNpvY5izlAbgfdQMUj6r3kRJkPj1eqj8/l+
z/W3LhUG4EpygMH7xQ1nOUfu4rtrrx7Vu+YTNsAetREjH5RtLBGym8r68kAM/rrRUdjiqCe5siHh
ABQcuhZenNCQk5woqsjwZ34ArPWYtGExTjBuB7z97ZiM1Jvj+EcfebQkW/kanFJeK2IgxGRkEc9k
vZguLZiPV0bfV5tK3ollXqw+vLExxqZnY9iriVGvrfdafR5qdbV9U5+xIIDiz5UrnwBo8/Nn29Ix
FmyFNSUJ7Y/0srL2tRhsCfJL2veJPMxpO8FPl9FGOcsivNS119k9DXtVKl7zf16qi8+AU8YJDD4U
eOX8jtDJ3rn0MKdfsO2WrQ5N/4WoU26Oy3nXE8mhzdHmg8Qlm+Gwvy3iVSPe0qzZ5tTD2Xk7boMG
MaQfswFE6tk/JYw4+MKYknAilFQQmaamS21TbDuI/KlcJ43eyVJHCchpLW9y3Z2TRwPVa+zJbq63
N7uRyWvoL+3ZsEjg3fMk2L5fhyCVYcBIaW8P5tF6lnVtZkxc9STln7hQQNlIfn0RsztIrvwDPPXT
9Vi4lE1c76rr7f66/a+KFs40yg8CSgyodnDYotxz7n8yHnzs+WWGznYAb6mw2LfRYpTuMUhqiS2k
YJ3uTBH7QMgXJ60OBN8TcnHtWE3R2nnTfBWKiMDIE+sh+pbhA4jzW+6XppQvMb8tqlOxzsgE2mut
SImqF2kIzx6HjFHRzokkrJX/aMHWSlCt6GQtlmKh8CYlfbGrxorYgFYWNewA3vrceksr3a8tLAuH
gCeKolNUnLkwoLCkQ9pqOYyZD0ZcwJ8gZeIzLsviuJnSvBfvhGreA50o9+7VRzBtHrENvgi/vcnq
8bfXYd5P0gF9Zdy/elV07ou1Qy+CZ5g81FD97cKnf73AG7xscJeiDVFdTCMKAioECwDJccgwRLsg
dhYehCWOEJAnRxenkkYwYOQPTIOiMuzXOOLulgn3a1kyD1GewE3TuTEzAlw/JODMEvpyp8QHWW8+
UrIClrVi2cvIS9W/DPvLeEEDvehD0mv4ZUW4kleSRhT3s1kGVEc8T1USmlumKmFX9Y5XseR0/NF7
GFBljbgq3NUWo5snPT8Z05vWznpQIKg3OC/uUK8jXD3+WCB4NpGYkrQL9qwXgxWMOqpwU8Ir08lZ
W9gko07LUUhOMvtRPQLk9yIg0ml8cBwCjgwZrTfhLuPU4JrpDrrJh8mrHnHjSigrzHBMq5sFjp7l
lop9iWNmzjreFngDCXLKcjHxgMFCC95N+UnEBlCS64AD9RgBO+wpq8AMS1oj470p2TzcNn2JQii/
BjvXf1CkbZE+vAv2xPhqU9E/PjW0wB0JchRtXij5NgYoiigyYC5cFhDgU+dDkCOuWomx98qvl2mY
3uQM033HRjSHc05n4L0UPZ+mlyGBoxedEOqqgM/RJMhdBZ9aWcsDF95bEmg+R1xc16L7sZHOiTjW
vmXcRZYxTxFC60JvY/PJSVklKSTs1C3RPsXt6BwEXikwmbsmcCFjfOYS6Ytg1T23ElySH0A3LiKN
udMFddX+C8WBpMW3jLghj3NsLcYqf3sRy1QanxEeYOi003p6igwEETguw6TNY8DRjosUUt0ru/ca
ZRC+BwPmMuZPTP6CRbwrqc349q71S/sIR1gDZYavou6ftA3BH5iYvQaNOeHCLcwwVOtfs8olIBsp
hRNK8qIof0nI9NwClsp1ojeaIbWMIuAb+/x3fRVPSHzbSTF4xteUPxtcm/uBgb2rcOahshX2WQ/j
6KbjaKGq4RvaY0FnHZ+aAuJtn3WQMkoxTHL/HTVfDJWlZlypgINpMWHdwlL0XyIJ7w2QgbxsBWUY
Wibs+uDicXEtVgDVLE75UVgxKbnkP7gwYHDuslIbwKVb5PLPq6Qq/3/8S5QCXg/CXBbXSaOteMd6
NYxQCoylw99gNPyOZjX6T5a1tX3DawR53iuOqR7qWgC7pUnbF91NDpY6OyWPAh9WSoqF6jZYDNIY
r6YBr3drsgpTbudet8w8K6Rj3OU1ffVvyxUimRiAQteio6lRYaOwKZ1oJCtnrSbVa82JgpWDOLx4
PkrECbnS/gDwGGfQj59F1xZTifusPa7lV0VfnPrOXPmjRKhHTqGU59k3wVWpO5n0xjLNioGk9yT3
7GgZLSwGxf6Rdo7E4qcwVa63s2bctPf429Yt5063i+Ta62BFtnMWKuKUZewZE1CV5iNlC9nLROMy
gZd67IT6pcT+gqwgP7dS5/kKSsue3DpiwaXsTumLYvAC0s4/BXS+r1xPNF/3BGnclKePjxw2mzUU
atdwALPf5jUUTaX/OKxKJkqqDZttrZJlrBYGZeXgSJimZGMnrCXmqHhsP4/G1vcqq/aYsHVJltYC
VMB1wDmmb35NzrZNaqXmxq0flF1wmYwjzr/b85hVs3uGnSexlMELYGmDGHgMk/o+YPfaHV6CYHBm
J3bKrCHsLkv1QSe8fKvLuUQ7ewBNofcE8Lc6bHskt8wSzflJyH082yPl0uBzHIoC0q4bdzFO7aCJ
qI7qLYyOCviHTQ3MW+OYqVnBWiBTwHlTRRyILGhsqdP4boj6MHIjHMO4Dlrsm/7vpReNaDuLWfqR
sw55MNepZhkIHp9CQ7h8F6dH6vmYAaVXCqoLkFlsPMcuDjqV+XPkGLkTSKiQkfdSW5oXrbiteeWo
T1nySeXdAJJDIA6xW0qQDFMTPRQlE/Nj5V2eFFE2qPUN5Wsk2y4CquBQ04WJCt8FnGJ/2QUtbmiO
cRMWRfu7eEo/A0jZ1PJvBGxThLNX5oYBKnteD+b7WMt3vVnQvf+OgHZk78aBHq1jYTzoZLsJRyz+
vQIpd0pw82lgS7fWy/JJh8x1e0LAJEESQlQppnhEHT51AV6M+RrhMNKaNnYRktcIUXHj2ufnF/l+
UqqkJwVWnMDtc4ln7HcJs454ZZw3puEtoVhZJ4b5WSg4ROB2HogMAnDpczcuQgxu7qHVqd3WnoeQ
UM5sGiTH0Ml3PoFPYG1Ud/vt8LJPbbANqn/nddUPoQogOHd/LxuxPgoeP8YN9xwlJM/Fzf0jG39v
BO7SRANr1nlv9BjEN6td4fciYygc/Iqcv9hjMHaa0LCvpqmC51byXv9qjuf8pw+b6IFf9Ulbv49j
f7hiYtSYnEe14R1rkEIfKviegZ1UYTs3TX5e46HRzz6+oLYIa0ZseIOrASQY33m9M/gTMOKvdxT4
T+s9VM8jpt9gyoJmLNkGjwBcA8dW+OB7HrWyta8DhPByPqYDjKBBFWoSH8eGJHkNmtigPoyfqu6s
5OO2hJTbpH/4TS8edINabaKC7m4dI8P7escWtzBQ3v11AF/K+mxwlvkiDOTi9kaRxkg4swxHX+Jo
Zn+7RmUj75Wr4Xp6dR2Ok7Q81DmWU8kbwIzotZtY/w8Npm8qLbUM1BjVH+gs5Cdaok9F/lyP0LT8
aEV+Dgu+ZlHjBvRIO6mNufmitmw5a+bP9Orh1PFsjYNmJRjMriMm/SCVMl/zaFHw583sN7BrSfFC
AZxHHShg55wAlxTozQ1qFq/H5r0ll2DbowAHTdwMowbr/z4P2NYt+syLAehE2jffV1aQg0Nk6O38
IEAsFe9fWuu325y7qBmUZiQcEFCuyNCwGaqHvp7nmLJ9OE8qDCM09BDwTDKqhOZKAfp+nzZ37z4B
MseZKL4d9we0bCVUs94IIGAnkq2zwPZQ7PK+tJehkeUmvxfvuMXAy5dJhK5bvJDwNrFC8QXLk3w8
5NAiuc3M+3MGqu0o/yBZTJ/EBDRSXlKwXp4e7aXsW97PoYfA6f8YfBrRoIzQEpBQjO5AlBQu9TFo
TD251OSkMBmd8HLXyFD/Cj2Gprv2vMCDhwJFgPa+///XUrkv9GaOleEudw+wVKGj5dNLBGoacs0G
tZRDhEdXgydxxLzt5N8OgP42USITxEabR8E47n7jgrKpDtmDUgxIkHmqIn6D0C5wDiGJPkDuOcQ8
kD6mQkd2F7pQW8wOZmjelLeuNILrekD283OzRrPA8nHB5gfRr5NVQeYUJEzpABvYKkGP3rN85BOj
LlGoqgzuoJuLUZTS1txXt6UFeoOlddlo/3fBiRVIZwR7STMMTVmcQOnr9yrKL1PASY9djyWa3678
HO4S31H1/9L3Z0yEjsPqb6Dh4W0m7VJ0p9hLTj4PEt5yr++RjjimB3wkLLK/gAy1jE5mAn1hPize
etC/ZSrC3eQQn5ZePrMpjLMzZB76EadGYgP+IXoABDKPMEynj9qY6cUx6mcSALHHB50tfQ1puAnK
C8RU5icvksdxeCjtU9BhclUKIUkd2DkYI0vg8vIKvwvOo/unzrWJjAJGbjeD11BQexAPVCtHnLUm
isw545V78w/zttGHkIQInQxRHO+9gUWGhEthbhWuo1ioWo9QbGhYxz81qVUueywGZFh+H+mV0WcI
9hkVdCJhXBNvYNqWJ+tpZziimY04VkbSkW176s4u23w9l3AdKpNBf9igRUVnH5XsHDobe4x4QU2F
t82s7+IgINke+RtCrxi+XBqy/Q172JBlHFEmdMJITt8FEbLZe4+nVX2xm0Vf3TYgs44BkIcjQyZ9
tDYAEZY7/kbXfWNtZuJmAEspXVslrNul2SmY+YoqtZjpo3HiylA4UZPUwdv/GqRKfIr5SlrEgE34
tPsUQKdctsdUE6HD4f4H00bPL0trfP7CQwop6HtMu5CQwM4cxU8/LJ3SMkCxdrW9RAHQ7V37VkQ8
uG0a4IpBZEtlmPYUqRxX/GlaJjLHjCyi+5htz3pAV8uOBKLbYxgDB5mHBusfgEsgE9Zm1dEMOW4u
fkNiQi8umbfWQDJicketKH/WeGZTTvt2NlLeA1MMgyBsKwLr36vWFqq+M+PZrXS1SCyFjB3SubxA
oERMO49C9YrB1doXMOIREN9oBt3NM59vqk+7zfABZ/ArWwWVHEKyAWR4pXc7vnf1QRtqu1/ANLSc
b39osHaK0F9hXHgEblRrWXUZ8T3osvr282EufIgGE1YxRiXNcudeRUJ3wHkGjuf0OZ3/Df9r2otb
c+OnARxjWfgUQTlPzQsmn4JN3XipDJ1wMBJJ2jwpXY6r7EZGphflhhiRrIj6QdL0Iifl5OPjafOA
BEvWffYzN5YalgL0ATDjZjc3Kw31FspO1P4FpiujNl8Iftb1YkWXub4LMLz0lG2lIly8JOLYR3+s
FL48T74rG+z5JVXyjP6RsoelkAEhcNr45COO6TkfuDVvuHRdf7g3t78WjX98CyZRZWi9rySOg5Pa
4CdxKx/dLOIiCytLakOqlmCrAQ4Zo2LUE3lJE8bNTxVMWmi6UoGIw7UWnNN8IUJSEYOC6MUSsdGe
NkLFqaL6ESJw2/nvpQxDLcyAAkeb9sowTcm9KSa6jX6/fsu/FWM9O3EeqFufFwpQks5FlhXd8Ixn
PxJJppvoywRwqaKmRrToYdeb+43nKpwotTKxcXqE4h0aKX6Hdn/F3mzxxl4e3aG7cb78k3y6kouT
8OAkW58hkMZ6OcSoq+E+Hz4B0nFEP5+fcTbAQtqmE3YRXdBsp8Bp3F8FeJqfE7OqPakLavuCtKKK
/ms91J5ZBvi0625WIYUV936PQhR8iUpSHc7wj3/fl/RV5gUF08Nvvx4h6mYbviBYtwLFfA770G1w
j/1LpaTaFy8iFgQ+Gz6gw/vMFeF7gL6SjdxKi9gBWn4r2067+0fDHIUW3IcIy4g8SlvvvXowudq2
tUaOmB91/8c36c1GAvVvmGb9XcmprrWbmloMGKoGXwF/7bNbtPO5fIKAXd3Kv/zb1YcYfYKxC7JD
+tkq2LdtgpFI+ncb6InwuwhyV109VuoTmWixPCVRCxHWeVgpvbPlLhXDX77xJG6YbLN+TcJzasoe
wzZ1fbckCcyzeY5xCDWiM1Tz+ZT7zmRorYA/V5Y2nojGmCh+Lx68FvpA59ju5xnqdyOVVmfTaNrL
mOvKlJCA09bI7hbhaBw9QsGbEF7Yutr4m0VLAZarcevGzcADQ7SRO6nnuZ2oR5gYIQ4qc2CwdU3U
NTpKwtP/K4KX/1qx6HbRjoCqsqPR14fY9HaFtfnNjVLVa9GX7zrDi/+cUl70lgC/0FfgMcGXFcuw
tjLJHPg/xuf8EHXbwrOysN2zWIEAvhj0N4Sc7eoH6a8XXgrLcVD8D2We4a6zxIfJAelM5CZQVFmU
XIuKxwydzh/7k6qBfJUu422zmVv5HI5lk3Ql2/8Gld49C18UG+pG6x69wBJYrS6c9EJttZwhgsKy
MjA7I3Z0JKpGx++O6U71MNTVn02x87gYkBys0o1NXqfvCesUCMlc77hm4KbWdIIc8Ej+/cga4JzI
/8UO0VYa7BhZMZbcd4P9AByfBm+DsPxjaE6SScbHVDySFu542ZMZ5FOi7vNCcA7xnR8JcnnmjEYA
c2vk2NBHknroPSdBx+DtkiAtMH7nqa4wMjwMqfU+S+o4nrw9eE6RD0eT/s4y6bDom6OssCtHnpuN
1z8PiTiynA1J40aT2oF8jETGC5SmTfHfqk5E5sBPUYgJih6aygN6cjjuB59sRxdBC4ovSmz0rhu0
BJv/7I63X/6EU2Olp4BZ+Lx7YNzQVBmPHib74xyZhyfwhQ0kXKaRjysKkxXt/RiDOTkgkwWreWJ5
F1NlGrjhcgbuLmZ8leRr0pXd+lreSaVCPT4G/3+3KhMKnrN7sHz2XjdtjGgxF9OO0AEmQ9FPxtpl
E/4485BH2lFhVc16/l1fmdz3q4KEOLwzq4WRogRC6F1flloWnk9cKaHP4eecX4jIIHHtfJLkwaRB
ZpxWlUS1J+qDgWhPUC1Bjpw4Jb6A+7lLjkwbrF5viqSxoth/TiBv9qoia/mE8xVtISXSQkhMVNjF
L/7C4k7deCcGciLt/YH28pgXp+K8I63eUVd0b8NDzIltwVY4UePQJPnOPiCagRYIlDC2/zVAePh5
YpjDUzT/2XrclLTn/XcY8pI91L5gNYZD+7pwkFh8LXVt9HkTXEFV2yTqnxb6UHZED/tDHvsCoafo
PuzCJ8wnqCj976Jh+axb5EPZyIFPPU6R4iR0FBe43YgkuLA+eJ57gbbMvHE+A9OQIXau17QbzMIX
c9ECn8tIuuDkbk9qc8N0pmhcK6zJ2m830XwqO//tkcaiL+DRayb149jrV5p9sczvW/QEOywPSH2c
utBTj8P8VVv12UoeABSymsh7EhZqW/0jTY9Ot0T4kQ8+w2YLta9fSnIrHxsfMnmLFSwNxOEryR4f
CpmK4mzJtSEQAt0ETKgwwVakfpN5EuhkeA4eRIagTrDqVZtuTYSWAw+1tkJF8vJ+Ih8Mftr2GYNL
gZzfGLLfg5MNrErCRoqfyegrkdLpqc/ktG+1a5abO2laJXqQRa0VRwORnhNt/gDNYOTCMrtcXjjJ
82dmu3udwOtvWVT8k5EHkjUtnug0tcu9fLv9STPbW8EuhJPktJ2V6v9c86gDXUVyVJfYvqCXd/1V
IHaQiUmpt8+rs/U+th36f+Jc//lTWCxK8rb9wCMiOXDwXGaA669hVIUBd5qagYk18CzH2EXOiZdp
ESF+Q9fqMOfg1SzD3aRTXO+8wsEkiC0ymt+dS8oIu0W6m7gMoUMAQFlMkhA52JjP26dkIRSZJi+a
dpm+8r5YMpxO4SQhObNF8woeLTUoiwybhftdtoDQml8KIa78STSB5hx5TDEJ6ABcnMswK9K4qVVz
i1UUlOgcqIJlRHTdIlFzFCTY4kdNj3QRI2JQRZuJJaAre485tEBTE0jAt76wHzzXzrRfHcMWDhOS
4+zyEtjV+hPPi/mDVdVbNScwEwindAlBpGLKBDkv8TTu1JWiWeMt+sdqJS7Kw2ObfCD/wn95kvPo
sZ5zgBchgDDKIDxHip+x+w4RnsVS6ZpM6H02SJrqW4A5K2hD2Djk4adENpw7jUOBd2LbESdjgjYv
MP8LTrnqQFXfqEF0moWJMu9XDuHBy1CI8S1Vb4kpK350h259H8llRg1hzS92AIlVOGE/jQTUbveo
4lqYX1IYTzmvEBboXlpUhX6kv75z/pT+QJMDmYi/oxMaH/3pCACza9fnDTJPdOnJkvqgbO6vHxl0
N0kFc7qYuUa3lQXvBoQ1ngzBJmKrOmqg3Tas0r5UhGwCu82Z1HP1ipn1UzjOVJPfOiPKs9tO3RnE
jWzO3T3b3oJmqcGfrQAeqKLIFUF1/uJi6PzVuf7BhadugrEUtkXtXgtAgmO4NAFRaUm4kdnHsvRO
06PEOYwI18rjuWJE6i0bQ6EiEZj82RZiKBLPqDT4iosQ1ABHVdgu/0KC4DxMKWaDX97p0HYCJZNn
muQ5q5gNEsEyT4FH9uBNukSprVTr5lCs1YiJMc3Qp7GuJkuBHszDd2ryJZhOI8FHEfx6zna01siv
aizeTAgE8SGMjLYcRtAqvpUFOHJy01EQCzOypwwZBimizfJ2LRJ4Pi18V3cGGuQs8V+6DLxVsWti
BowJP8xLzOYCJl1lMalViZq+0OqgSHG9aRHEyaPSNE/BwuzYDzKj3+CuR/S7NBYOLLPZ26fOP3Hn
ORQKWpjJufnz66EjGxQN/rjrxbyVGyQiVqpdIW/BpeSWC2PdAU9gNKdO+9xznvSoSjLEMpholfHh
1zuzAEdisCnTCFfluhLXHCjJMc8rO/wo+KvchhKP1ZE36TC4fo1JTuZ5A3mP/MIXKiYa83HASGsH
58IowkSEbLWBT6ss1Jjsa6fuleT7opuMDO22nbi97Pl0KGz7jMHW1KxWSibYVUEPUg+v5tvGKNO3
av/aUYT/W01xsnO6iLx02GyOGYvJdBiF6pvc7C9bX9TbUCXIXuZZgnxKRjeVRCpXjiClZ7eN2lJD
eSL4/Y1F6arKDkRaMPGSmFE1JY+i8r0PVQUTi+BuZbmloXCCiG6V0eFquM3XSm+lWFHyj3zDgJsv
6oINQO5zwh1amNVD5RmRtMGmw1UA3Nt5U0i32PV+l0MPpHBzkSgN4+wKaw/77SwdMiBSVwOd0SAe
4VKkWkSrqk/6m1hsjVsdlrWfv1jEJ/vKLOF18NwsbNYwqvOoh42srggdOJTgFKpXJJ2MmVMnOA8W
nmKT5E+s9bywY9lT9oKi1hVOvP0ewFI7nGrudmsWo5r5gXhXPLh96a5LapCkP7Dgyv9yhDCP7FGX
5Xdx/GQJBofnAu1v+qsdrmE/9pUdizGNVRQrrsZ6EzDLBM7OfuijRbvZ0SCTNuF4kRAdIDOhkZwF
d68VDqKWvr0fMHeKhRBQBpowlNXrdoYPOHMfhXtYfO+CjvlC5uHHg6b+eGYBSOA4Pqqc4BeZNACd
pDKrRmYr7aq+InmzucqiSbDOnBUFSJsiBMSjSSRxB+5ZKb1KEALQZfM4spFMVgHZhz8rfHLgBnx+
FCMjh8F5mxHsklJXkk6w8vBLs8nQ4MY39bymXr9u8FEqFOLY1mQ+jaa8PU+zwukIgGz2g8kW/e5/
7uu4a+251Ffslk2G1Hsp8Z6Htp2jfGHyweaapDXBwhuW5FCnN59Tdz6kcED84thtgUuEzHINRB/a
oyma6XwfESx/UHrrjIuKgYEoeGvt0FJzfXpphrkkM9FNDGjAOKiAMDmgSZ81Mh2r5U0R4wiM9mZ/
1dB1uIM6RW3JOAu66XDlckMiPKTGQ0eOSWOKvRrXe/u2TMpIrbpiRqOKMYxpK1FQdCckoq0LteX4
axOt6NHEu5RITJ6KcV3shn7jhiSBnlKnBgTtXqqIdFfruj78ThXyfnDYL/5euM2+pbh5AAVKTxbd
6aS5x1Ffh111x5LGvYAOMNN4WdnluX6XScPNP02bymBigTPlQVWV6mw9YBGmh5lcKxc7ZesSXXpv
/k4zgqOmpHFvdMpBX+czk1bvamsU1aHYpbYwVaom4dvJfrIXQyYd4MYjoctSDTyypXuJOitE2mid
CN8pjLrmx0HStULvd+eoRyAePqi1vRpFEgLSaJqzDaAcDZNtWkbBxD1vSykJbHOGRIO5OD2kf6aZ
P+AahyxLV000nZErgOrOlhEGhKIsaFSLxuveLlivApEFqbO34lnv3/gAgLSQcjDKf39IhqXEZIar
gGoE18CyWYQhJ1j2bqk021OWxpQQxLCMu7phwjhjUQpph0fXcN7e9VhZGVKm9jyNEBYbAORxtEZZ
J4+TlHBK1eWzlNbJGGR4X92W44DJ28vvYNDOT9HG34QQlfMEpah08B5u66A36ScCH3ZniLQlg/P8
R0BT4+28SlxRW9e5lEU4FXjGD+vXOoTolSNfo2qc9SydgTpxm36TlD+vn5vaPvRWKjXtW9vLiHZx
1K5hy3mu6mIzZ7wmOl78WNek098jH33NMvjNW/xA0SdWTHkyRXXq99Xp7Ak6AKLVql0YMyAPEatj
NqVrYbsy384/6AFdFehTg/TvxuPQfwDbZkoJxTPYpeANPi3Aa5YZE+P1ig/1tsSRM0tZS/Dy/isx
jyU2ddNm6wRzwq4iEh8GCmFmF1oR0Zb1pzx8kkQnLdomdioRC0MH7eTk00Wauj22RnQkdhXfcoVg
BHn6V52GGqsxJYdEAVit7bNE5tk5VmpDUo1YIFW5829RettxsGaFwilo9upQB5u9Pj1id+vLMGiP
P/im4P+Q4e30chw7es30wPkItqCbs1fAljsMiCVy5VQl7IvXYuhFMcuNHQ2SjdCy9Nb+Yc7W2G9e
57SI30IhNtav4bLVbp4kkn0tuQC1El22e1ZaxXpkE3vzxTLtrBbzfWUly2A+J3lF3NmAnfUIN7RX
2ULo1873moj8AMlO2RJiUmv9S5n7Sk4MLMtlGagyvTMCmGEI3Y6HAMToQHb5t8K0IN0kyZ14Px23
l9yrmv763+kKB4klK2SrQEk32OC0nXZOoEuB0e49ayyp4ypxp3bU9beWMbtkrbvQdM6NoW+Pj0sR
u1wNRtQ3iyq0t2hre3ktby2EJTXaHQ/mbk12Im1h9YMgQ1cPT+ActKdH4i8vVlxh0edjPyCj1avk
dR/dNwgPxl71780VSHDv4Wnb4DU5D7V/Mes/QGZTutZH+jjy593+dLznbmCghogb0F1gx2+lPBWa
iidSDKI0XdAZ+Woe+sZbpX7a/ZclBt8Y5ACskuXAgpW/Fwq23kPYZ4EEuYdvY9JyS2h/N292fZp0
+d8RWxw+ifPzMavM5LUT2jg/UUZuvEdcLjs4EL67UXKH8CN4p2SUx5gHfpL57zdzKtWxEBBDHpRJ
oF/0UzoxXJLXlSRViDdDGhs8ZY6joyR5QDEMLV7Uv0UOwaghO/3dwEf4x58vapayke7KpgG3UOvh
pg+8rVGM0ZZT1KHx3FEXuUdLe4YfVckGeA7/8K03FBZ/hKvWF+37gmOaxF7bClzidhNAC95CXKyt
Box7b4DPM6izkkJYLC4fPZGYKwAe3dnLpo0WAoLeKtczBwPx8elKm73K7aNu7JJPIqxKc4P1tSP3
nI5Xe0r0WAJdYuNxyKpPprlG9b3JYir5QoeN6dZhepm5Wg4aZL/2HIJNMCQmJQD9SsVc45cinYFL
J2SEIhUJkkoISYQbVa/q15qg0Swsq+JY/FobBRjCdL8ERidfJ3jSMY7vM9rPg0MJmbpCInnI7Xv4
M4ZFXLWn6lk9h1tk8lLDCWvDZLCS9mxVG8jROnWXFc2m84kzBVmWihMYmiJcZYk6nNc+trKusnZG
JHyf6aDXXaJTumYPX/yzC2moXrRn4xMkXvX89OMPtaYPAJDBuJMnG+ByEoNIMN69B87dEC6a7etY
EhAwfnm5+s2BYuWTtWnVOANhp2QtQW5jfc2aXquj8G30yamYcc1UkGMObxwrZd3i5CIdnHYCMuJi
ATOnJCRQa+a5TER26cJdXwIFqkNWTpBBSmPGSkPpKrLPoO/AxmX/EPd9mZVCmHZGDGejvn0eLm2H
G/pfgTtP9Pw8s2NisU74aIHsnxDvfqHzhMz9X6f+qKJNcxQTNnP6QE5qO1MkWI2cn1yxg2/aktfP
UA0Y/ojuYHjOR0eOfH+z1owgd31YOQjgPcPsjYa3TYrW6+XKWU4Qy5AOKSGV5nMU7mOQ6tlhxWvh
xqmrSCrG9TSt+a1yrBDR2sKAzwUxJk/YXGZh36kHhvwFATevwi+3cXQeEjqzok+W+Lxb+79e8bwf
afD2i5mDNGbkDgZwbkAVZy5q2zqFDjYsEHd2jAxpTcxqPIKk8W4XKcPEsDKM8hlu/p4UgBa0OxmZ
b5wvTm23+X92KwZpZYdg12JKb/aMwm8BslTo/9WwErFdehhfgTjbBFKTACjobUp4W7OUefDCsvOR
2Wr/9xzJsIkmeFAIhtmK70YYmDyuieStLipbxaNuzRSZgIzxw3EI4RbrWXDgLLQzX/oMxihC+jOC
ZbNl2o5MDDuQMamuIgVTAlkn2a0bQRYU+VIqh4wxVdKW2+vjHl1BOuJdnrVPFSdkZmrP4mcS1cps
rh3gw1zyRI0SQfVYgo9LHOFP/UlJ/qR5uCugrQzMX5mp1WGth6nq2QGOWeJ6WG92K9mLsfVD8JIk
VyucbQgFr3eXnlCwhfBe4As01c2d2sGpkB1uO8Ex5Vt/dX7pH/v0yvoy+hEEf83Kpkf+FXaksLNm
EzDYhzsZPznmR37KkZc0MRGYYRxS61giupMR1YLrmpG4BeK9SlWzllbTlTy6Djpc8wHrz35vWax5
f2SNK0QXyK0Zn7k9mU+hkXhKN1Ph2vut1rAQ/7MS8NEpIJ0ViMBPLZhkMkVPXagRnEmNUWDDUuK2
hyIDXAY3kzyKkPwxt3JEePhgBQzQBLWCZjLPaGJDbo+PVv7L/SGlF+CYfMlzN4trrVEpTWa+GB4T
Llum6zwaWxeQ+L9n0mNP49UzVo9WuvLApDTxyEKSCrZXqcRefeQxUSSETWbsBg5LFVKZNJ+c7lCz
KCCSZw/PGv7FRFJbHrI9PXnC8+EjuSIAT+5Qtz58RilZ3bYrTBjUGQiJIPKdWTHuR949a16OWyEJ
pOCLZTiaqWhdANQjPN1sD2g/ZOXlwFJENWtjr6vrFKFlKsF/v8voTXl9Uu026nNFCD1UNRPJpE/c
/MyZNyYuhWrgBnFqyr45iXJqY9GmZJbndD60ZJFuwwAX6aBCoweyUYwjAzfvjEsWXH27TTFSegby
3uaPibWnIorlwj/bDPJeLIxihk7sKXpKzK/2jZ7EOQ1OUTEO7F/G/OftGbKvJvvwWlZwNuZe8utv
eG5PcEnlLRaD817s0aiU5U+oaj4lXW5arwY+PY5jIo8ZvFfV9Q+Kn0lC/aTwsZZXFW96qAhK1RZz
gBjzCPUNWdJ6jkwnSIktG9GcurPVQkijR31slwT9usFieTscRcVNDau7BSTZbZCNhGxyH6ygr3OK
fgPFNSxxx0/4h2tfi4Nbs6rSh5sdDLXFZpVUcieUT4Fdmnlc4TJ3P6Kx3quWtOQMqvsClLDwOG27
EW1PwDTa+wn3q0Qo5tE8b8hbWy0y3+0PEvr5YaBBnor0KuM+YoiWWtsl1wLTG2023eZ5zWDwGBEz
0LAKNblU9WuGyFhv4Ty0k9SC0STPCPf1yXVMbR/ym/h+Mcd38GE1RehD2H3FSRhPHVeGcfb31V7n
H71lNpsKMUZxKjETdM0ZNVEGyYFvu9FwTnEyUAwEYTU793DGvEeBQVi8qTxKovpWXaeg+++F0rmO
MqVwTMLqzD0k+K0q0FqcrOciB4V0/zEsLGElCg1ItHfhzbLrX+VNVZggHipT6Fayl57BJUmUVwtQ
jkoGp4xVzdqPT1t+eNweqYS9bTwDcESB9DC9EI6EL1ClOYPpDrCMfG4WSX0UM1vYbYAjLMAF1y9s
X9Q1XL5GoWPMuPP1b94mmWMLzW0lI5y1Woq7mBe7Ubjf7VHtZZEcOn2DKHyKL86jDBhJcn/7oxfJ
s9RYEkL5TtLseH8ZlmcZpmZecMnrdW+4pAh3haSOqFoouIe08s8taztxSmFZhHftcX898Vi8exDS
K00bJ1bn4OOw9uakAs+/NJCeISKn5pMdsaBYZZhloT6drsPGQ7SBJl1OqN/ZAYKZba1MjYK+0VM3
SXo8PfzaO6JQRKfREMk711bQF3krsbdRB+5apOtpYj+3A/EEeUeqoZOasEayUq7M1JK/drKjY+dO
mPwTpseEVd+7BkSPECCubHNPdExvXE0BAcn205xZmOiaCsXYLV179SMCo+UqDFluFWLcKGfaVSHg
bOX9QtYfecH+XhItImLNwg0XYFIh+i7KpUYSe71NKhg1wcCufFnMIKzEF0l4y4uoznLYsyrzWNjq
GHZ/UzyJ9qADN+ool50hBQHZCORDF3qDtOxcif5dDt8ZccpT+DjccAzIbObJHbUB2n1hlgre/RY+
yrnLn5Y1QA85Wjg4vkR09kcdu4wapwEiqOqTEBqXhTq4xcbFo20kMK6DoOhd7N6OHkt6c4o1DGAa
aALBSx7eEV+3HHQdAJyve7fP0hXWKdWr3EpKG6A8AepOWOUouDhul0PAwlxFFd8eW9tzd/TMHHcD
QcVBtOHLhIMttymmSBCjkDQKLVyOnm3nIAUmHDmoA76OVNL4Tl+Xv/sacS3YG6igIpzSm8WPtQii
j43IDqD7QPmMitfYhZeHeRUtiC5F1Ruh/Wv57mdlLFuPUFjkYPqwkV1UkufDzUG8uFuVb8C5/RGK
l0ooIeDMbCqv0Icp4auXDipAkXAIvfL/L7klR5wsK48KGL1QLGiqPYvkFdnpObsbcAS88BX2gSFs
9Rbd1d8r7I5t2f+5fE3G/R9beVIx/Vyl+Mv+Pk+0VuPGQthInjiUrB2O+pIRrJGiAbaj/nPV+1DU
5d7lEGiRklg6cGrLAHqLxo3mxmzfKb39R6mytZRafdgvHeRpzEUvF7ST94bjB2JGJXrtbdElte51
GeDRCNVFC3WWi9jdQFIon18kEhTCrV63xkM0P1ZSbVQbgz29BYzyxtsX586oeNmYAN95F04zFSb3
oJWYOLxiewqteVfEJS/K2Aqa9tmyo6Yxg6WP12kAwf1mw0ggXgn97w1QBLAea50ZmT/1XEQlN2Lc
HsxHo57s9juF0zSNTTqKdBrtzBz1EWlSD/7rintaRW1Kjny5k2WxT4FkkMvucYBsCciSG8hyxMku
YdxLAwEjwGgdlNtLV1ATlz8/IqeeA/plt45uT6tGZm3ntTYYjw7e5tvCrbOL1aKAK7dBidLIpohl
39lMiiqHR0eNVORLZWTqRnwqpIcc2UGbSDNtCVjB5LEsl7oed35wVhrttu7RQVKu2/FB1ShbGbc5
gyzury/EyilBjp9bkvphT0ISA8MFVyXaE39TjnEI48yvons40AASKakHi/bNg8A1/wHRUSF+pjX7
N9Hf8v+Tg5xhbvOa4BTf+4PpgIFwyyKjdI9xriKtkMduFwb+2SmOWe0kXmY2pEBmmncscMM7dq+V
7cTJew6oze1+LKg94Vp1C/FsDuLv9XxflnJs/PkBFdADPpBy5s1r3RzSUGDjzgkzUanhodzSUvB7
vB13DYefginkgUozh2Go0XaIaL6A5H5lGqOfOEGIFSrQlNNtiZJUeiRkvQIllZI8K0kKJFe1BDpO
KnRzdwjbw4POD5u925SXoPCb0caqSFGV00yyM9em0zoPrfVIyKiwrlVdqarAHUHVDiemeEwDcFdO
eNnYiNrOC3O/ksxslzzBbJwy7QImAJNSXgHkDCU/YigvgvohUhoWmSQLRIw7FEHAeSmkoNyuzbKA
tBqZ5iQIm1CIX/uQaKd1krDV9FkLjtTJT/+3zQTZ/BtSgTtICBAExUt9KqbzRS4WCk5I/BIuv+KL
I4f3jwASsV8UXG/Xz7Jcifsdw8wdgB+1Xfbeo7+DijqFF/Qy8jSCrSPF837Jpd7Ok08EgvLNlUzs
N6kLzIuxdSytBImJeoCgvihbm8CQ44XLb99sZZORG1VbY0EZO3j21e151T+tWiVjZn7cLGpP+lUu
/ZOSj5U1Pbh7zCU5dMuq8WLHjEQIfExutEdgYOmAEbA/GcRIPCjk4OSQGlWFaVS9BZKITXVpcC3y
Yn3o9pxmwM4AUmjRqQuiD1iuYa2JD7t8lt8rtRXzpg3c9Fk69jxJb441rOG8HagOErfFFTJyRG5S
P/WZu0PGg8J2YvuYMWzBD/zo/B47MZ6fM9rnZ3PzqQnzmo5eH0JD+ZzIjmv+SgvJV+qIwdCxlX8a
M1GziDzxSsfDX0dZ5RCGyF94WpzS8oyjeiXbYd94IS7T+LgO9XIjRDJ1X3QbWL/r/LZP0asEJGgh
uYxkniffTgx2+npCGpxvmiawOFaJvH2Hk+tzi/fK73/YUUZ2kYFCJDb7b82j+IUJDOLUpu7w1Idf
32h64aTJkiPZkTmQ+NTmsvZ3LEoNTy3zDxilAp3J3Il+WWgw5U2ZUHW8yWG10thHqTM/XE/iUund
Sr8jIot9WhJiKRAtLzuGrstaG77Bf2Ek5SE1Lqy50FCmLpkU0JImtUfCqYp5D6FJ/6qO4mJ82cbI
7iiConanrgvITknyKPK/zpaH2/LvyQRBANYtUkzYKtzxvmPVueyCQUtMnyWFyPW6IJHAFeUEr9lJ
0H801D7VZa3+MjV4yOcwh0OhkyyYxgqtEiQ1hWeG+mgRPkYnNzFK8ztq2Pa9t+qGVTA9UiiWsbyb
FVNynGC7jK+Aytnf1sf/QcJyf5VtQkOoHLPSNe7XkKkTmpYU559WcpQ4zQU+1hm7ctekgoEr48ft
KwzmBcaOfcCvXYQoPs19QTauYUFhoG7+yfcmp1oMSj904vEKeXbkdgBz1phkr2mmstVtxchgiVsI
wSH8Rm46+OimDc0hDfng2AEa11Ee56yiC/ziLfwxSs3R8WH9qo9ruzKfYxSeBKv87hg3V/gPXoas
W8hFLvnj2uVbDWntr8gIkSXxeNDisQxWrvJPmURVxAjkZfvu30SvlxL/KQI9Xw6ehXUvzfoyXpl0
dPTbFdb/Jtex8x/7L/7u35/hsl4jZI1qo0PJiVyENRTgpD7B/d0RPK4FyOzhn84jJcEFUX23W0hO
uFOBWQbTM8ziAAifi+hvYa/Iakx2arrXYFnobWwqprdOdhgLowJtRIY6irJNrS8Y8OybQJol+ghW
vJFLXZLpiZorUr2xhTPHYHAHUSSjSOvZjJLStVlwIA8eezpDlyjbTnw2gB8X+/QrIp44KlwTOEfD
DW7oCb3yDZ5uV0zYacrbz2ZgBLxWuezclTYtww5Ag13XUtN7DCn+kDbWA77EMpZNRgSQkdsPblrx
/Ehkjlj6tY+l5T7oxGxNUdBRDCoi3NXtYKW544glB+EFXMtT+JAdFNjDl5UE2yEUjK2Ww+T3KaGc
tiIJMTwusWO4EMqr/NBOQwv+TnjGpT2uEoWhOnoFEKIIu9FKJG9X86aH3W+mNDzw1PPXaBAS5d8s
Odf4wgAW/z5UA9HN5SRuDqgdgDQDgcWslcinbNIORiNkejz7VHil/RmjDn3bUCa/ilUiw6zQbI1J
mjOjrpts8nlG0trhxUjVVAcHM7Ps/sHk/g80hCn5qnljSvyjnPvpYdGhtwTrakiBFJxzlCnCPfIz
hKZM5GSh6oPlHCF7MFLB0Vyhbi1Eeqrc68J8Lp1E+UX5l5Df3Q88plMCmsIfEvjpwYgT0ZGIyt3v
XFllFXT7ZRmMx6UrK7r3GxZLkqgLpNJzg9CL4YdB20B/vqAor8dbCEfUS/2Pgpyknm0QjRM4ArVs
JvexT07y9AJJ9yZT/UIi4K2zxkCYtPdbcU1i2xMx5yQkv43jGNa+FNl6b7IlnoNOW/z0lfEUEitU
B2dCk78TIem2PRpqegDH544QTZu35llzs6ern71FAEfEar+cUvxVj/j1BXgaQXPpR/YRP4CWLBxP
Hn0I/Rj8N4HKjlrjcHIwAAavOqk1DfZGAUvtxDBa65Nkz55xKTEtXKnHLPrlhL9ESXIRTlE7m52s
sqI0r3v1Ni+W+GeBgwovlwuY+2Xjy/REp3BP9+88kOZJXhX6AcETiSEqHvyewvxtaIy2cIclYc2v
acgQ9A8HJSqBR1vZE0rvudxFR9hU9nzyVt9Xd1sSfFDSr4/t5gIV13zR6pWz0PN9dmMEJ+1oELiN
WwmX1Q98+PtLP7qbDPD9IRAYr3bojrO76GLuOz5AG1SVlIFbRy8dTnJJnJAtKmdutJmELGmBac7s
dKbzsrZrbzfhMni4FIIMPB0aBXVMKStsYuYPErxuLOYe9lswzlAHpS5xXiFPPyuaubwSL4JIGD01
3rlV+9+jcQhuB2gzQTnQ36ZwQbW/9T8Oocq5FDN5miH0KgoOA89UC1WG46h9PryVVa+j4aWlJZi9
BV3dNgQB2gevCR5uz5vZe5FdKsgEHmjmdCMSSkIuxO/mNXvIcG4xIpT4O/eV7SI95aezEHmpmVMv
aat0K3Ng9VuVLkjueaiPNav1V8Tdnxe/dA0x9vEQ8KB+nj3pLh+PWlDciNBNbrW/p6v2Md49MKQK
kG2Kuor/K8PEALIWaMQ/odT9bQZvbyxtjWScTx4oQYLhu8tSHr8w1gv5ZJoJpLSqSGqlup2cvQ2Y
rgRyaq96ldW78pTSPz6Rumswxi2AYI51dr/TgC7k2jsvA6MauRYvWGQY1f3YsNrfQqIA3rx50SeV
3tL1iFkITa420UG7wo46w6r1bmanWLMs31lU7bs04Aih5miLZhBqtpf10Egu1Hjno9vK5bR9LvZZ
wT3jq8K8uoOwy0AAgwig/zNoppa8aXPkmV9+90IZ87TDUsG2Mn+iMzyQ3q+eSHDtWWdPJv5RwN0o
2qc90O1sFcXSFvcbpTsgRTrlBT16ZBoEXyBubFd21nlPDP6f396ZG0JzM6k/dOziyDy/s9quRbiS
durbafWj3RVe8lBZ0MMR5WTI7e3bgocCRDwvcL++iOhiRTw+Dr+Tgt2uHoPvnOD2Ly1Psif3UQG3
9TdsQAOomqWhCcZT6ZyjXFh7JMmiR5oCl3K7hJJNgufVv2ftZA/2onGRD+cH8QtALjOQnnrk2taC
waQVbjCi8+WgdC5AlV/88DcXJHikqJPKI2cC9Oq03hThOBWkeMOjUeHv5FZq00Lpscg0/jst34ts
7wSxV8T+jZzB4WErdUrqydAzyRE16BMT+C9gYo+KVu8bMMHenGH95ZP4+THUxjSSa/FN++6HV6xZ
fyYjVXnlewX6Dx6aZHENdrTQ7eyeBCh50UWA5F3jE/KHCeQLGBaX+dRTIeNpdXThBTLMYpzhMbEb
44zUGUQgWK3aM4awveOqZKkxSg5p7vLJL4H0Qv7dpdb6X3uAxDxDiQvPa3Daee5AZTqS+6e0E5z9
yov7ltXYCLZv/GCfmWEfr/TwudR8kG72hm/VVWQJqoHELo6GgwcNyWdajaYx48XHJcOqDUByma1V
WPu0TU2+rv+xxVb47zrqs7NW/JpJ/rHezz3oxK0CfnS+aw4NYNIxWSk2VkSixkHV2IkW6L71743U
rxDWDhZpVsVwBTu+W5iNwQuLpfjn8f2ytFM3LhhlFdix5j2SB8rm2+88XJGVADNleibex78OcZOI
0zg4eXiRcPkkdX+AfcEwnkmovqYMRnNbWgN3OEzO05P/zmWZZ7YXtzkPlEvd/aDuoNNFEazvehYA
ph7hhUv/ZYkoyvd7jrCT0TXJmpXbrjARNxfDRjQiKF5XAXoxU+fP6lzr6c8R/f6sxkzArH9TsJ5T
AyGCoRbfVnxdCS4HOIoIVnsY9gCe4i5MY/J/7cyQ+mO/u+sdF8R0H5XzwPxlrzxteLxMqhg1SWEN
2bk2ddCzwmc7Vxn0EE3C0aggVYP8g0YrZMfLGqtNf8V1JtmzkdahzAVOqtVA+IRI+mgMoncOEkE+
wgpzKzL61mGNyJ73UVnoX2aR+kQs8GPmFmqlN3dIvRBnOogmDEc/r1cbukSGsCOIYblZ7InYbKXI
iDjIj/KD/9cm/LkodxlhorVxpZaJpATylu/ACOWVdZNjIVHLhZQsxc1mxxRIJUWDeRKdfBmQVXFf
JqIfigxRVPKlqhER0k2bzs5ehnz+4ByJMxQ1KS/DFxYavZBYsA6A4WHCX88nLffURm9TuKcD2uoG
ZXUudcdHDZfiDVQEjDGNIVxTUCo8fnGrBHvAboFuxAjBjZ23M9ccxHcIvGNfK3jfNryrP0Ow08B4
N43a31YouPLaHFHkZzsUcDhAzb7XbR99d8V5/sr6RmoTlgKVu6prtxufjh85Q2fFPMATkXs85qad
P6FEnGm2ZzxXb3w85m0CQmsc2EP9oHb15BmbMPq2SlCKLHzQiXtfNHHWf30ZqBQFqWlaH29r+1mu
teJUkIdVCbDnw0fGtyjwFsyU+sTeRKOriCLKLfn8Ot2SB2l56oPimo5gbss7BoDgd36Kbvg+EWY4
FR64tA9DsDoBD+5vy/LdO+sReFpkAfcTHVr/QPKg4O/TI+xxoKDFU1JD0w2kSe+g3rB1sqz96Da8
7ej7Fzfk+mQNRD3ZidUQ77463mhZpoeJGbQkjLTrwr7rGshZGy5ij9AOJT2gvmAX22wdfwMWqnGU
n2TFjNw6wQPM4NS702hr+1NIGVMFSkAdglPURO89WIeBvWkrQJ24TxIiFBOgBz/4QK6mAhT4jz8a
ELM4DK66cjAdT9cSEae83sFndIjHZOyBmnhF7kNgnjQeBkDXFFVVk20FTtwIW6uSl5394o7TUnqX
nyCg92emT8kJuf0e3xuwjw0V9OpmEJw2cjAkSHyH8ImdtuPXSBS2ko1cn/vJnhx/Cj83em4ySbpl
1dFjV9sdd8keM3go3G2mCPPwo4qH9djQ2E+ql3X9JDtzd20RVHkuQSN+ctA01UAPuTMru7T2Ju2E
buZ1kcbsrrFno/XB6eopu92d+uaTifIfxpGeG1qYBP2WDS8cmz6JgQ4jtc5NRPIZ3z7mHP2FJLPq
oDwQ4ueyQUlDliHsROKg3iPyLndNAysE12u0i3ReL/N1Bx4YyZE/hEX6HHsDx7WZVXef7S9lLVE4
T7+WX2/JGxtdRKDYSpRe3ia6KFVCsWvwygKQc61VEt7GzYGio8KIjdH/TwGwYoPv7UttUNwDfgM/
TOXyYiJDQx+omu13PyZcm8+YW+BNtP6po5gz/d6DDHCfz91BVtEzYSPmQxK3LSj5ADQLO4lL6iix
FgdmrJUFpAYZU5FPdfONvw1h7a7nKI5+5XsOeeXGGaIYoWI55xnHDIK03A4kh4llpLAOVqP+TF6I
1rYQW/du5tw16TesDqUK2CnPeTZMePAGJjfOp/xQ67jAG9heCnlP2+wz2Sif27rZA2YJfJT5imL8
HBuhMbG3Wp8vUjs3CL9UJm1eNSA2vDIN/5ueMcAgcKrhgnSPB1+yFzVRH1wqKJM12A5VXY9iJrIn
D8F1hTRh4j5do2y18jXGXyGjaI2t1nhT0v/w+mzHIB7OXBy06+eFhPqpOlMcjgnUsS1VvihxipQq
LUxy4oqbbswrRywdtYIhOdvXnlnH1UasRnucmAf7qW+0oCyaGTv+XKt50mivMVuQ8IhdyzzBSSdC
+WKQ7qLPk6P0GL29kpLOcjqk9+cDf+Ik0BuUGF1otZ+gm+GACkSBaziGVCuDF69+GBlEWojKg03K
enThNObxTGCBWGg+ZHL8NRIt8I9o9WaiNxa1EmTwvF3F1CrMVH62FMK1OOgIDRWwViHz6/f03Ve2
BzVRQZj1xTeQBTXMRY/qGyo0NdWM2/tOjf0nrrny3BuUeCmdBw/BJdbRUp1w3FDgH/wI4Aoth5Ff
sBCr4K9TWCs40+MqRdHw86DYEnpMZ+4s2EOHlkKGuSoTNbTQ6lj+qxfFDrH2w1dKuYXIBGPdHQQd
JWH0WOXyKK67q4f/S6iRXAZix0CeKxe6kQhkl3bQW4yrxOjBmldOwf6YFbKZscE6BbLGygECinTg
nPthVCmK2KSGEXDxCsLaInvhi4Jml+WSGYdNJYy5GTGt1dWuKs8PVA1WIPX15+6IFUO0UUEGPIG8
GW2EWq/b3Em5IWc3+U6GigrnQXvng3hPtCIWp4d7abnqQGiU5CcOjVL4kax8vv8EQYmACYX66Aw/
GtmiCvz3oVqw2H0T4JhTrisujdxK8Vd8fhl7ODC2BGwSNTZLyxORe7QFOK0fSQkyWsurK7Ow5sr9
bU6GH9UyNECheQwjti36ajmVl4AtPX1MRK6zVvOFctkGOo5AHtbJuAgIkkbseN5luZ+IRKPsl/KS
rvxsUo7+0p9xVwIgzSiipBKHsFekiM0cH4rZinEI2dEUfHEjVbvdUPXATrebGtlOzRe0SDbVJLxC
YqAmUHde1R4WyEAHhP72icK8dGkaMOzQYzMPr+SP2IcM97QF1SM7U2ha5fvJ9v98qbh7WISZ4iMu
jgRo42JpiH85WBunWO+JfdUKVPinHVME9rRP5/0hx7EhVOHhIvNx9+Cs7jl5bdV26Lw3OAuc2GGK
6V8nAot5Yf2U1fl1nPjJ4/gqw3QUrE0BUMFprMrzwWXg7KY7hSPErGPfJCOujbRhWBz+mq48eYiU
RFfdX+OON4XQhb8Wa9M8E2UE9/fZCo/C6IKCwMCNI70k62ecby/v0PXEbGiPPKUTwkcVWGqdfyBt
zvkL3IIHUDmYPlfmbwLGH8gzrM/PI2vNzse/TWmNlzmO6iBlKy1yIBxFSBNwidkFvZSavxLDpTPM
OnfiW0BsuHW9ZHws/iVdb7LDhV7ZOX0A9tXA58AUDHCdmqutNHokAIGyZWLdyFXGCa87hjfjGXH8
qd2hY7WaQCG6MGsO5WVPRvC6ytyr2UYobtm/EeD6rJIXwvm7Z1g6NfunZRFrsO5QsOrhF+nwTqVr
pdNsT26IwSNKbclWBCKH848NU7JduT6KdAaFCUyK82ZcHpbh6yFWSIQCV1CLBCBNCXADPONc7v3z
z1faEkLstd82ejszI7S6FqZp7o3EI2d6nc1bTQNawCTq2X1KaJm39EZQk0fsIyLIWOMhcnV/nWyZ
NyD91sxPPYpojVew66IEvX7K9DasMDC8qY6/FHsxY2nei2Gky2W53OfbOtCreZINpJ8ZAeS+FezB
r5E8raHq65565cAVSNawp/LP6t4hZtDz64TVC6Rx1BZaKUOa/Dlhd/fr2VeN8XoYkdkRKHbvANF+
fe5P5GJzvZMh6FdJvjJ0ojVQmWR7IuJnHT1ghdIVKPVdHhVY+TJwUsyZpmqgBfw1b9AXf0/xdcS8
wskvZx25iARRUoJRgFcmfPc9jujJsDy81R31GufTriEh5l0N0Ij7UEyfq2BMzeXuBCz7m4p8NLTF
DSkGgcFdxse6ohMu7ymavyNJ5lEnjOq1yYWjwYaNcf+MYRVKOfd8G1/Fqgr0bw1TOPopCYKcByRq
wRLEVNlsjf+41n4cUBeTJ2I/53rHT5Jr9BDUMlljmhbZ2kTjl3MBJFg8PxAR1lm9tuRKcG+4ezaL
TRI/t3+2Av5nSIxNBllGsPJdLpZTx+k0eWgIejJE1lwtKTEgY52vUWZhW2w7NlNk6O0Cmgt0HZrR
dvRXdHAz9xj6uNIFfEcYjkIwdaT37BHPTHqwh67I7ujGmjbZWRotBAEKXRIl6sVfZfwAO0LrPGOy
MpZ8s1re4oo58ZSRypCjFmrdPyEYTPq5ZDBCddRc5QuhpxVo7Oa4pGOhBaE6ggqXGHyMRf0X7pW6
SaMqNhvxdYGJcuitIHpzGrHDpiDCvDTpPRN6DjtXPJAG4X9YmuciZhjI2VQGSz2U9fEcfIWtZa6K
TWbh1IZH1cmVjfEUJkXrTwdcMuivZM/1UfjmNyOCg5FBM4EFNV76NdggY/di8XA2mp/qrhmOQcAJ
1NfLNEBUe5iaCOzuzotG+roiqIisP+ebY1e0Wqa+Ny+7ydFWZMtVHV/mQYIYhhBlGYP9eVH6pxNZ
r4cXxnBboCHBgv8JXSAIGKueiXbPAKjNJ44n/AnUxy2q+G2qbL2Hpge4UHLlixp9YN70zwTT+mc6
VhPvNclwiiukiqXcs72xKCQTEsBKAmfXHKOQXpYe5q60z6IkkaaA91CINYBWYhm7HnSNjnbmZSL+
Udew+3JdpuBZIpFFk/Abb1+baylvRX/kKKYbYHb/OnfwRHwQYrhBZ06RvzLCNvwJySymYT4y8U2Z
ZjSvCyGagHjNrwNyPHhhxgCEOCCxHJFlDjxQPegfuFUNVEFyv7lw+oavtAKLFhM4AK3Vc5Xy++8e
AHqGSmMSloKEW/z/wdheQ4M+V04oNDq2tcdPmWer6Q7nVKyhtPY1ZfVUT1JOcjGVJXE+9gp0RnYN
FjUsOs9j8I4R34sCcoTYsbNDIS9u10hG51VBINZ/DKXkXSWEmLk3sN+n683gVSM1nWmtADtl29h4
WSspTzLFqPqecLYjpxwYi0fUWIFdYdAjTDbMJgfGdXXy2AyEOCWYjD/8ZUk1KsFn4DBfY0cYHRTq
4XJ9nv5CF5yRUEXzm3dx3NoRF+t2GbHGu13BQR1kmnWn54fq4CLX7s8HoySe/LC9O6a7D/oto46E
L1cO88kJ8gvxBDkYd0EDci3u62loZCzsMkeXFrtRq1I7afbYLaDX04RcvxL8AT26yzN5Rge7GXIn
xQpjyl0NUVYqPFUnQKoNztKLg5+tnMCO7H+ma18C+ITA2cO0Zo/9UOa1/9Mijic6xK3YpCK5+KJW
YOlsD/7JawMNG9RsN+ogLFy+ciTaXA0qfp87rjfme2ppkBpbT0RUjUyGC8viH4j5xqkOS3GZapRt
C+mZ7xy2mR44CvxM3HgAF2cuv1fa/yXlyUxxHZpXzjbsHgraSix2WzVq3RiVoy80AHIqwQZ4w3kH
0T1DKUF7CJrEPkQkqMSqF9lkhtpensZbiC4HFOaCdvrkoY3aTrN/bxc/ayX4D8fpWagOuL5gYoDb
USjk/4I5e8uwEDfDhrGDHVsIhq/SyiSx84FOlT4iCNaxMmHuCgiJpWiJhM22HOtp883ah+Mf8S42
KxVWp6PouHiHlUceH6WB879MjBn6N5HWG/YtKwi8twrwYwYW75rVloPAA1fQW0lxODb0OAUc/IP5
Yn+jeZZwLClrvXFZCAwxO76idxpKJoAc9MX5CUdgXud5d1sFnZZOHFf++XxtK+771ffYSny9KX1o
pKQqJTcsYaMcjzzMJNAZ2tRwmy7XfPsnnl/M6nE+LlEhndxiy6g2VNSKK/pbhWzCbo5gMcf5FW4K
gqCRbzabxynqJu11taGTxerNJbxVebBOTO71mcy2NW0rURL4hsjkb49o2mYiHTiCY2J552PQnTS2
GerSXw0yixxRUTKVdi7dC3j4yvsgZUjjKJpLBpx2NW3SbBTS1kNYVXs5NVe2pqx5oJwUfWuuW10l
sHdO33fgs0u5y0iRmOHu567icnDMx/aF8u+MKGDOygsCJ/Ap8hPYvONF2SIbGuNnRD6rQOwp55Rn
ssj1Wo+78qsCYLVN1e2fHCmEbp7iVn1iYe9OOD4LrTFU6x+Me0wYKQmSNNDw7TeOyKyISmiGnSbY
VEkQW+1Eb+e03eEFo/k6aDD+xIkhoSQxiLyoIIGE3AgNX2LJ1j7vqvIf0Kkc83i2HqSpI+k2NQTo
6DFqo6rg/tAK4l9PUwTX9z5aIsRwAf4mqz+lp0EMpZwJS5meP8AK0pQ4AAq3Cc2SXlz5Nxi7BlYL
/ZA6yEz0buozV81js6KRsQynpYytXVDX8x8ST6AIhGR0BdnAYBB+3ycyjt+k1/oypB2EI5r4AV5L
8JO/QeiTgp7CVwlOUHSk48kYS6/Sd55iSQeUp3MsuGJZP0nCFul6UU/72hvu4sWwh4ef/w3FTzWR
2zJYOkDgPwtHuqCAsmWJYruqLTnui3CQPihxUdPuui2AIGKrmkGTxZUl3sqWqFEK8+YPINJnfmEH
I8qVSK9wW+0iTX1qGYBOGVLK8aDqEsXSp5B5ioMCsI8SW3LmhgtugXSI2cevVK3NEqdTsFSdQXig
nPQ9HijSQmBdHY4kic//x85kxnLcvdH4o1eowb+wr6dVPJaqYHZM0cGZfmp04jiog+5Nsuu0oael
ZYUVyg/VWmS69krsnrJ6EhbpvwsSxlc6K8bTHJFvRn9kxp+q6w0YkBDDFx3OCYd+iMiaYSEmVY01
5LxYhMhXgUHrFv4NVsDp9Q8Ny79xGYj+6keLB/7iSoPJYZhQfqxpjbI0PS6PfZb51MeOOTaf+Ukl
fqzRb1sRuZarVr/nkzol/5qNfipTNrtZ/mIOW3MVi7uwdgokHmvQuNuzQml/dL7CpLtjAAZdZxju
XQD4Nhd9iYGG+TpHlTvqawlZFsBXgKEelKAtszWDUlkX6Q1i1+kfw6L8b42Igvgt7P4qKpsC8jef
kV6c6/Xbwto6+3C/kxzPto2TX+Bc2IV3ug7g7EiwpP8ky9gvudqzzOhbiYJMpwlGqcHJ7upr8wrI
LlvFBvPhHcnl5c555LzlJMjp78Y+wlYUUOn1au6s2voB5zPC6zYYsy84egb4vYijCYvHzpnbve+s
XFWLLfrJ6X8f25qh/tHVjehKvCY85yT+BW0CflW4BQQZuK6IhZ7rdbvwZYwTF43h/OOazglWlzX7
wH6bG3lGihpajwvWnNAPtBJQVotjVNYp8+9cmg3Fru5A++SzVep7G1ygJrWJHF6IAtfdPs7ZZGc4
xlQzBqjHJbOH9sN+wO4upQOwLzS+MWJ4uYlreSbFO7YC5/PEH6aoVHOH4CglSZ2UQmO2dC27i44q
yXZaxBu3uQ9+2WMXjMqF2DfABp4U5BlxXH6f9c/JKIaywGLdlDf9r0HQsWa9eT2OEKXsV39IxSVA
YdQ1JdRHFlz68lpJNWUi1HFwAQNTW79NusxcaDbmfGPO1MO1PvSltZobBUB1UV5chHrEtkDJsnvy
PHqK6GY1fkP9sLhOgYBQ/ivwMEzInOWrUYQdhEw0FqtQgmICxVExr3Bv/hlhnvs2BIfs8uPXMqS8
NEMznXjvX3fAEWAPexxlEO9WT9jdxLYL5Q5lF+YFyMwU7wvuYk34qnyuFX11IEr2nqC8TvyKF29X
K3kzVhhBlPBSkFCtvqVxLD1CZzqXvXOpH18b/VzoNO6PJWQEh8J5bQ1o5RI8q2xrmSeFhN/01Wo1
19XMBp0q1YbJ/Xt8xDFdN029Q6+fjuggTDEG2wpj27IsmqgGW1c3HvcfkkZ5yjINDICWHp7fkuD8
j/0aVrIvcPpIku169u25Ikg7EYsf3J2QYGF8J7BHLlL696DqJ/o0jtPKFyPlmq4LLc8NYBqFdk3Z
rZArhosWES0PQPaFQW/rG5UFyRPArHZdPRIy4D+O8pKIJncar/yPoQutG4Ank3060N2qGYkJulLY
xMYm4T1snf0sOaCYbR7CjTKnZA6BGEJLYx9uOwEK7cHSaROYq3kaNXF8dK00ZJN5UIMQsAnDiIZ6
gSwTKOBuGoTMSDCZP90FcTFIulXs4+aBGvCAxb2Uc6km5ZXrmdN/v27bOzTkpOXiXl7vndrx6LqY
zXWAiz5xwr9KVkK4G3nsQ2iUk2PaesZgXqFkI+vUjzps3T+Hy93CyLXFIrDIZMLKxaWvkaMI/pOc
YwnK02jeNyR2E8B1mOkUqfrOW4AtiffoytfmXTswjK1I7swSD5MKBjJu5klC8xSDIZDtHwRvjUsD
U0KNI8t/qH3mQs/PRyWSJQlAQ7oH7U4CAUh81M37dJnxHlp0NujESB95EiU8Kh9fgJ5ynHowR5MZ
uaHkRjt69eoGT9CVBEMSN0ual1SL7SP0Fxs0Qz/ULpWmmAM93sa1r+KhaPevIP0jj5kakM4kEGSO
kGWORUlHrFhagheXi6w1wJ6/FLuAnaGXIB4J00ZCzmnDy7jQKfb5SfQWsU1OWMYV9jZ9SDGFZnXA
cTmy+JhFRcuxdJD94QVUpjKnu40fOXUmUdHbd0u1uk+9C2tnfsa47q1AifxOgCPftjkv/RsmXAVW
Lc58npzYwAyOGeGhOSwsNECit3t+mDxUq/s8VmoGVBBNgJ31WfqcWwZN/eifGJl+mJE08hWQSpYq
NPP06EK4hLLhaJ9tK+26nnfbSZ+h2Ws6lH8rDuydS6o9qMqly0v4ZAXrjFTyBGpn9IGGE0H0HEkh
Q8SMvauwoNe/2w0lL+8fYZIw61d+WUmxecWzFEMbqzRYqCqvBQkoePr6F/F6Wws85cRmCiZ3PIOx
yZxP0eg5+k1Z1AYgWyZ3bLvewnYpITax27v8qDJz7wgR2LIGayRD8KtgpSkFH1DVmfMwGvVU8tkf
mgw20kgnJKapkIsM7TXrE2Ivpqw/e8jLeUcG1M5vtYTJVRH6nufAm1r04NDRdAlNmYhur+yGGNA6
yT+RrdWnJoCKCeUKZM/niRba1iHDsia9qYapv0Ku3YBBqwoBW9qyIylDemzgtFJuI9vvSFcTRjMq
/7AKyt+jGCPt4X/IR74DrbxPM/mNSvy6q6MNIPbW65WEpVxAwrKdFry7x+rh3+3A0PiBUpaPuhG1
eAdIkiFc06I69tNA3SsQQGFS1+Gnv87PXRpkY+ClKl5Em0hMwr/qC4XSJrc7sByq0Se+0lIeGWCb
SA/Gwg4AHRD3urjNKbeGVFQUZKRicSakNi6Z9DklccUH+nEEFRA/ym7sozjpjFgnB0SncwP9jZrq
hqgS/PwzUO5wc8ftQBLxNfaNzjQgLvlvMAGnjZyJ0zbDO6gkwoa3qHMAphMYfCRdUi7doGd8xWct
2BX+3UgQqUu7ghzKUvQ8KMvuE1TrMPCWXp6bcPcrqQFmTnpI2a9w9q2OtSGdjVxtOqUdSiBpeIrk
LjITrUXbf3LSpTfh2BTFanPRA5aIQut1CFV6rrWdriEDyNQMubohAByl4xjvdIMo5CQ1Wg2AUNZ8
ZZLNecuAA7w2X6CV5TdL5AYmny0gMFYOy1SiO58g6pAk5dmLIccxScC2spbAH/JNE1ijM4cfyE6b
VCRlyYZlCkXFU7pEbL7qj6H0P3749Rz06mAKZJ+kVapIsErri2tBdhlpDZO1gxSMJyB+ECPp4OW0
8N/cMZjqDwzPwfzAjACC/beOeAOvy+ZWbh81W8rwbUOxiuFqpjddN4XShGiWCiI/+JI5RixP+Syv
YCUXz6Kicq/sw7iAMmMjJpAsnApB4a5MXEQzdSjUkohFB4FnV8r5shLCXjoM162toj/C4QNFO4p3
rnOTQF9G3+eToIwz9c77W0pX+5JdNARBfREh1K9ScNDLV/lbd/vCqviTadrNidepPl1zykwAwYRN
GRHszsYkDA7K78fF9Z4vyHod/kw+TUYyjjGJK53kQ6JNMR5KJN8ilIVcuOM5Wzdt0gVXTE9pJX7o
Pg25SnpIijGdB/CVlVVJ/pAQhRmZjDS0Vmv4ELkJ/gL6u6PyFrzg/kb+C21AktwkN8iXGIzLB4yX
zK5YIO3Xy05yNpI6HViscHRIEIxmqWEPRRPPzKA5/Fa/LKOAkA66kFCxHEy+Tldjo2hmHOiYF3HF
n85wqOVi1kfGs73f8vDcswCQrJF/pUU757D7Uzs14z6Ec3pT8/mPQNueBAnQpI0MgEycWSe7aW0n
BtXqnL7Zx9S4ZKF6+ND0z7oWKtTz7pRsZgcgy27gsaWkwhiJdW1skbGEpYIir7ORVLeplsS9CcKA
d2FA/0Qi2jxYzDZVDA2ORHopxCmh9S8Rk6PSTDGWSCfO3g3RwNhtlxX7nFd+Ezs5zik1ta4zBXSS
4YGx5xKdOjTBQpl5ne+FRzKtKpL1iUrJhOlAHnzhDf9wLVqwx9intB0NsuQEVnXUeMh5ICNMURMO
+OFU7iINfQkzpQ8Oy0p57fEcDuDrJ6eouaO/l2Sxwo4uLPrKhUTQv3NCa9RGTLNhiuCuhPaowk2N
jyfsL+R+sZXoUdwhLtJuhXOD8K2GlONVuNg/TI4lEqlYHLjbfgjzSZ5yRm+7fQL+jwhifskmqZQm
S1BfvRFepT6vABh+GJgxUm9a+IvMbrgzJesCSnrqMW7Qo1d2p5gxCTuqK0LTT5ng7zbCd22Slwpz
3Uzw9Y6HoUHFWFNHlYB5mRWLktfFQXSjGmcnFZ/vjf3C8RBHFsaOVvMy1BFvsrXeZqIrIArKvBiK
2aKsxuDYVUOEeKojS3BYUGqz+fS7kMm228u6pjpobNQz3zzUX13wsCpIKHBmqsLMmsML0lPYvs2n
o0+t+HrA0DU2pJiUtS+CoH9MDOeMTqaDKm2C9nQSqvz8Gv4QmfcXuDrYApMIYUgC15Vvv+rkeOBz
XGRLVOqugUJUgojYTyih6m4wfaUSir7G94ztDJ4EXWaJ8QqCI+oh84WReXda8JUdlw9swTIvbo4t
s4SSB6Rz75h1skIRTDiy3s1+2y2M6rFGyepLHU1RZV1z3b1q5yGv3uHvYJ/1oM0dP7ol8M5iUbLC
JE++GbUxG0WLTxaLC+O6pbpb8xRSXC7YVP2Ks1Rj+teOmvIh/nEjlUhs7+ythMo2l/UhTMi7wWXd
bX07K8QMoFSD/9B9KANxyYOZ56YGN+LUVcZbbgNCyXpRtdOGffkmueze7oTRT9R/IQkCloRGyJZx
ylCKcprAdL9WqHPZfMxMBYcySDbgBVcNdA9Z/UASt2+TKdO1jNo7E442G79hXKx9aFiUFP8BqJBg
FdxIda1GLjkZRYM1WcfrziDw4H6snJV9RbUoTxoxzuMZXDYZSewCePwttOr2+tdNTNl3ORNM6GdS
jiHY8LmaFfSiOtYQQyK0wIegV1bot0PWI8WVViHy2/Yt59zI1EcFbfWpOC7Pn1lpJTxX2SWdFPrr
f4hcyKBUf9QFIGY9fZuRx8nP/anjkh6z7aS9xbecaZ/5T0Hetdv3KwFSlT3pP+uCt3ofefE/O0o7
86T+kh6aD4wzgr3SgYTJyk2zw1a76gNa1zPQJ7UIdizjEvFKvva2YFFjzuaTG1EjGwU13Po7wSIp
p/0ST8i9gzbUbCtJVMnBqutw/UmkZA/4M0aAiIu2OUCHYnEaIfZPMwM1n5qLfBLxssm7DoEEguAJ
fmaCucEHFast74DI8ryo/20rMSPV7FNRqWspNPzd62lzr1sZWyvgTbCpf1/K/eVsgf9rjR0pAKM2
u9eJq8EIGcePKPHvJAMWBtJ+CmEjQia651jw8dti2tVTiaHSeV1dECYFnZaoncd2ieh/LAUnp6En
JDVDGQjpkEMMoVeBE2nngL35UWukJhhBG8bttCZrKmzfnELgTRUdYcKf12VgRCVTqiPyLHPz3L+w
ll1jPLGJ+pX3Wkg+zvGP/xLCLjlJ40EY0bNHN3qBIacX/4f64p/Zh9zoH2kyZannVALHFYkkmztK
W9iwfxUJVX7uRylPy2Fz0Sz0TTtHc+7ph70mGmmbpxWRLsgV3qrnZgTJ9TEyvvH4Q+o8OJefG5YK
YrxYv7/LgkJjSPBDCq4uwR2SwxbrRslsqqjB7fOy9FUf7wd1Ui0qeRtPtN//9WsMsiAPmcClTgFf
fiYEpCFEYO4hXrRvioTcsdPxaxdwOFSfjj3ZXmaWXFS70jeYs8AvMyttrmG/TAQcI5Wrz0XyNRcH
eNilQsd9Qq2dd5MT1hidXXdsBDNsxhKu7rFm9p1bVYLE1h/pXcRqC+rAomLQZRQvzhQXyHtqN04X
3chzu014qQkrRB28YnCJeSa6ZdZmiwFKebXR38BHVJoFNxqlcWEfEFAXEBiHffdb4Jr4URWb54Dq
5A3qbaupFWJKW3noeRQPePDdVVGkjepu9UvwSx215Sz7hCdRAuCJE5WqedRSmza6CzhVREfPVtiZ
CP/qvsHRndKhioemwEOqsIaEU5z6RZfgVsz/9lPxL7QcxESa/AmPO8PGfhwH39zJlKeNuKrRqOAk
cYhem/WthHBpjbibH+mBNLWJXCHe/UGLCFgQx20emA+T1MFxpiIug8fW5a5UgiPT+Fv+9h8XPqxA
BioNB4oUGOpyIbT7Ywtvv5jWikz+huWcQpyrwVo0bX1caVWqFXQn6XX9H/7hgW2sA02SXa9sWiKo
T+VcpwQA2ae5rlhVKUbtTni8rh3pvuWyR644WhiAQAq9fspWZ7GckhVZg3jXVYfByK12KPmUn5A2
z0EBtB/TW0ZtUtWlQOE5VdXsrumy+4UvSz7/7yw/jSSac9kTsV0gLa+TB+zTpXXlEImV7vB6yy9h
DMjMCn4D+IiTWhVZguP7pbhcjx/qp1X1XQcHvSG1cH9TAmWFuaVx7Sc8d/aU33uic6YHi6ZRKhHE
FOjr40XweLMjaYkJuPpaG7J0zgM8oi2S2Q7V0lxueEGOMr4u6qj6X9Mm2l0OYOcFfmXbvLu9Cx2t
eP2M62SFCRsLwu1/aaw4MrJWY8zWbWPNguMDC4R7UVVoczgCFMur5XnwZu2st8fZ5l9fy8xvWva2
JRVCdenKjPCYio2aJiQMKhXN3Y0pETgW5+AUgPr0ZD/qnzvY8C2joEyAOqRL+HsWwD7joQ+U1BTW
X4jntQgkeqrZbEYDUmQe3QVcnntKORWiyFjWF2LwTUHKw47qIrM9rM7DxMapPBmMfnrOsySqaoBO
NhBbn5aD280SdS4XVEJhKxrZqTRSz957SuA4BNo8Jv8FAIqrNUHONLH5QvW3sE9hOqwqciQysQ8F
rHoZaeZzakfjzj+StxApnJyAJeIiWJDQMXE2wt2JgouhlfJfQxjbk7zOA+b45O5yhrnt3TT30iLK
xrp0QvSe4SnGThAYwGgDx2GCmep7Dwu428vBCM8F+qVRPhOihQoo2PI0Gxy7/nm8iL4S6H8Gglsc
oCUxQ2qyZoiEKcPllOPS4a4pky/YhRXG5B0mxcjN7PZYZLt/8xwezHzvX6nc/4WpjF8eCZhasXWN
jUj9KJBwtSlMhUnv2veYP8C/h67Q0q+SOY5Y8p+kbMqKSkl/MYjgAKYhdZIYnQdqXs3A2SDqwNHw
Bils1ylVf+ilS4yCCayWlseLpa+WOQ6FJWbke+l/DHZuGFnwH2IgfTwy2dxbzQcl/mRBI0tHinHp
P7+BkDfHNBj4135ltPV4WVGJCA6TpubHNffyPfABzPlbcpanwhb5PjlAnMQ8jh4TBPAeJXNNfeoB
mi3CQB5Wzuef55bPwKbSmIsRql5Da2PCxTXNUVrueZwWi2hFTXL1KZiwv9/ndvyzGMbwxtvZK6dr
qfUHr/qTFoKRdhJBUBqB7AGj+Y5m3FVhfHylq1JW2dLdoqhgW1nlDty9IxMVP1HZrv03V0SbFizQ
vMwTCtsOAeQyxvo8Ybwfa2WDvc+QuOQVxnf7LAYSxwyzIlNGCCa6pnylsFiW1Ch+zsaecyfGsRjs
Jw/OluXWiB1t8RpfID3F0lBrw7H0S6Jx8g/5IGYcvGqy0k97zKFhPOYl6p7zMtdbaP8iGXIkb6OL
BSZEEL52hbqMvRuwXQ+JhPeEnbC8SViQvohk50hmNEAKtdnNTiXQWjda/kry66H0EfX7KzwmI4jj
PKa3P2rzokJagnBJMH++DL76W0mZ8jzIdBRzTtF3Bag/bJD7Q8z61Vf0WytmSsO5WzRTcYYge2KM
tOvQg9q7YSLmfZevcXIveU5I+RAl0LCkM+XYUtqtX9bSoz2l/50TPkX7vqE1IzUe1FofQQJBVr5F
YEHhoaxNTuWPGwnkI7qnsJ9Pj3SWcFb00fatvoJK5dBN+jhPWIeDxUfORP8Wfv72BiHRKFXamj24
OuRlR9RbdfWFZHy+yI4fkAsc8jDXs+KYkvbKRsE7DVBVU1ScXqi76lYGU2BYLt1FUYABjpC5Vs7J
YPW0vY20vUjvNW4uqE9SJCb9dE5WxpQI/Xu3S0zB/i105LEtiOcKBi7Z8/9epVoFgSc538s98aNt
/E+W3asWd+FnbwiptpaUubmgCCKTH/8ydVlxnxTQLgS452ecSVbBZmPDJw93Qzzoe3T7Da4uHwkm
LIFZhBXkRqvTpN+oamrn/Q8oGJeDy0nxPpzJPF05ljdKdK1RMJwM9061c/GFlNr2U4GAkPE5Yk7A
9pKO0Gfc235IZ4XW8pBhVLiMQMU3Wn32hj582+6PXLge0VuDiyKx6Jwo6Drq//4tesgOBz+dQv8D
Mf1jQ0nkJWASDGjULZvKsGCXFOnVtSitJD4AnnUPY8gP7SNcwf03j3QJ0bzMJloChq3duoKH1fDO
r8CTUi2OHmabeMSJMo2G6G3caYIYWynRvmDvqsslqDVheWi40sSs+N92euRVa0FBtmWWhaPo0oGL
qJkTWTkZmSTkZ8f5pC7gHXTTHcgq7coUSaK5YFe/blDfaWBgcvpC1xvb7FggM5kjoktBQRcOKRxM
DOxcf66LHIMZibQkhlLU4ZRlkbk+/OcFsS3jP+iHYEyHdLOcitVUcpxsQwsSmDyGViw1NmdkAKd9
IN2lxIT2iW9LG3toIVnESA7Hu3dqLYZ2IpDeHSS8PMZjGElRCRoEfiTX2EAUIJ8aH7WDbCfr0drY
Oa6CF9iBG7oAaXLUGjNLH/LiYbQQOOjufqiCn5nEaiYwx0pbBnI36KqM59xY/dNvUjpyQ03laso/
J5lLsX6RfmM95WbRhvYyubUSTTlHJtwzGY6rx4n977Aqj+h7frewAKA6/ydJuPKYRpwCwQbU9khY
FotWpz0NA95eus8cMDZc5eY6zugaOTL1k2TreOL97O5aheBuN/seO1ERe4PsBpV1+ovxFau8FL+o
+3jW6mBqkL5bTRbtkPZiqB/yRrjvC+fPoEArr7cYdfB/5AcY3zATCNYRSkdx2n/6OTYfUHBIP0Ij
57uhJWoGujy8jVyA79SBa5WbiRh/KWA8rskky3HfsE7xaNRA/zsSL7BFkM9wwqNLZRuupBZ5va3d
ahZdcaSOiCYVnKhjLTH9ALwbBZ+QijDmo4G6Lk+alJg4Q1H2x27PxYURIaU7/uLEpBqcQZpwv/Zp
K8fg+FaP/WiygZU3LKvkdPFJANiyr2Sk7dIgvbQjE94HakyENEkK20FqDvldsrKRnfHMEZtE9uQ+
NsHoi9e+yeY9LudpmVT0NyjFxYUlj9YVglDnCjdwmtdH1QKmbXmoxOcxlLrsY9OW5/XjuofJl1Bp
REpj0kEb6Y+GdYZU2KF7cq0zO98ujg+guDZ2dPoFfUu5/wLJAxfty9R8/cQuxIiNNlxD2N+eYW4b
NrlIzBHpxTRa0iR/FLLGH4tfrV6f9RUU7gj1cUdkyfjThGa6BgSKR5WjtksQLLyIztxe9EYjKb6O
5uOIrb7XHlpEbWTXX5kLIm3B6FbKhtZHHTPGDABb6gAk2Emncztf8D229rz3QNUpR9ICatSYGBbP
4TgD7JL/5OhrCyy2h+I26cJYWhkzdPphlM7davuYDYC/PdzYvvFInz8Onp1k+akmpRPoaZYOku/u
CBtwxkQWAK4pM0S9kUrZz/XHkzRjJkVP4Z7VYUh7vUqGMBR1+Eugc2A95VThmdSefFK8ucrWINe5
fmk2fD85plE/SVJjHHkM/uHZIscB4BCOxnUoS+2cbDOZHJjgsK0+G1BUDbp59PB/PaPZTTyghH7c
LkAwgfDgaD4cZcIWVKPjPAOLsgScrpybXeF2vWhoLv6p8ESVqURM8zFPUeXde466HdpKiFvkF8/1
uJgGtCGNcqCX4B0pL+6746Jb1uGVGb+MWg2/hTJ+RH3iJoDUga+ULTtKAfnIzTAZqbfQiaLIDbD6
zkoFW9JOih4IijXuXFpG7edYzdWISPxGfjIepNEiRLS3H6FOTWnmT9y0VvzRQp/6fis/GL7J/ywD
E7XSezEn+4d83nMfW7BFGZIiGtyFSwpebzzbDLyDQcubwyDVHsajJfHu4BqCCbgicrjsAgZdAPu0
brR8AX2zY9gY5B/KIm6d4JCoPMDicFzBFC6XygdprrD0AHBwD+bXov2uLsJxc4bD++JZijE5OUTU
9AuuZUeYJT7GHOP5R0EINvFDHpCcvz5Lvgd54MO08jvT55vUxTOHIFaEA38YoIu3yU828ndWCTYB
K+JUu606DuHY9Ziex9Bh2IHsxXFk05Ltpr9HCbEKNSiaXlIYefR/3BDoCGZQnP4JnaGsNZjdh7bo
Vk/3lnjxuRmaA+h38q77kcEiwPx3zcB5xmBtEETOqEnB8TwUWhVdo3KSC+E6BeTLx8UnQhO+UyYY
iTmFQiOd0qSfOok30G/CdXOZ5ynuUUxw2JWARFVUCyQheMAgMUQ7fsoMa0qrMsTgYFOIs4HIrulh
8LkEJ5EvoMxNNtDsio6C5T3aBlvVSOtcGOO5OzaA8mMLgUlLfoAs8h221Dwh2H4HveOsTNsR85Jc
0aFVqnX4OZRTP9tqKyZgToAL2axG5f8+PRabfzuT7vpjFeIMne8Lr7QQDWTZO7gNFIIBhUymCk/h
5dV21lpbRera2/53VppXe/x2ci6Ifk+7HgOSDoGTn1XsJLwdSHtrDNn0zkGhNB1NE5BSzygmAq3/
bb7EwIN8VSIKEt0jrS3ozxFUHxSSC55PhZnm4U8ifoMQrFhCK6brJTKyR0TIKYbCovTo/xu+sHhQ
0Inp0qcYcecdleXcL+9zeZjURBck4Zc1JpqlGISPr2oPvL7jnapYTGM54RskUjqWoCO0ELXk5Z3A
b+biDorzvU+aox8BFHRu+niBIdxWOdMdmLqJv2HjH7chHbDweXaJpJXVByXswkRDysEhF3dVTF7d
0lqBeYWvGPvpCkShfv3J4EcAqghDOss4ss5bmTpIiEIgFuM7j9Xt+sdeTZaoXUBvD0h4qedSY6RE
y4Zp19EDNUks6/XoYaRH/xp9yFG2UfqLdEQRpwB21nliEQSwbBt7zIxOouwVjTSeRaeQG19ouEXB
ExOY/yRMmZWxv2cwnahnvCn93ECxEgk58tbkRoo/WUrXIO7Ym/oyHgjd1UJRWe1fwrGUE4qfwOuT
SsdnUsOMvzb4GOs2ERVKXtNVUperWuoBvia9iM94+UZePgz36hHISbfC1vrivVIgc1HFO0EaGkXY
qKFSEQ+p0On/v59scOuoWr+Tg6Mt0d92I2NsKHsr7Rt4XI2KyIdZOUHjzZ2iam59gHbch87DObFA
4yAyqi24My+DDOLw8IziMFcKwSILhYWPYcysn6nUO+5cxAMFfA1zUHnExaL4EHtXwWUEd5icSm+H
L5SLx/+aM3eeQN8S99JI73SXb7PNWNn5SASfZTKa5ixPb/IvMbbPn88KgGfeaI5Hs/uOyz9i3+ZT
IdMTQxlVOCG0J/J1k4vl1ZgUY0ePKLDFiiwDA+Nn4xZtcyyLjmrtnAnRjQnr5DDFUS7OZbvHSYmZ
5Ta15Vig/GIpSv3Jn5vFqC6Aa7HCCN28mAOtb4tcER/JeqGB/tTEa8iioOqpTegL3z+dEhHz+nS9
zYgWeQMKdwHA6d8JdbiuLT11GZuCYMZbQbzeiSLYbHHiDQz8nJyXD913KW+fS5ntOt2qe/9FwO7N
3YE7tfx7gfiifXnofiz/xO5VU/WjDi35srGECEXckRm5h8iptf2WBCAZuf4i/g8GCLC7IsOw3nSV
zvQ/Yev1lV4z8xBEJuH/uSUlHhcDrMINZA3hgbuqWECqVt4oqLw2+GQ0NdrMSMh4j2SFnBe0Wumn
3WJ2VNcns+/N9MFeaYZBfa+m/Xu0rSGZjmnYXRlxLdOCXgmqcFS6UKvOb1BFseDuBUOG1HtFc4vM
pU4JL5hFLfhlesB3RPfX6SPBTZV9pI3WflR1zwqZ5LlE1TmtkTD/cwDdvbJgcW4lY82pGioPMbVz
aTiVxrQKdv7RyJLZPJ88Sg7XdRfoDk/corBbcLQIUEgv+ahlIS9jeCCqbefORWBmD+N/TCrkZLIQ
ylIAnEey4E30I4a95Thp0iy+xVRx4+CTcf+eRGvSYhH2kfPgu8pTz7iQufY5I38U2TQoEX5aANUp
r4eDMpamtgEyg7wp/mWVBoBwoB10m6VhoN7/7TJRTiuEChs/X3O5dWr5gg8FgRLOlsG6WPuNP049
loybAc8iojhs5v0JBs6WTqTFlVIGUJI6XfTyKVrr5HXGnQZD3yG6Fp9FXHBQwLCehSk2//iWV9yj
kRBJ4kYnLTWxhKpt4tV9ysqK3p8EAPUsgS3g7YZg0GwtICMMxY5RfqHMn4/QXBZVyPYJJNua3OP5
qXNcLB7WBaHRdekodYrPSdxtgG23USpRl4Om8cAWDwPwGA6384c1XgpcmJ0Q56DUQiJfBbV1K7tc
Crk1XJTUb9xZbr5huApHxbx2keY9x63zl2yG+TaqAp4DqRxg2WAjgQ4dqJckzb3yZGHMke+eC7pa
/E7rqquwaK/pO45wupMpK7iAK/YKGErXdHo2papcJr7xKDoEXiyUyzKOt0u/LZlDF2ZoFe/2OjkE
bsSRUyaA6ETmwRNv0/VrdwYs6tdKhjyTIz1llSTeIRjbCF3C6klCSoTZA8mKA9W4eIkHJSJNwe8N
b6Ebeu+fXNUraufNuEodPIh4EFSKMcTkyz8EjHOwnW0mn19j1v1rQQObcnZk/SqxhmRWeEtvgejV
IBC0jvOr7qFs4haKoPqauEyoyCww/LMp44RW5s5Zk9RUyFKo4vhXBJ58S7Ax0/jLAyK4EoUjjvCf
U96rScv/K5meMY+nfA3J6PfSyIK2Kp/QUf+THED5v6i+wvPf0KZspxauBksisDNFpjENxRwtTu+Y
CcaC4GViX4mY0d/svmeICaxkkxxTNErOKy8jTWRW1PBXV4kjAJm9N20ySS++IJxUv95lSp0VLODv
04bXaZOnJSMykbAGjLEdtjRbEBduEthlpPxZeHF5rk0YR/qAe+irjMOdwzKLbh6KM0a6KYFXqqyI
+dC+ZlvcWJnZhxlkUon79B0UVxw+hMDOFQYi3miL0cJAbogsuX58Lq9yk1nC7wBp2hrJUGR4K2ke
bfQqJt1+nJ4kcFpko1QjFkqcvCvtgmVFFKaeRu4aQoOrX5iM8sZcYhimgIdy/01hkweKYBZ1XK2m
BfYiUXQjEUCcw/dUP9FUjDLTheVihfFHAV5jr7heMOVKsbySyXc695JcoK3O+Ct+b2YjQzLgjJjy
2n6zhf4MhUxrF3IegpE+3O8VJ1WSvvP8YWLkPmGY9VS6W7I3FJ7bojeFaEX/Z7ejw6H7X4UMuAPr
Sj7TPG4ZZmmhJvVgD/R0DjZBVj8iOtvm9AuHCVPfq2PsXqOBjLsVN8F9rfNOH2JlrZ9gjk05a73e
RRT6uIYtQMw4xJBphSTsyikRdIn1RzGf6SpUpVTp5EdKhWPvQlwedRnn64CM9xrXn68+q/Duq/0b
QqqK959isQmpOHTsPv6RF7s2CYEbTsZIQwEhJwrMoxkYtv+Lv/kzJxVYiao3A8IOaToJrSuZmJKV
lG5RRnhzO1Rn6YXMvuu+UIJO430l4CaJJ9Q/H3jWGiHri5nsePqodHssf6vC1BGQQY7U5py4z2J/
eZShbA2WPpRPhob/1+LJ6paE40OLYU7xOWYxmxjtekPQL9iKgJw7gw1hXLx0FQkAivGT+60pYfJ7
F3p7ysUtYV6DNyJfh0Ggw0B3JRi2RgY4YqJeFjI15iwWn8lDfxX5WXY8IoU+sQsRw5aMEWf4cJMw
auF7DD7VHQhmJvW9VICoTXJ4oL8i/4EnCeDTimg+05pLQXGKXoDyxQKH9vMA4M+WgGtFo7GaV2je
8XvO98yG4FdXhQpviSPgHEtmixuoBXbs9I1i9mPmR3Lq+heV3yNGA5w+84Pbjn0DUM8wWJ3vqPnC
KZCOb/ZCD0qMvH/mlyq7wZZX3YVDlhLiTlhKLtLyml5EXRbwnCkMMtwbawo52roRKYOVzrFTYntl
bPski8LG4nEyFhlX//E5Kz2ue2iicz1ULqcEVfZrizuIJui8aTG8oxqKeoEysa/mvdY9MN4b1mMJ
HkayetB/w+cq2zuJRdvtstx0s4g2OOH3jZ6FKcuX9YvKONcg3nslkn1D3GdK4dT2w1PAYFvz/90U
C21/bcLLVvFuBMcgrrFQgIBYMdvngUpi1tASiXJ6YEEj2EIVWQObi+T9qzQ2EeIl1911asxF0eZI
3D49Q8FszPCpBixO0arjaFPbyZ4mZMGfoWTkpzaUW4nBClF30JPjTHHK1W2HyWE+MnsOVXfKPanc
rPOKjOc0/OIDea30bIAcNQ/RUuj13wus6JYo/zRg0Yi1grivshP2oCkJue4k6NFA9pLgsIqx2F4i
3Qg17rVJctXg4nZHNUsyfjEfhCvmqBINLZ7lQFTmH5W3Ay/Zst+5pl/OSw0oxFEXjLX5hfhDJQtc
h1RjXM08QsW8H8/u/+YjsLfadFs2m+HZUoWfkvgqqPvwOeoIhfwuL4dHF9ym3RCURG73AMge+4HV
4L1WnNT/OpYtcXPEVjNIKmRlAC5HkD2PiB/NDCSsRWIj/oQx04/NN1IMbP9EAcV2owfQtWrPYdbP
54tM9s/joBlW/PDGe+KER2k07NzOkR7DGit9OKasukZWkXtO8jKQz30W940dIWFiOtN5E1g3FXII
eQ0obVoeZtDBSd2sD7EWn8bGm/5VJDCilwiMuFRvbolzWYogr/9jqhzbtRbhB74qeM9qSFsbboaG
29gykKQdhM0TP7bnJRgpghuA2/VxknpGOou514UQhYq7xwtQheV2cwdUfbGNpymip9zumg37todF
KQzhPOPu3Ck4ENZsvWaIjh52r/TiRoiaNU4O7KFSjTzC+YiGYU3yejqS5bA5PXuIGFLChJdWa/BF
L6e8qDvtsw2uzstFm7GRFQIOh7FgI/qNJDEen8OP743aQvISg5NE//WY3RUAXiN33iJ+aX3aZ4aL
WHES10lKUz/SPqTd081Kwzcw9PDpKgSFJ6CQeSc/qdmsNZzBIRweswfcU+GKCIY0wnUu0/wVnyb5
l+YIf9qi3EeHJiun8M/0GGurSXfc33CYjZVe9mJxeVHYiTmKrBEhMwULmbO/FpHAqhI2kfuHK2g3
U+/bVzsLdsHWjHErFH76+rVaLa9/9BQ7YHcNsH8KFFnc7bTSsKi+jqKDVfF6n/PjU8pbPE9r7e9X
2z7eqNNMcPhAGOIY3JOzwa69K4vG0QwpjNJ3EAXGm5FwiT76uT965//EpLcQx0x9YCyINIf/Jkkw
MVPkHJMI1zNusoGJ6OY06wIGzOJtBLruchRoQ5NzpR4tcYD9vh/vT6FeDbjINhOmhiMas/W/FGrQ
w/OSEzhml9fuq4Ie4t/p7UmQktA5J2w7a/4u1XpN06RZNLgf+fGPgVcMbavn5Mwc1aq9p/ba3zlI
TueDc84FQVp8ZtolfiVljxTfNhUVkFv8CU1KV8/I6T6dc2ftQyXEPiJ1JyHWz3phcwnARaGEOZgt
w2ui0/9df7QNrMoUIoedBCdLSHr0FfQHc5JL2gzrZjlzO5PYAiQsEwpR25oUS5m72+DFj80davLo
gLlnAuzrvUz/tKs+N//feQYpXomqzo8Tyrl1k4cQ2HQpZkEmDAbOyhFhcjJwuGFQjIhrL5m2GnZG
PmmTlqy6onoWleETGnBz+uC9u4reodbBBvS0wWmtlQq3Q0OtM9MJf7dqK5dT7cRQBryRcrXoo0s/
BkAinamnezE9lrL60lg8OXZvv5Ts0A8LNSHXKYbS6Coh9EzAspgHM2chtALC7UYnDeDA0ML6+xcF
XymK8po9dJpfQuEi0nx8jimgya2mafncOgO2BHuCxTWcHLGHjEEIrEnbAqRx8wxZOtT/hImf7VdM
Ni0MNf+Y5OoT6+9qUVPNJQaUNvJukCs9H1ZqoG8wLaYApgzgGy8VY7fqPivvqX37hJGCmCjnRAwe
uIHzod0DiY0ji26cPOgayNM8unA0WAZXuUaQuVhEq+xTKoJcSp/Y0lPRzwc7ihWKxOBAOGvVb/wK
e+FvKYCDGbz0VtO5b9OPyXcgZbXvXa8P9dRxXI+uNaD9RYDUrzO9CxdPMXj+Re3jf7zOr4z1hxD0
6auHnbcgDFf8+YclNcVussDdiFts4RgcVywgVlcrdxXfiF9uEV9C7m8+ywNBz+w9o4o9ZutVvgCn
Bw0gabZItpB5nj0B5RBrva71KArKJPe3sGQ9+Pa0UXYyZheGpHyC8sEpRvFT6C09xt5a26nV3kJo
/1OvnW0JXALpZErRoolKR8dbDX52RklFhcDZJ0EGr425OerN29eRHTStVNHv/cg1mqDTWff9e4M3
w4vT6ttvm2ZpGyIFEryMSFXM4l5W98yxyQVhrR1baUJfPO13DSFL20kvHVjxbcdAisb0NaWDBYvQ
Y9OFtp2q5KeAkHSPzgrVAgKq+VerecGSij7pAjwH5KL4IAQYWdTikWwn2NwE0vzZ4oMQ+hunouVq
BiRkQFLAxl97CfeaPGEh/BBsIhW9LaKz+9YCtvsuFhN+69vMy9sihuarfs26CRfoajqQTMJAsijo
ZQonbgQQGIZOicCcSH6owSZpMJbHN3AKMRr21kuZILP0lAChyGoFL1/YhWb04FA1vYNFjTTE6Vf2
RngwHHazJYHHMas04DCWEfGif7HVhpqn8Djnx3gABt80G/6TwHOMeZT+UpTIofguanft1g+Csy1E
wMrKBdQjjsM+CZKo2sWNR8xKlqeQw7r+niutvyf5SKnRzG8XakBgjj5SaArXa+AaoOKkGNlRJm2J
SVzQcFmz0lYxEf5sY7eD8Slb+LunK0qwX4a2PyS6l5Mc18njZq1be+sjfh5+BUvzXlnl2zjYV57f
j+CGIGmHYZJlG0HbT184Q5fjS5sxP2x6zDwU8Qi55v9Y53TfE5vvSK78+B4wodgtpBL9yfsk8CXi
nvu3MmS+6vjpvo4fuf+9BgV05nYdFzEZTsUUC0Uhgi61JYHgsoauulIwvYJyJ9o3HrvkJJa7zE/m
xtcAIPH/pTcvHrs5VrNYlYWUR/KCV3pEv/MT/mYVGkqKKkrWqG/BNAsUgGw1Gmh/Q6tjvoxKJJbL
gOVZ96k6zIEdhy5P2FiJu16LVC0l8B+Lqum5PklxTR5+isnE5lrsGVqLTqRCb+83++Bn5begzpu8
m0jA89IJMSkyNZROZNx5aFsqxIwWLhwRciuyvwYJFtrQ5+slZDXgrhU5yeHKSgGcumcX3bnbwinU
qbQcQSgjAfAv0NI56CWpHwUwBUUVBzUkW4e6Zj7y0T8ohEFtsTyMcZwvi486xNypDCyS8ufYsqnd
sWm/5HifijWql4D8XS5h3ZJQmwD8lGBBPt+GxV5jP4yAWxWHCgysBblBYSvOIeM2EyP6C5ySAHf8
VtHIeWySsYfiOi8HJdqBBPCpLCX4+pCbEVg+c5sOaKL1VEJctUIbAzJEjHVyVgLUB0kueaTr5vgj
K2MdAPoX1qgwf5JNDJArzupg8f4QW599/4/Y3fZ5p9Q+DhH7ERIlspNPU+85ATH2d+aESY1wUgba
viQe3q9I7otzNImQPtZgXs2VKJfGVyYbjga1UjtUpRcRMY/5K3NXcaAtCzpoVv2utOfqOM7foUU5
cJQkZEIs7f2d3wysqRo3BeCUEpArSw61VRixQMC0yMliJ9A+OcKJ9ciLI4EEY1Wk57Kq05cFFO3i
/gjx46x/wRPKUoAg7G2ma3IQbg5jV3IhhT7Vrfpsku3lM8K7PODT5RWhn/JUR2GCPBAQdmX5QUqN
rlriaCHOTB5H6dAfLaU5bUPeKgHbTBoJyhhSfsuoIzjGm61ITDRFWlTCJboeUSHRwCyhbo1g+XkU
VpwvqUagRFar30PoUnTMA1xVPythkupMKCB4XEv6KHvncKTwPWJw8VFAm3ufCnYbTIYiBrcS4M4U
BXJ0IbumHJfNbwms9/kJSjBlIGw92MV4Js79xmogGNLS/qyviaQGR9LQjLpUJZDrxWtax4QWNE+v
tDmWb5u1sGBKKw5V2P0wotzjpBiKYqNm8spuz0hr9o85dYnDuFHE6pDnGY+W3AjvKJu+EAKONlkZ
02a4J3PatOLlp58pAtkjPg1qDJDkWvpyAJRwAVKzQ38s+UDDDci2C/Yh4TCQZ6/xuBXc65pKuQTp
HBdkdCPj2h8/Yk4g+CPLya3NgeJUs6PHgxWxf08bU1vc/t7C0Nb+cxmWhmHPqKQhjc6mKyW8rY8u
ILZXm3qI7KD5QDSLjR3IYHl2Jo3MBgRjiGJ8MPvYJrgTSeKAUlReSJoKQHsy46hQQNNZPabFOsH3
Xick8ZfE8lUpyzJ9ce9Q8CMsWf7Ip0eY+3aQR+uJm3bWDPBeRBStUXUFgfWlVuQe3XRfIdJgG/1K
9ND+m+hKykqv/cmNmGw+2QVs5z8jTSaSj5E+AnRYSNmzma52ql+IH+Elaqrh6qAgVQ8tkc0Sn50d
fyI7DBty9omwAJ4NYy1eCDNut2df9qoZk04sVJd1StaKphOakZistjP1xgkUpq2yAh3XUe1iSKjN
/+Aw1WoDSq/EscTuDk900OBkdKFeWVZtRYW6enPGb6L9A0PsoVD6R52ayUW44Bm5sbf+AOJfJ5ty
NXmSmdkWb9jSRS/FR7QDD8FabMH6v+yELKb0uNVX4pazEdlrynAJ/TRrc6o89hX0ePGzYIi2s6eS
A+lO8QtRHK9BO0tvuEGjXoPw0+sf/94PMfaDH8xbS6oXSbOqEGHuBNZxUDxcas+3g2H87MjA7/jT
jJzsR2ZpptwFkfYM+gC1SNpK90VdkmeSeed2HLOTIcsAIbAwdzOx3LBk8dzVuGDrSsRInRn5DYYE
wquOfc+8cI2VZ2pjyqkXvyWFTszLM2Sw1aOs+jdww6Sxi9wiEfDVdFfJgVDpct+qsUO0Act0JhFC
+HrWBA5IECD7g69VfnLKX9CzlIbAYXXqi9Oh/RSxuGz17LMnGSD2v5tiYoQIAoF70mIBZ5LABrQl
4HblimjoVqvN6sGPMA76bkb90bmcBy7Z1dYFdkgBbXHO8RyGh9MMtrlzPdhIybmYnQJBiozFrGYu
diikdUd/SlKLlAJDOAASrUqOHZy9zKyORftzbjR7ecwWwxl3q3K3CNEwDZEkyED/VhZ9vtnA07QK
VynL93hPwWdrRYKb4cO93OEgIjFjYOI1hkmjV80F/qTFz3HXWGG075tgqmPkYtTqHzN73510JhPL
lAqcz2aQ6ziFB5IDsuks3BccmPUqgNdeigZgv1txj8vDXSd89k7n8eJtSFLW/wmmYVwElw1AgNKj
HnxNB0CxUYpinNuuY2zLdSETTkHRyenPboc4m1LHEuRWmGBok3Ch5XT+ymuNIzep2PULle+/9dPs
PYG8hSy2J2K58H8aQZN8qoj0gKNjQxiMxKjMgwuV3jcPl/QmrvM+3LW4FG7w9SZOWSFabJFowspB
Uf8PliXH+PZ78nEhlZixwrIga6/HoWiAhI+TwPZ2gMi98s0r94juAygBCsJCDASQgpcFEiV0TMow
nKc4BI2+pE8CIJjcJjVXPoaXaXYDH+R/z9viNRRL3GIzWXpcM1Fh31Vi3GsCcLZ3r2iVxaCJg04d
7kCa6jdS6s72nvHGG4Z6B4qGgutMAtyz1ezYPW3TQllVLVDKKNIaQ39RdF38U2c79eeHHz/XVhc9
DEjkdSUzMDKsREzVykxV47pQ79ELUd3uPedvTGsa/sFXBSiUM1EgsT+EWupaoNMp/+S4/SdJvgCM
sp/kA8IkxIN0COtjqWpY6ZnBIm/hL/k5jBAHEo+X9F1ZXX8lKA8lVxbKx5WvUEcm8PhRQw55x1aL
N/MJY7kCNZ+jdAu4sNNg5sIA1RQBukc5nyXvkUtSjr7idfxwc2ul0UB1Y3vkU9fJzoiYHOIgs4cC
cXHrdXySwUq33FErsIZELP6++J7NKH4FJBuA279HQRpuwDF/EwAMkV+iLq1th462kYFT5BYZO4vH
kuaHkmZT6Z8SV4jFf49coQ8+cpoZ5UmCTKzhi1U0m1FMU5aHsTI8+XbPvmjK1Hr43wOFM5UuF1Qk
MwYg2ow+t6GfEELbjkPL5BxqpgugflnW7c61aiAoqR32ZO8pAuxZprFnAazyj4Ej+sQKkMUuBbRl
ijw5SnSb0Mo59IxBdAWKZ6QfwSVvtQZ49SUz/rw6eFylRtBZSBGubjVz7BhxSWZ42yjDpOJkbpxZ
WfQQy4Gh+a3NXbP7q/aYWrBBwLXFa9Io8MJvocV1/wncN34+hQFDqXHiKuCLMacXxY7Pjt1FvmD+
L45QD5iHRO6UFd9DPoULYjJ2ieyDgDV0tUnE//4PlFZ2S8cOpGK+VzMrFnNWYQ6M1H0PBxO7paeP
Twkup606q9K1OmyyPdla4wF89EzMwBKkZyqCBX8gB6QL5we5RY8AU475e3IyOK9sncNzFDl6LNfM
SvMKvFlhx1o6Ml8UD3aVp31wyKGbV4WPngbeCPFh40klGubm9kG7Kc5HNB0AgG6dQ7wCXJ5nzdIo
cMYgI5mNGTy6V2oh+0pQl1mWh0wUHpFiBMj1Va2+duOVxKbjoeYNHAh86skGKfRdyokM5WCtaZlm
aJDSk6DqkKD1eWHCCYmstRcR24hpRx0CKgeBYLaesKZ/pM/+eeP5KECk7/Mu33Gbrxzfmfg9fxHf
tsaqqJjXMmGkaTqGEj8RzYSG6zLaSw132A0AxfOZKAES3JKxxVFAy2tUKz8FqPqK0pHQXRDMq/kl
fq+IjDFzSC8D4r9jFrxrfHIMyftVKeggpIcM3P2UXmFNG/PzGCfHFO37vdFPXv45tXUaFfVibjaG
iKpbPg4nE1HLBPrpDwg+plIf8wMznmPCxZz38zUEQ80PjbGTCdAutgb5UaYVPZiy0GxjOVknwR2K
cHpfIgDcly5gG7DlkCl6LDNYt0iEXerO7AJpj0Gx+6vKq9md6nC5KCZk0vnUbSPyMLAJJDYAl0zj
Q08kJQ0k+cIBrki3+3zMSH5/+SCM31AXx9wv03SUTjB1KBmXf/k3aZ52S56sEipCCTDMnNrfIJAK
NEJn+YTCRT+6YKF7gt/Z/URQKdjs6UZZHjEkaA62DON3JJ5FLsDPSObD7qyPOCRxilyp86UGtWmf
WyUaB95ZUYAtWJ2s2TvviAaiqAyo4kamzyi1yVSzPX3GoLpV/ubwEIn1ZS3HZ/Nl5tz1HUMR3ERm
W3JNSLDNcfZcLyY8lbq3nFO3lPWGa74hA/w6LJIMuq480lrbFB1B1E4nkBKVfJVVBt/yhItejFXv
/s9KZGP3Wd4EX/U18ChZKCPG6BE38ikmIfvNlOVqCcNQBGaqtU2xjenJCf3dxr6QLqI7TJw6MUdP
5JARzDEZMhw57ObMnXJOd29EyvcKHxuwFNb9rc/56GYKxtdVNkqJyEPSZ1rzC1dHXaeXwf17T20S
XCoDIp/9rLC6cnxI3RIfs8Xx2Qllyd3kHEHcey2A7rX0SOvNfKZUKS3wMEy4YMHCIl+Ml/ihwT6C
UOCWpv6AFDsdohkvtFjwgsN/4wlIOsaQhRVHDUvfQqTNzthtofSz1HoiYNXjkcWo4xxLgWCPE5MJ
F61EfPIR/+j3Ggy/TA8d9TWuEIj0UJpsTKB59oSoqp8dpepk+C/hd4WeBCLrR22dd2tRUZhBQLkE
NTQLQuqFPabCDm2BXXqLxoHwLaftsiw7y3fYcHDoIkiUJYwJzNSEHTJWg22e9kuxAOBliuCFTtZo
dosKwz+zf5XUJKAVr+ka6lh9n7HHP4D/YlGCmHVi7UhxYksdjwb8pugfzrucIvXoOCiDme+9c6oM
D7fXt8og7MJNMJC4dSLv8sGXVRE0Yw/Aw45Xr9/PvOakfnqhjGo1KsbJfJtoIkf9f7Ubq55Pd7vT
1NgcOatkr1lphDUi37YX6pHK1RT25tguWdkBOSVtJkHFqQArBp5gjHlmLHb5GE4s7+X6lDEwCWbY
XBWR4wc6iyw+KZxAD06/PI6RZ/SwyfqO5w+Zpmaf9XJuWbj+Vc4wOo2lFfFKDm3kU9ovRMkaDXMf
Kx2DXqD/PYzLbqciU6z9NQjWKbEUYhoJBL4477Z8vophA/wGsbsVrTgXn8BUVovRh7j6BB4XcD9/
Y0uLDG+6XhFnsH2tKEnaNWHA3k2VxiGazoFnBmUZ5dRAY4R7OP8rlNehyDcoYat+fn1wM6tiHiKa
q/HuyIsfLRHEjraS6pMf5MbuyVVxlDaWlBg2xuYq57ZqtgBc83mvLJOxT6AP68joGzyW8xRzlGTl
ee7P9VznJTdC+ydD05duvidbtB9ouT10Ln1QuzfEBqy3CzvmrcLPRG6qrZAfO8B/7rd4Go4uvG9a
VTg2WQgdEx/MiH9oimoHEyAUNnBNQQdZq34LWoSrSCqpCb0lm6iCkVEstGuN9avycGES5scLVTHp
lROGQMz0LC5ZoP09ZLF1R47M2T9+X2I/jTzO1qWhy8YN1d/a2ylFV9F/csow0gtHWBB9hKwp8yzH
nb0lDqROFquCTA8WN8FYwqW6IoqXPJltP+Pr410kfJGM4aeLaFww4OgwUs8h1Q3MQvzY8FNSNnh3
oE9UJ97NHHehHmYH7VRiB1q+MUEtytjuNaML8rLCSO9iQNSG2YnHDZ+RqedYbnDHiNnA2VVlMSge
jtqc503BvgJfKhksH8sC2i3Ku2mdT0e/QTF+00VvU1J4qJPQZTvthpR4/uPhM2WbTZrgT9+KN+Gm
+7Obshb+OsdDbGP1uTLkjU6iZPeRz1g7U0vOH/SsdFqQgdcwCN4ZUlQgCDIK6zixa2ZgNlju1eiR
p6ebKm/SrLIk+ObjPJomlAnPQhiSxF0KuAZZ4erbmtRctSex2u0J11sUydLh6naBnbXVebl47JHs
SxzcW85cBU7rTJa02hSrE2dW+8ORx6gD8ESyLw3HsoYkxjZKUMo+FIaqjRZeSk4WrpmSxZViH196
9f+P+x5qwfLlPbSiP4UASLB9jF8huRBZpX8hk3ljb9InnqW28ADIjWS7ojVLPvHz1nlr17tvZHA3
h/ylIBJdUS9Nznbhc/5OfYWpbihRYHbyAosKIDMmywk26+Hel6QXBH0FZZgr1kb4jQXtXAWYPTDS
CKr7bFFwlmJVsPblA/xF0+cHGXoCDVBlmauXmQsLVK4lh8VGNreg818kHMxcJNqNsmzTJvog5HWZ
s+dJ+239YAwrdSg5d3lPbP/qkhl7oaMb9K9IR+gU6BzXq92tcWqPKi/fovsFeIRel7o7BYpF3WP5
VPzH7/eJzhysAWUVLPDaPM9TC9bcG/R+kQ6O5CPZInC+TAUqhXNAkbcU1erqqmSn9g442wgP3Y9x
xs/zReaie9kmDcxZjVA2BWqOwLjlkZxiA6jnqWbIH1mmleKfqPNZk0WPOvRhCKsErQeCl+6isgIY
CUUDDSlfN9VJpTtMWpZ3EammLabeA87uaDG1YnZRrmMYynIqN98ouoWHIXHmdsT4fjx5PMJ4QFzc
Gs7F9MKuQUqh1ApOF7Q4XriMMdJUkJd2Vct+rx7+e5CNOSIcO1b4ZF4jatrOxOg3PkECsTDPalx2
Ih1YpMVkEfRIkw0YNY3jIyowm4Rx9urRhQ7fk/5kC/zA5iUhgOyTJLPHObLZqsHCqauiQB8gqTno
gjYX897AQtro1z3fcNkkNqZ4Rs1wE0WTrwfxU2zh2HQ0ctkuRlL2Obof7cD6xDpa61Uva7XNFQns
qRILTpVHhJiA9WrN2ArzjHoQhsQXVuygsyxr7nLd2EseKI7j1MZpLIIpRE7L8aJbniKPGUHy1oth
JLBwZ9UlDFFfReluBuPmLiBjLV6g5EFKteT40SRiZBmXGCh8aH+lv/xfq8suOudBo38zVBnmDX1z
mbrs0bs8KTLWOkEnD06E3H3fpigiLXIZqIi5Ud3lEsLFxIictFH+dKg1FIb8WJeCyMpHHFGFJsXt
AKN+i/EQ7gHYvC3Hhz/oLE9SzTMbOTlF1U6PXynHMpAzAdWebjq5JAPB7P+wggYB+8sr/qpNxNS+
Gs25DX8S55xNENxwUfi6oOLxDFsuPb7d3Laec2YtVv3hYwBGB8tl4XDa+0/1G0vQOsD/H28z0t1C
gwrYYGIjNror721aBpSWFSsVSuC1fhMSsap93nzFQJ3sJGFrSj3gHjUX0dut+e4xCEb+TFxKpjac
WrD2XoTsRmmDWug+wM3vjKIls/FST8A5Q4yCkgRgi0WtlBHgGooKYqu8aLDASAUsiH+rfDdAc5Tl
9saGHeaUqtddPVPk0h8ujBWXtwCBoB5y5UWCfYLrc76uO2b7NO/7kg5wTntvOQ2AF++kGl94A1Dm
x4I3VtIfB/QuhIfVRST0QYyEtM3UZnekYCEaqXls/QVe/Wxqgf2azVmADudZCv9UU9NYv2XVuxQP
nJZB9w+1ZxpNB2MZ2mGnCsIBV408+J1VrI5ZFXpkemrs2uekKLevlEMBM1PbY/z7uaM9QSXFoPcy
XxCG6eD2MTIf6ZIHpFFP8ehdpGczHef8H88RTa9UKjaK82Eo2wI3EiKU0ucbSrObENNTl0T3+6ox
+THuK9Dm52onWXJabKHUTIqP9T6K3QhroQ14jTGGc5+aANNEd89kSoV5X4NF9DGyKb9Z6t8YHaQS
Fx/jDNlNsjNifLVfVx/9CsTlFeqntDs/Yaq+H/cLInCd8MhuWmMlmL/kgMfR4zYINenZ+uyG1Y7+
2HPP4HOStJsyvMDfJZXDBo9NZu7gIHgOvE+9QujzpyVhGmHEzDhmvSlP15THMkYNvlW0l8gAc4jn
DeGyTpVUv4xSXovEhl7GSoSkHU2S35+7dv1obJAv+KBry89tZT0Hq7T6vr0Ui7QF9GACfunH/FUV
0k0HutZpb6IY+9UhWBGECO15PcGZbiXQwkoHloeVbiY/96Mw1vcIOBwS1efRRec+NrIdFtiPfCJ4
d7ZLIDX4fXigclV0Plk+Wplq8rDfDxWQ27fZYAwlR4adOZslzBMuX2S4O1xG1Icc7tY3LQ/pcXj+
0Nlxad4I0ueUbAZGNPYWQ6MsDBl76sYopEJTpy9MgcBb4QurD9MCK8AUAreS5PVWIxfjOg8Stvie
S7dmCRE4jNuE2NfgFyS6A2FoxgVvKyprTRp+GPv7mH1AGpL+C6sxiw+D9nBJQuXCxAQCXfSo7LPi
rPsWrwovbbqEVu0M2bllimT5+EPHxjDzEiTd8UmVnCnWAOoDRr/q2CBGP4bZrXHeIntwh+MV2Yy5
BE/wm6U5Q0B4y7Fgli+y8GItj+49HsUI+JFfXK0VxVPT93J9oPYbQQ/itTg2CMjf8zBTXCQTApPs
eANYJP8bdPkW+JMOwO3y7ZzJjkrY9hq6H/ZuLAFMUf3xpPyhdh8BqgyfogKLJyyunvYBeZiF8ee8
9wuSujJE35fIS44zzygsCV1jtWYa6K8uuMWEUbY0UHqz7fZ0YMR4gHolAaAPN3+fPy1Dmm8ZHksN
Mropk9aLYYdL9YIAFnAHGzUUexX6PMgQk1+GWY4JOzJmJ/lAnJte+vNZUWZyDbYqoOpakRwVyZcW
kszB3bOE0YIWdDuxk2goHl/K1tFKUplzlS+4GJ9SQHdwZxl48dBM1LP9BOF4bWVh3aedyZsywwQl
SL4ZCfz03QUypB94jvMv97oFvWetRl4OVwAA1uzTkq7XBGV8rsG5wo3ogjhVRgICmGhXzxkiV2sV
UjRiXSEiMQCHWxxyEd90AMJCJW+6Bq/Z1gJfNTJ3atRQcwtpTCA1kGaPRaNO/2lE3e0Cmrg//Le9
pmuJZ26oltO5XC6KkVbhqrMPeiVUV4xC6XDMMz+N9kU65X5wcHdZvcCVjVP4t7+DY6p+A9IqeXjs
VG5Iyhs5KU4EHqE0kB1U5sdvl5hJDQsJjHeueOHj5wI7U1w7tLRDLSefFzy8E58+PuhZLBDZIAq0
Hp3qM6B33V9HGfMdjPYX50sTZXmGlNSDpKvSIgVeqgwgxm6QomqdXmqClQaEDqHjpia9nyfTwUw4
Fx3roP6ZLdo6Y/gECXPIter1yDZ7LaEKVSZhhQz6HhvsIaejDLhhdm7idyE2L0X/AWtpMLdOCblg
LTDyQHHRW3rg1zrcjQI9ZQ7JNTvtZvVXY1Pcoi9jTsCO7N3V76WR+LzD7o1LphId0iWyOjIlHJDW
fQjyQT54zEyHk5R+sCZ/EDAy5Ho93PXZVY0kHx9gZ6B+A+Owwegv4qTq/+sLMZl2S+wcDMKzvOFM
9tYnmhV3YBOK5Oczh5wQJhPLYpnBqW14UO2MDeSzwzhZTlxoToFS3iISI/CbMocicOhMHmxCGgtG
pPf0E/tlMY13JlXRV28BncJjcfD7iARU7h1VGDyF9E9aEqSIh5o7i8BwCMfCY4Fhwqns3VHCGq8I
GnIdg7yVlOBCfd6VUapzXyOfEw9uHBVz2EcuuTzLd+9/78c7JYzyIE5lcibS/RU9v52x5YP76E40
zU6fRbO3dsrFSNXCWPzFukbMyDVh8l/FFX8kN3dPzgfgmJPJV+bKzzYXQsKPlieI7B0utoBlBUZz
yghnZd4Xq/GrDM+HKBlk+uNXaoejCZxzcgGWWVeF6isrLqdmMLzDTAxvuZJSRyGUvvJv5jI7xGfY
MhgIHWdYW+9RK8Xaj2ief8XMjHYw/kZIW8/P6hSsSZ0jGV6vu2KsT+JnuJ1m2r0VNRa/9i9Ju/fT
4O1ARytw64RJqnsXy1Jv7v6ivftD+8kzoEBDSPXStQmxeZSdp/mnQpPLQb36x8kxtnIdbjoM2BGN
yMb5yeovUG/VEB0V4x3BEpyIR0D67AKe7REeIHIMPFba+rltKvaFZcBgQBYkgpHd2Mt21h+vYHNE
OWUaPuNAY7i9CS6YhIS319OG36S4oVMfBn5fdgLNodYZrFhSNWMAm9YvUUDMvAH8aqFofJuqTrNK
kS7Anx5NzKM9wJw8ql08yjAMUiqN6dn9w9Wet4rvBortJaR82AF3iWBG2OO76whoNXk7XMY3379/
aj1IFRgCbsA6LUBNfZqQ2As0Y7kBjqeSzxmD98mtt0xvx4rFcg+X3R65nz1UtMJUiLb7xNVyWYR2
orho3DdpcrO1JvqXvQqlMQbk29FvPgRbS8BzRISr8aT4CmTKsntXe+5sGkWQdE7gUZGOhYejH/xG
NYbq4fgZLVnJz7J5GUgGskYpRH3inpzd0wdSkMwgaN2SK7HG0bGPpPu07a08O1GzT/ah07pqqW76
wx4uuY/kJmp779PamQzMPld16rF1YZbMIrwg5W6sTpxhLyScQ7GSWsDJTyluqvlDFer+DUvexb/4
VauH2ZgAYqwTWT8iscny7sRYjwF0QqlhcbVfOdIlpCEATKHwPm0W4mfJKZg9LlwjTuWRZ9mcViU8
H9eDcugwTn8UG8NQ4ilSylLfBApT8Nlg5HnyxlFHE2knLieljbmY1bcm+5FKz24MZoYn5Kf7/zve
ZlRZMR9tmyo+C5ksxYzrOpzqhq6u3KtB3xh5bPF1yOfkCyshtsO6ZLwO+pL5PEhSmZHb/GlXrVaQ
FZD0tqbqwFf2RN6JO4UzyE0h77F8qIKepUK/Y+2p8o0cB6ERhnH6PykQhsVtERIGHVlghRCCGfe8
NgUk69gWWIl7gxVMDH4VDYgA5K3E8Yh+YmN/diMnhDqWd7Z8roq5BLXz+9wKi0WIMAy9GdZpyvoi
bkQ56oaR4gMiJpfJuTqlqCQp4MgAa6MuV3BIsTsU4hIcT7/X1hEFC2P6wpiQ9n+JsnNCOCnhM3RO
rzh3ZSPOggN1L78EO9wwS8FfT1w2CNnmPiw+BDyTxfPp0vX1mToktTuVnQrKaULGF32DadleYQtr
9NgDEAEv7cC48zmDTa65IZEl2V3UZYaIDmpbSbao8apvl95Ik0XtvZ9G5pMoiQYnVu5y4h5+zscH
XfHmz37z/uqdDenIwwgthFUg+T4du+J0dXr71kJo1o1yUSaxAweMHD4qlq6v17liDtsiu3N8Nx8k
I9g7OSBJL42+v/EJgnXGWKYcPT+iwRqFtUDRWWTeMmYFPZuPXJx/rwj7kXesDieVEwLWZ+8xdLYb
+/JtTqKkoSdOcZnf+Cjc2SbhnEeMsIUdAXG1C5WHo7+RtHuvo3NsBv7qdFR31AGgPZH9MFgon+ex
tmBJD6hHSm8Sp85Phcmx7COENaT9s0Z3sUpsOLAX+TDr08QHOVilQ+mcgx1d8MkgUZ5XQAuu7C/R
r4zFKA77RG8qxdFsmpEb/jWDBUnu0hayVDhhu8tjy5848PMssLhrDhBWseuiWCLglRAd+ZnXNoT1
ORtIu4Aa03t9cKGGp67LaMNolOWzM3VJcydWU3CFP8lfkk3eLoEVkNPnWC0ojFPenl/MQ6aBxx1P
ji6AFZlMFbwlVLL33hv80COXaBQKZYO9v5aHAZV2ph3QJsLbQNJyCVeNrtVayFLSlyIdE/Bu4iDm
uc730ZBXo4PRehymoMBwcgHvxdwgpkIMeqxPDxZKgBGmXYNL4cW9JbpbGP4iChNVheZeK3e0goAd
LJ5DGlcfnor5FpaXPEqlirGaG0S10a23dLoCJqMBG+YCXoKE5mVwWCvur3y9dWoYmrQcniGjewPs
ZNX7dyQzpQYe0Q/HumKv5u5Qwpmikxa6D3qTuzBNNijpdQvrcTLcMiWbdjGY1BLh5s4gWq/VW7/z
ex+1jkUvcuDjj64+4XFW4d6oH44MBm60DqsCocsVASN8BbdO7If7Rqkju8DIAFLWtjGrEPgCg13+
xOq/IfWzCy8MMKR8U9tUgjljDz2ZLoKl+4LkRE5I/+rAu/VWBRNQCk51EIf3/zSfaeTOCj/sc7OH
9GBgM1txn2ox7TvmFGtwQCG5W2t4FH6jL98O3smcf7GHp8PzMpdkjCzF7tbV0rztzqJry3wZXfmX
blioAr0hirattkBogYovKboFWGgEHlWWJ0zcHyAwYazGKamYC6+7GRlumBimWWvjHmkAl5g72PmO
teAtfbd9G1Nba9+hmX4ta5rcyDU91MnED35MRRRJnuB04od2YTMYWucaSJFhZCwrMSttqMdKHzhr
4lW69/F4VuKLg65cZ5Em2dmMJJnbnGFCR2s+mFUqFhGt+e9vesgPHemKY3MozUEuwz+vWwyLE/7g
qB3KGbptXOlqnxYLR03JFnr1zpn5M6pp01fodMsXC9K50a9M136jFenxLAU755vQQqhGxzZteW+u
dvKp1Q0zChrv8dL4vjSyk0A7N+xosKZSCzPX7xMbiqSLRkgI4eIP5zQwb6uPmCuJ0wTkc0X6sT5A
s8LBaHfmAND3q+QbAckH86W4Au58oQQEjvm3LWMTudvHtt2URaS8JEmS6L2HDnKayaPS+dtdETrj
fwVN7BXbBQhJNMEXGm1mqWTAa/yj0NsoYaR2IHamRGhWoTHQ4+sCSwvvZc1QMlZtrfppQ4D85Amr
chUZXqXH9l2pF3gnJWNaNh7dd5coqSamALr7GYQKRaIaUBoJucfTo3t4tj1xB9WwXkI0MFc5TS37
XQJJhuJ1y1kEgmraBd3ZRMcB8d4EnqtR33BUEL2yJT2xKCIjOxq2HhqhA7nmCfsA8BWQOL/z7unh
/UECy86Cr4mVCBp+fCb/F1p08jqQHBKcOD11nA6U4BJE2FoNoV3mtShfDUu0XXargZ04C+O81GiR
Wh7CeVX3av32AWTYZPFB7FO2F/eO2JAC9MgYnb4QhZCpX1ZfU4Yx56gliac12N+zYzmm/XLaS+Vx
MGSUDbomkjoq+0o53ggFtu69+5EJdyXWCkc/dleYQal8uFFK1K+VQ2Dy5zX+flSnpqMc8BalBxD4
NE66chQQwoAYcatqOtnrwDJvk3LRBnRw+YcQgI99unaBJy1XV4OXww364Gc/9sW0mJj6xlKrJaE9
d4adtULnaxhg2HGYPS3plW0ukjrxHKM2ypsI1e5INLvUG03g/kc/E8eXziM8yDssbHSssa1V6OmG
2eEaER8DNT4gw5FiREUVizD9D5xJ/EaZON/MOABlAx8DHkBhAccPqEpmak9x0khBZJhsP6s/m17g
w1RM7lpqLzWcCphKyI41OvVrAnd4d5V23JXEjtIkH5cF66Cfa9OZb1Hwdn+Q9tJeaDU2kazbaBAz
1BPQxsHNcu7Dr9k8nQ2NW0Ovd+Maj0r7W9gMWirJ0tqaXqAUe59pq3tum5+36bN4DfdIl0xfo0+o
cIGxjpx+d0gIur1Bf+O1ZpRZDZ9BpU4wONmwq2Is0/O9b5H1EtLPiy+V8ohBZQgcGni3t6YlCaOE
DzkH82+62+5/IM3HPlcgLFBh3XcyR1ALAGuG2sTDp3tuCO64V2FehO8Zo/FEd+nLJLRzjrfzUyjw
TdUy/TVHLKKs4pjRTm05YU/mWbPbs7QgXxyesnADppWQrNzq9EdIfrrfvamlJ8ptLAsKevdwBN7T
XAvSM6LKFYTjOWthfNovi5WavYi943ED+GlZhrZNyL+EQu2LhxKKEEBmK8gJH6Q+KjBgAX3SA8e8
OUaY6sAG8JGVi1HGIZjVB2/MI1tDkLps4waK/W1cnl2RuK2Dvt7Zl8lTw+gy2Y4ryvSViPw8dl4F
ngjV+YGrl7x6voK+sWbN4R8Z+N/qiZw/j8axzpnsKEJzJ0hsCUbHKnp1J2sPsiHpeS1KTQ16E8+Z
Ea/fOxFdRAkdWxjWxlOrUp1xR1OEX+itjX8O0VKkB9DX3NsU+Nq8vT6J09FBOMU/19gDMt5NP2W3
BRqaNuq8pIfWFWllRHbP2aZ637NCUAa4NS0UcP9EY7b0KEcB7zNB6ohzDbUF5DcIGHrrOwctsN2o
4JwM8u4JiFSYYJJnZnnCOwpAIFGIneOPLl3DAZHHyiMRe5cZQSoQI1k6Lt3xXZTyut8P0C/qqHnf
K2phNHxUJ+pD+7F6AvVkvvWrwgjd+dYAy7pvHKukD/xOwR8/IeNaxXSytcPmFv27nVlyxWwPlft/
GsnK3WZcUmIcjAB6PiZtjTWjSXJUPrJ8v6P+1UX+47WbkEVWtgyjEdcZrJVXMVqvmDUSHo6C5C9b
JhDM/7MNaTm8ykTtuvgeXz+X4ixcm+EI9WiYpfuPiq0H277X6+IrLCCmJha9nZILSebzQqsSSp41
YV3e1lqX/dS47WXXqTNToeED4kGh+1WJxSK81F+SU9H9QNqHJMil9Wp4E0R5Tzi6qzSG/CNRjanX
L3VemWr6nUZxxf2+EmDtLZZJYwvmbFMjMp4+HSszDJElR02jvhphWOpkGCUuvMRMqJXlsFdoBbgq
Gkbi922KcVLRqDRGtLxZCKtdkFiwsJV7YBketlX8M9/FdbSXnNemhIfqU9Ti/zf2eMckT6Si4Hvl
mFj/NJ//hE0Q1AV05B68XPfiGILdVh7vpvxY5AHAFrn/SrOiub+PjtQXnhfUHZAUrzBxdNzBcAd7
kf3QzTYs/PABj6kocKMiDzs4H0ZfZPsG3SXtCPbEMD8LCZP/oN/OsS7VBf3ZlE1YSvRiiuzD58nQ
Aohw/ak6Z+udVx9XQN2XGwqT90t/LvBUZnX1MV7zb8A77nGT6Kq7Kq3WjmwPpIIGjMfw7bU7aWhF
8sz1IB/fOyZ2J2ynyzP29H9skgjp4Sn/LIMLclA6TkhvMdc2MlAF0XZm2BYSYBIKF1jQzTmVS4dq
6wAXAuljH5Q9JSY1aEz7rfNsAyWiJdVnSoKmOGjpCUAM927IeOBDVWBWAugMUjZMok7PR2lEASZc
AXHymycwvzFZndDmgkH8cMeQvrElPc1v4dRNe5owXJ8pa5IxqCUwyj8pxuA+vSg51XVlxuSAIiX0
HoZBoinhDLfNLdhQH2E+UkNhU47wy4WmhJZ3eZgfW602JKdVZL81FEtvBLlF/8O/L+NU5x5tm5I+
X++QF9A5mDpGD/sT8QhTVP7vkXFaq8jMXMiVTSKovY2925Ym8qc6F2vAMvusS7NBc3wzGA+AKdWS
+ZQva8XiX0uNLzjTnd4WlCnzj094fnggemhSNgTE1hXskMp3yF/4ZsOZvJO1oQMDCZdyyjZY46kr
zMGtfyoI+ktEjfiHdXxEPbNR+X3aAl9Teny9yyPPn07+N6QlZR1nDUmIAyDIZnztUM+sAUF+fpPk
dRvBKE0nUS6iEZ5idu/a3SQ1sLGYhRDxk31nHdizZKa6PNoEnypLRYKZRm2TvritP930CvTtWoxu
/Gv1KjLObslAJt+TvlP9fH+t70xtt9woiwZSCsBcxLg20a7jq6pMRHnfACSbAw1ridAVkwLoHXcB
oXDSHjTHjbwqDRk4ZydDw5SAKOeivchghhco4rNfXAGhbFn7ZO/OG5wE+vAYujcNzF4vyx0/ieLe
qAarVZ6sBsmNbFh0SdGcrky8WI2tAqOfNfX5ksSsXpZl4HRyOG2VActH0nUKqxoNPd7nztoH6E6/
4eAtkOvNSup62fYVUEeRX5YeveOStIgHVomLi6scPznviIwdvPOvsyvqFpv8mwOzCsH/pPOnZ8DO
+/3J56acBoC+zrqOLCTK5SdOO1hfAsyXvqbQqo+3Rm4bO2Wir8BgvzfjSfDOGHBaO3/HHxKP8PRN
w7iDrlOxp1DNtR30ofYrUKt3d5uftODke+1qHwKp+fkH89IZ+bTOApurST/rxKM4TcRDs1pwXQaV
zLHsxplNJ+4/t4tJDuctLUOyIHh0S5Q68JHKMxKW1pmNEWcPjC8uRvz2jg2AIy0drCcttqV8Qr7l
LDNHkXjIw31+zqKefTTNfFTGfGBfMhfqbKGzLzI/swdSDh5Jk1u1NKDjWvOLV0us9grjz5arNdeC
HyIyzLI/ez26HMZA/qj43Z8kwQ1hfjd560bsdsMcIhIGHEb8fihxu3qhHnuKTw/X39f1Bgt1Ohh6
HZcxeCXYVk3pM1GGrnri47PRFMpV8mv7/GIA7WdPMGNE7aHpTMBk/y92wHbjsFJNL0ciyOXYtsuZ
ae8fqdWh+/us21yr6AwSWLqmYCyF7tntk4ffjoNnKzQC9zTcXeSuNyu3/thjimHIgXrW8myflPpK
Fktl1++iG4EIqQ+oni/O73AU8xCyZw0fQMInPxz6Tfz0OaLZxH8tZzEekmiZP7+l8403Q4yPmQ7T
+qV3breugtHRM9BgOCYGhk21BPUEDmdgR/bV2LE6pPK5BmU5plIcARmSoKaLVNpNcU2M1d0a8+eh
OE1bm5p49zUrKVc1Nd0a4zyW5YyVpI+VkbesBvk1pqbzYNeMI+Tqh6beMx/gQo/P8I14CxlQxLcZ
ZgcLXQvN4v9Eni3delWgjnJBZwBt3ZLLxmqX5mzyRiDTPBYL4KKPjxuOfMbxbD1P2HX/31nTQ2q9
BhHdunVtNs2EU4wdLm5j6G3bZik6bzkQYvQyz3J+bMNI0Y2jgU4dZPGe6XO8abaU4097gHHLjwdO
GX9FnSLAjP5GliYiwAc8iGpOUErbHKFgGkYqRrc4WdJ1H3D3S3Q2RV2a2DEpM30PxGqnvy9bs86p
QY608OKsEr5dEKqjrlFPcIfLR9o8Tscn7LlHpwI5vb1HJLQVmMxE93+TZjRRFtl69TmHApyR6KY8
CmtJfOe879YDXZXEkwedME6m2rMbHdkgER5avNQSX3iqRL3+aJEJs6vZQxgKDmYZC1oOtn5L/mTy
XHzrLhN2sxkFxNNcQPR4rLagEf3jKHcWjMPbP9HrDhHQ4K1H8+0uA2C5wf+OaJCvytTbmYq0KVxy
DodPTRSuMPeV9d1/nPjJmzYIh6ub/V0GP+YGBGNqwu/iXBNgZ4S31jEBaeB8VS15szIpqP0sigmI
HoqJQ+7UYiL1bVJyYWT+gl1aRv6M9L5nNKTOH+EQbSNf0wZWbtNpOg5uGgt8kzGvI+s0et+6dVKa
Mj4H0P6ITAofpXJg1LjOnf2yuuCbZBR6tb4OB1hQ/6nYr5fltDWP1Ia0Dlb4TS84q/unAawg1zHN
A0b62UEj7er5wZFZOGbr+plUt5oV8YfYQXVVY4wq1T4FlIxJrXesMTrjVSpvxIitkFAfbHdXRxtl
tap0c0XleT4R4vlpxFM0BdE6JTz7oH0qbqa+l3f/kKEATuhBpQob6fEdzwSk85kq2foBtvuiWgIp
i9M7WvO/sdb+n7pCb1Ebh7SazlORvSdCOTNofYLphWy62OELejkZrMElf3luQZK528tnz6kUv0Iu
msCMuGgvAvtGnmhtR6xX80AdU/YzvAeeOP9BR54VyR6HJoqtqADzBvk1QD47qEUZ+bguVRBuV9e5
BzZ7Lfv6j/0JQQQznMYVcTZDZTDr+AmKNJxeURZ3oTQva87rLONK0H+SI/oiAMiaYf2CRiJ9WZEt
g8w41NAkChwjfGs6iquZNmhP6zE1Bg8dpJAJfZmnsbyOVz3c11+26Ahzyk8tAOKBsBKXFch4XErU
cVirrMkPP6SuQuE2SNXhXk+YID2sxOBZZxzSGJEUHWjuC2sxZVHDraHb9nHQuYLqorSO3Y3WTD4p
XigN/Ua6TypQM8po0hmZ5BSrOxiNxxuoQoLzfWXjIv9MP7qhYjL2xgFkbU4LhjJgfwy7Be0CE91X
pYZYQ4WCU43oVPfKQn48ca3axnh0kx1OtdZcgZUVhvajKqd456+QhxpA7pa0mIDPT/85sxh+lfQ6
DBwETnnDkz9Dzv1VVykwaWqQdVAsuOeo8Ei7Spp2G8IZCs1qawx5Zx9EKYyhftNcxswkQVfzfdlW
TGMXlrww8shKCuR/OePkH9E5w79l1DatNWFpRqLeAjL62WHklWDpGjKN48gx8yZRLi96sP0DbDRA
B1wmJ9BStsyozpRXDnl9Byr7X4gY/hQFbqTxu4N9doDQKHYnJ7IJPvjEFoCv8oFCauKIDOX1VcIE
kqIKC4WyT9LeDCjiiykeOK6FSdR3oamS3rKJijoPQyrZFmG3yKv3kfIkTsp4D3Sa/ShfKNVf200A
/wjmXURgqfuSG2Te8vAZ1F+Ev38Lf8WBoZAYgwxoL31T/E98s+0bDV147Md/XX0Xn0iuQxmcT1c1
2AAey/UkMVRjoM+KkPjR0oSNV6hocYeAgY6QVtWByOvegNYG8qB/gwFx6bn/DflPcaRbA/cD3CeV
spLFNdA20QRnhgsKN8Z/jc0PTkJYb/a4xk26nfxrC7zth0mYjjJtYCpqK2daY4K8L/HDQCL2kOuW
z7TkJBd5HgZn858xxStzxrClUz3nLtCx1eBemdRy6yc3WPF5Wq5wSXHOcEkr1sZo4+UVUvxIoZXD
10p9dGxfbIO99bBel7dscxys7Je2waqBBa3zajNWRcY/Q7fPZO9Ad5AiCrUotpheJ0HijkrD9XZG
fabCiOH4Rhc6BEAeFjz4Kjkumsj10yytv50UnPUnjPAh9sOT5D/mmRvBUBmJ3yDkd4drhljP5zsV
Fp2tnbfy7w4hsYuac33uZPPTyLEKn9IzM2kaiiO33v61KAn5pLEQL5L8dZlJnGjXEDCK3TnqMOEd
GuEnsg10oUfZFmXubCmkX0O3PKFpa69oBnuVUBcTkZghtfVWjjKLQvfKxxqU2UW35NnollMOweb2
ZatnBiOuNL4s+lClpO6XKzVS9cuo4WCV0pv4zSdcK3qLGCfLdzRgrxLiDcUUVgbEBm+yk3UpHy27
aObLfoQXNzPvR7Qw7R3f1J9AHI5eD/4cPwEQxs1HBodtHtybdcfbs3X7oyJqGFMuu5aVsGx1ePCu
S+JPQpO3bT73U0rHm6PW9NT7HnYVqz9YEQkqnbHpGWP7q6KgPhUm5qQiRn8BiULLjC2MVz938UjX
NTr4kmjVUsGDFIp78H8Z8tszOrwmOxffM9JrDtsbP3AF+kG+0y2O0mun78+Ayq4rqNCKgfYv49qQ
ZxWBHX7b0LjDmZJYVcghvOyD82qmKqkC5CxxgiCDV++CryZ3EyFd3U3MSJ5Y1lDZY/lRVr3SUTYP
c4DOSbcf3JRULl8OO/+M+oZnrR7emuiorprWHff7Lzhn+VrhR9H3YX0fswddF0AS646B/4mP1lDR
+rUrdgNc187JlNzDtjknz7vMr9jv0NpwVib/U5N8yRpK0Ge4V4xurxTR2e0w1HMw4y8LDHB9SiBS
Ux5C9WGcBadTg+6sHbrZFA9MhOH++NASc4MzYSylql4URJet74CKxnaK5z1FqB6Fmjm9hqcli0YG
1TplBt4BlhtJsEC/tTw9UywWFqWqZFBHdY6tv7bFIDBYak8dzLTTpfZA8v0HrePBxeQeSWsM/lVW
ZAavlTX6ViKdCnIoj7O3gBrP1DgrRAghjmWSkdEN4SyndToW7kng2h29nXxEggXF7ivnpmuytVbj
QrcnEGvcoKDLyTXlYTk4wvR0XuBn1WCad2e5NncP5TPG/seFCcmGh3HpPsPr6G4QC5ZXBBS78hSA
xjDk5WPnFCelkwGJwp2LrrLlpaWVEmpNPpFd0Ml89onZgwgzS3PK2/MVKOSJqsvvoGbzoHkc0sA3
xuRGumYl0KuzE5A9EL7ip0SLu1V+aATRC8XM7hoSKg0bCDJayzdKvKOTc61O1immKh9LjaNaHT+b
rTKfWXfG/0X2gz5mPFr1Gmok3Y8VxT01coToZh2ilYPL/ya2FOhdlDN3hVs0LzsnAagg9aYmskIT
q6vkzOYxkaccRmID+QEtLb9Lt9IH3lzX9RYNvKOLHOPT/MAeDaZBNxpDHjDuunH4GaGATWC6PAjv
EHPRH8xxBAQoPn8jeP4beuYbG5gb8GVAF8AiV5+Stj9Capw3KAdmlC5iVSbUJCy1wpNvIzcjIsMt
coHlKVnilpsS5MTk+lYBTA1pKoRu8InZ2ROt9G7QN16KBJ4G4oMvDEmJmhGw67MzNHvgQaQkyP1S
bGd44lx2DFnGty0t252VKHFWVlZSIq+S7gOWCbqF8OJUlgG266YXEEwyCnoI2CoIEvjyltT9THti
vbQm3G9wAJlqBn4DReyZEzVL/+hlHFijYZ5Vf12QHHdm7h9pk/7WOhxRlap1Nig0xYZC8LeKQgIB
WMorNtntmgVc/XRtPZ6WRFwMpzQidmRibwcrUYYuxpOPLzgFFOm1REwLKpudRHVjcMaKDivQiU0e
PVXCLIukJJrVAS1pZi3oX/qOU/0FdibUpV/76Mg1oqGZQj1Z/gc4NZ3BrsR8ckw4JiA2hV+cguIM
XWlDJrcNoLydxBJy4GC3T7/d5mEuO737b/IZhHEG6cPSjdlFykprGxnYInB3f9bnwUa4sKoNQnXn
mOOsdK7043sOJ0N6y9qL2GMyR3LRVjsyzYy5BRpbxFv+zjMbBY+amAqvtLuZxfUIBNjW48BwtnHu
dOCameZG+ohPBisJ3aNT4KN1M2w6zsumjbrtQSjxe+sMJss/qZvbXkh+sctgDZaEfXjmFEvve4d4
PzkiUwSV1zg+k1Ruk7JP8jwNdoqT0gVdFUTvr7Yco/J1ZwaOOY1z5Lw/PtDvxt9y/0NChQcpBVVV
lpUFmL+wabL8Cpx3+LBlVrcyPkQ38woeeYR4D0xoBGHe8Q56RhlZbQQ3hVR5hCr4bURu3Ke2pOjX
brNGdZ3Sr8kN2ANqVZMTlMRt9BDWyFj2KVOwcL488/YWg6u+342GpREmdgZUCKBAD7mjdphXEO5T
IaNpMmt+WpQqARsh5dOojqZordy7hUMqvCxCUXPuYNPz9CycnO/6uRKsLRBIkLY7XZ+MU7p9ajXl
G8KQ7F8E6lkL8MBZ0ptyv8HUSQ6nw3/G8cT90BY63fNMLzm9vOK0egNMllfHqq9bcbSuKcn3TRO1
xbi55PJApwIeCI5mX/RgpaGmAgsGhcJbZU0LStH0OL60lEjGktLUwdvX9PS3sN3vGMP4agdoaMID
A1Sw0mFBqud2SS/IhtZjx+0WOoDu4YVzXkutzjQ406BZadcm65QZcJbpEKWurxFOT/Dnczcv3CiM
ZTmOGgUkqxyzxqQseRw/15aGCKWYcZ6lloSDtHhtb9gsAV6S2PBXt/U4RcRbsn2Fpigb4u2j3rCG
bllcF2bsEwPDQ4nraehmNN9fbxDZdFrExF1GlmSe8lL9F+PPGyz73uMHHgIKrX56RZKrOpUsyhs3
Hrr9cT7qCGDp1BNAUW17Gh2cug7kAz7i5fZgrnGoJs4WHNqUqOR9xn+5vCOu68+TPuHsxYgECZVy
XvoexiIHO/4BJm8kl5XGvXw4hQpR94G9t3jdMzdrJTkHwg0EHWcrMjygsJ3+tzz5ZxwUu12niSkm
26lvEx3F8owI1rIIs6eudEt5siHDls+uCvqKcPpc1RTckoaqBwTBavXnUU7pQIu8D/+GIPuVNlDx
kVpS22eYNRAj0Y2/YNULQH83Nvjsrhsx6Vo4SUW0C5TeIy3OmJhgLwD7n2v5VYmzMacwIvRfEt4G
nK9v9Z++07/IH4/NV7dSXCwEvmcx83TNukOFvWzYZHMtDjZ6VYunBRuutVdjnFiBB8BG7Ed36nhv
yEruxsA5g4wvGpH2SoKjXUNptZ9He9uHrC+MoqXJ5rXDF35YV4rYGqAiqSme3Cc4eVa1xTlcqVHW
atH3eu0xELheVavftyQkkJgA1OyT24FsY29DEgk/tFMrv7ehXmWyo6JPw9BGrXNfqriIZ86oKquT
pbm+FVxmTldTl53lh+opY/Jf9JvfmjRhjuhnolUHUcdyHqfmMUGMqm0nTBYPjdroHk/cDUKbVfFo
TZIvymiKfn0C67toiP8EPjOMPhBQ98LeafhnmAMVDkLKo+XLSOXoqybikugQZVR3vUKTQyNPmi/T
kXoE2ure92hRoO92Z29XwplZdpGJgk7UrDyo3lD5zYQA7Sh/83JUS++idDf99D8x1Zh2nRMoCmTV
9er/eqvV/oEMMqbr7p6VgAIBNTTmSJOyPHyURxex030rcpvNiqcl6rrXsX4z8x+gVUX4dkGkfE/n
IB1v4mpC5Sv1LdMlj5c92Lktothq+8FbwfzCzmv28I3/V/FuPhsaVwaP9In9uSk9y8n/oF9+okd+
CKF6cvkuwzRdhmpOI3DDNY9zOX/Xs0zlfzaIKokBmzgWCYBxCLELLbzRM0DBR/fW7U0WWYaRL817
XSpqAKPE5egic3jf6eJ6CLegw5RwLLs1WPiUUWJmoyqQGgL4ejI0Gkk4NLCeEPVt9OEarhiu7FWH
NFSUKlBnzk6dnN8tnygJYH3vgvNXGpRM4BnFxtCwltzdr/GdVFiMudtH52KKRDVFYkRXqmQBZz51
kALOxeJdErsv8KujcJS5tZVcBPj/Ye2YIpv4AsyJzCtLK26gTwrkunPkPtM5vWTuDBYiAsY4FyuI
utqH/F70mMTtKd+614yIwX9sbm5FOPnUDz/NYm3owvtLoL5oPP+GCbB7ZgRCp+Acw7IphdJaDiKw
nUC8InqTIDIhA0iSd1/aTkPXZF4mUX1DXvIdT+jMHFAUiEP2PUATRYb1jpOolGAfZHgoZOxTVJw+
PSt28s0/wO7lpIKVRnFiEk4KK48uoJ5OrbNBvC5i6MMjApuTnKEUKDPSatjWx6pCpxGkj7Gq8g6A
/6IXIhh6lkyE/n8HV3QWCuuP/DkSYKo6BBLPsI4nU0+n6H8EZn3rBa1snNKTqbOL7MtNplfXotIY
77O/uRyDUruFz9EgoU22vsCymFFF2h0LqumvCd+y1jqezeUWjWJe0obhaqgnQBQFlQ4AJ+B9K8C0
7VudkgFol7tcplrMSGCmSMzwkDo7AGcwZPjH/HeLSIJ5Q01UDWIYXJeQupXkFrVQH+liLnUhhrWX
QAEY6g/ujw2Y5h0JZjYdgm1VX1WTpz3moi8aHaDWJ5TnvSfaYJ7H3HYcp/tx31Qbu5SQkSFYSagK
YcaJ/C5gWFlxOAwPcatu4E8ufauhUAQF4E8RVnl0irceqVsr16wd703i7u3+GYIh2PJVbSFMM0QE
/54b1VRBsEQhvEVP5bjqafVgRaabqdhuiKAfhP0SohM0s4CHqBQ/E+tmfZMwNXSSzGNXUj1x/wI1
nEIl18XLR7PqIca0wwMSe6NYprxfBWsdlvFm3fFLm3pqupNnq/zDFUta5sF0UQw5rdwvcNFSp+nO
+yOcUoW+LcfNouLoYPDYpVTq9LOM65KIOPwy9Z8XO2Ap3eUPjTG7+eVnBLtumHndBXU3fMm0sg3P
cTHGLZbBvL/0+k7Dz3/nPZKZ7nWNEZx3Q8NAqQcnEF7RtVidfT+COWd7ow/NBt+r1SCYfp6mnaYO
FEQ5BP6nOpY2h9Cd9P12vypdd+yAf0vp24oTpMF+ji82U5rOVr/eomfaPCsF4IBfpiePi86ZLmEY
/BSrMDzrqV+My3Wvr7acJNlAI2LJX4EqDTiAgC0/13o+qN77mMDHV5XRz0wMEQ668G30rIZbQFon
hmnz1kL99FLA4UtWxg0dR3oiVpfQklOookJQirE8MET9VpZQRbgGGk7V9tcFOuGkMGeIG5H2Q8RY
RI0/CMqtxRww89nygyE1xBkDiSzRnYMIkO3MLKTGyh2SupJfAVPfQOKJdCs7faHd1nRkXPqDaQRw
yeWByPjcFybDtCNgThUZo2GWaF2vmKZv+Shw8A6uGT3ESz2XQpINdr0rFrtkOA7FH4qA03irobWy
qTFvdsaYE/ugWaJmCQgkqlk9qgXlHK09HobN/2G9e43Qjv+pq3VtTcCoWLzMQpTXG7DwpdNMjw8D
0Nj2gUzmjklzOeL7JJ+Yrs0yRM09KsR09OTvz+sUlovcyroC4DkBgeJkYLa0plzFWUB091Y0bryW
JIrOsVxENshMs+tX/nu5DVYWPovL0kfSMdJUGNGbeQldUlUB3vuqb/syCwKfBL22mdl20szkkQwF
CPtFzJtMpDDTKqzidKgM8fqMsX955IZCK4GxVxqBmI8bMseT+HaMAZDitv1FbwtPAYTMUJ5wxttg
WZDXWOhIiY4CiqHAds6mBNvD0U6uo8+LFfT3eTfDaOl5cGJ1jBPd8vaBnh5HxhIHTb+QZv86XN7K
iinfOLR6hyuDeX60JeoUMNhbdTX3E805NmrpJcxtc8hB4YRG4oC/icwqvuU1RycFM+6Ey7I5Nv8l
BBRvWcabZxANP1IsD4oP6RujTMv83syCYOjC2WuQFVWs80OmSpN9jXf+SFtDnww7RK5vNWUYnKkZ
lHfC/pWI7NM6O7U7HY9GGC/F2sLqtBdr4wutqo2aoifDOXMT4DWZlMBjZiotnNsxwDr6y/yRs84E
QM/5EmSM12acaS0tKJJcPcEe+3XgKgMP3ErvcuuM+1n6XKaDP9+ldllObUZPJaX1h3SjA5WRIW0z
OaAiwilnbYlULi4EgnPuQq2BpZicHpCS8RP8NO/3HwojzGR3qxNedi3yMgAdXFvyaBsopWf6R1LS
GQIyhkeSNTleAWjQKZdXnFl8HCDu86yW1cGEPKenGifiwawI0m/XpEmuDziU41Xpdplsg9l2kJqh
cJOz1wexLkU/tllKtBxMhGaHoGAFWXLOvcueoPfDFeMZ77wT2JdF+Ikz0ehhvdG4lPJODe0NpupO
PS2fwgn/Lb2Dmd0iX27xKKKRk6twxhynL4cFH8ygOpJmw8AMfii6dqhLY7hJEI5r4xBy2Z1eEutv
zXpN2FimGLebAImjp4grXR4ppHPcz+EYbMXCT5mXtoj4S0F/UtFYh0XyZ3EcAvdMapU6mr2w/eej
C0WK7UgfT9Dk5jU3WcLnjXtYe7M6sQsVxiuBgpHDKdnbjggIEPD+EjefDcnA9Dnd274j417qnae4
PmQ/nlnUjei86YwxbPDmnu1qq/n38kjm5AFq8sM+y3EwhMhWXFguZj6ZUXjGR9QEt02jKJMCMKNt
fM0+FO0pH2EcoPzpZ6a0NmnV1kl3AE4+TwT3IhQ7Xv4K+ZPoznYmaIgxut0Y69WhkZXx12XAaCUD
oMPgNeOQ6y24nh8kiD8dr1wTKneYpht+7hRvK9x2zXNgX98/erO7IWiBhZ7CkyStAWd/VpSng/Xh
rk2UR5yU4G/PK0q1ZB7IQdzjL6fNG6rAzOfI1cObwQ69fYiaOod1sjm8zs/wJV+/RuHz/udx8dnh
YiPtLA8nckwblH4b8RkkMHytm6jjxhxrII0zok/M93j8pP/8oaleNFOH+b19Qv8FnnX7Wu1PR27s
R75bYidv+i8U2tTiO/DwFxwWCarSUjj+wG9bH/tHTFztndeNB2ntI2mA66bCB08gGbwowRwvHz3S
vJnyJyByPnnX0iImJIML4ya/NQesAa62+wTxDbPX40hzfBxhbs49m6HZNaAeB2pG310qH0W68rP2
aFaj2GCOUuxmis+rYK3eyI2lWYLIkb/BEYDpsNnR8A2AGiYINZunjIfd0GCGZ93GUarqoQrO32uK
zWJlRKAgwqJdu9CGdozepV8swoSn0j4Jz581NiG76WqXapeHODJeCBlBlDwbJBmNtz+WonLQ2xFp
Yd50bSsg4XSU0Pc2QFfB631A8fYzCiVSurvJDTTIEUIMUWjXUu0x3qmRgDTuSVgTNMOLIwft/9f5
LT50CQyEIrJDWJ0cSun2GBWZu7NacZt06iDep7SH8nxp/k6/pT9H9JNdDS2qHRRM1qVMM+me05Eh
7RN3ao5E7UqUWQqlqiePcfbgcOR7YjrKY6JryPuXyDHmupBg0G5YSNQgr6H6WoZ67zSSZf0pJVSb
xbEUM8t+6nol7Q6REUQfl7FPYhx+F+GR6E11aMK4NXm62Zm+4pr3tAri5635/xg0Lyl8Y8//4gO1
bSHqwbqGNFajlDKOZrDt1wOHZnYVb3sznVscIm/12ePahXtjGK616Rpu5SUc97CskL9fMx8MsDnn
uYmLFKPMGutHdGbbSbl1lZmEzhzdFfEtPbj4T99FmYLIZNfalbolQBuvc5hTGgZBU3z6SbCeIphR
0V+MUzxEnHhqjLG2BmrH2JIBfTXqf/AufHj5YQDqKEgt0IR7syQ0BJdRfG3yIZkcwXL749TFZOSI
kl8PKd4YOVBREZJiguhCuWCOsZb9t9kel+ocT1xhkxgY9ohfxlYxMtZ7NXU0E6vloQhm+s9s9v1H
yXQY2GhsXydqdudYRV2kjztjCbHDDeD3GMgcyApU95TO5sKs98pfeVKfbbz3hUncgWMCLuZ6PnlO
6KG1K3YknSq8Bwbkql1rRiOIRW5AzP3VTJj3puEDZd2OdbKQrtGdBwgPsk+ohyx4yEGI9d7J/Cq8
weDD/QNHF/2OOhXGZ2VoYrUdEOoCVIi1sOYq3iJj1dvCP+jEL1vChDtMpMmQmKLnUCytHjkKHqrc
kr2F2qKKF96yXjW+vK8+mWVy0dtjz6MQYHV7VGMlacFez+7DfWWzCH2BXXnJNkYdjp36Ys0s4wzJ
r2I+xdjnIrwT9nt4JijBVRRTsnpb/rOs6RuKAXVyq8eTwa/rDqNozHMkq5MLy0RZip00ixG9mfLC
BJ0/CXhtLqHL2JswwhuBLCsrQdxaHSDTjMgNqcCPfoXz7w+QcxL8Co7gdZzryMWMCmIwHWkfXBQf
UrHmUZRxZdn7qM+c+Ps4S9wpp8w9HyCcZgq8+jMmezRZ4rQpwydh0vpZiy1rOhL07WN9N3rhdK1K
yeEIN7xaDPaeKT3mkToDg7oo7ynR/N42OyfX+kC83+xCUaR9qhnp6fXORnOuOyDdcFW0SAQfZKB4
OmoaHSkTXBzu4UhTLR5W6i3LYudNKiCC/0KaD80kj3N/bgOshO7AUbg7d4HAiUDkmUcd2x50unr/
qOuyeY58pcyO/vtf9WIRhudRDbSjsVhDHXXxKNbbHnaw6HEdXhtDcONo5g3C2YLHXgd4bASonruI
hZ7W8zHaOUUdD9kIiFnyGMxBVmEmQdgV6Tpg+M5rnZzIHXVyGsQq0tavJUpJf+7NKAEwWGVs2kAp
RPI8s3P+37MTmUmDwPH3uhMhDMJbePSGcFYOY1mZMPJu3pRPpwrPbunbhvsk+xYNpNE9C+s3++rl
zR1GY0azOR3KCHhS38ps3vW6s2VsuDOA4P4AyMNZ6ZUYTPSEfLSnUA8R10YFoC6dLSMl5xfW21Pn
j84HG+Ds0CQ4aEzhKp4ExDDiTu2AnvFz0x6a42ED2dIwdyadrLP/omhqksqRHLnP0ppju7Md6Q9d
jCMGtphFDxGbEF7llmjqIMF6lKvbOK/VR/l/FMxUrnQMk1QrdpfyhyXXI2DryCgcW5OtQGWc1oy2
1XgmDU+zpCTaIIgWz996K8ipFNpA+f+WAITYQ3leh6l2NkJHkFARsa8Dkp91prEjwME1awSzGD+T
SF7q5o4ISsczEFfdAFnu5j5SWeh2i1kzGzdi9S9E0hQJXaVXq1PpJEYw6jPM0OAAX7oJCclyKGQf
oylQw9UFzq4W2PAOnwTlqCO6HggfJTxrTvY3qu2vlhuh5ZRkzCffFUwF3VTbW9jfZNLoG+xQKRea
u2G6CZD9E0JtB0m4MLNVuWaZnwbMK6sK3EzxPMlhMk0UjFUD4eK+C742+gWgqYolUHlYkZq2duMC
LXKL9brozD23r98rg9AVlzSQSz8oXyyjBo2cpQ+ZUGoIJq44MxvUVldZElnHMXcTfEgg+bxdixrm
+g0lzb4/1NbwQ+XuFWH3g4NpVt7cS6yILJ19JDODz7HeMlrfey/6qraC2aIThkyo7MQda8yLllYu
89P+AcryzcoYvpmw/k3CU1uJloQccQlTMgzz9Q6hDdAXsaU36n3UCboT/T+gTuvyJTii3cY11dys
Tpeb+MTMPad5kXjyLTGW4EX1JZlxW8pk82TLfSCzbVBstPfZTnVR6OpMFOZOuSqnQmaEcxuBUVik
tBD7I8ln9ImRl0grXVlSzl+O0WdV2a1kaLQ6l6+ApQCu0XHj03ofBylv/XbwIiRT85RWsI6aEzBV
DeEuNilGs08oa53o5UGrFx5FHi6een2QGpAqVGS1GSqMT911B8fvoUZszijhFqgYwNaRprlhpX62
oArDwBPpat7IcekErkem+bkaJT2o11RJROuX/hS9CVlKuAlXZlEFiVakOpMai59Q9+XmWN3plgok
At8JMVMWaB99/2oQgzS6lMbowj/RaUJ1k3u/x6b4Uo5jO5O6FpFMBRuVGAYezW/eG0Dpz88AXabo
myz/pbQzgt2sICizD++P21nsM6ZcOoZU+HQ6nTiFJGkiU6SK3sc8FgR3m/YKDOxYxHLAj7AJ/vpo
vyMzzyzWdbYEtRbWQXf0t6aNPa9A0O12xK76z5ZjvjCJVxAaJSXg1kTGGwb5O5VikPmixDgvUlSb
zN5AOZl9V+hnH07u9ou14h6Y/+qCCNYWQpbc8RmnOnvYerGu3WyXC1FoeNvvWA8mUWyzVY2UtyuC
cbtc61rzwy8LtEWv+FTdH9pijjHJPDzPccx3CknGIkGseVlrXpSFGv/8UmpXmqI/dS3wU69UinZ6
gRTKKTpYyPyfeRbzI5JVZOIzlXa2k2dKFx7Wo56Ul1XMfeg6hlQL3wXX4yM9qtk1a0IXr9e+OiDs
4223SAeVK+VSKSb0DO4kZU+WG3aFPtkYNxRuAa8NnkzbotHjYsN8Wfk92wa5873wD3HjT70sS+ST
LSaZJrUOjAqYImNF0U+cIzty5/wBbjDp3b3BdziO8R9ozA04dtYImPC28SlsID4w9Gnx6FWY/uB9
A10PyFfbRFlMj2qqUbguGCHOJVwF8f3yfq9znrpIhs7ZmrugpIwyXlW4pQrkW4tNaROsuoOfUjFX
vpf0PySAH/pTb7vwuq81UNv9iVLSWMeWlKbw7L5lAq5iZOYb7yY9q+UmbtCs3oVxMDRmDIF6DHmM
Jb0spBKG3Wwea6+jBdYB3g82LpJutL5mA+D8BiPp1WMf7OaLwmU+FyNp3B+N50Mdo/P772K9Se9f
pVyvzO/sw25NekEh+QASYMFx1HtjRR4K4teO1aLgPfeAeiMg3EHVRdZkoxPKEcq23g+6Qm/imw0M
OcwV90wL5fLfi5STiRE0cPf9k+JGVD8b5b4z/IqHfeVlY4Pn/fQWElTQaxknFdee116LY8WGm0cw
IULtMTfUTaET/U/JdUez+hdXckDIWE8dcYUpa6cwqkGeFh6XdINyQUVWFrR26ECfz5TTIC29jDo9
DV7gd0XSwQPZ78mG7/SEnnnqgGLRVOFylOayIGsumi03SGC/ETUa1CX/j49KpQeIeSPcMu7SQ8Er
nooi1ZKbIU3Ns28K5KPPB/deQ1N8sxA2nS1Z3mnn+IvMt7JGnOxyFMPGb2Zrdbt77/3XHOHpGGln
wfpZuy18i2DVQrluptLtRq5uMHPzbIrOiTZu/m28/8gi+aw1iDe/sV5vAO6T3yVXUu0ngHum/gN8
UZV/M/XQkHStkWDDoGJiSgTplzhGpGkuft9wcJfUuIe4wxKctkAc0UQ76JGTbIgIR7rh75nHua/T
Lh+KNcDtdFB+MyoX7R/89SR5fu+rEUCo9sDOAK/MWcZAOXAEE2gBqnFNI1VGePeCjM9Y7ivbh+aX
oA3wJg+PgCsGYG7xKTVUvHYHGTi6LBM+fA5HoUzqKYqBltLxLPstR74giFenicPp+6fCtuyXs2Ny
70whWyL6irwB0dH+ziiOmSNdrrAN6soPrGC5S9Sevp/mIgHczxHAyqSfVYWd7BLiyAglRqWmyV7t
Ri+a/bSmK13VhqOST4uPvFDTDOfM/8XxLUGs/3JJtNrj/oUXQAj3tzD9+orcNgWsaD8zybTl2kyS
yGULOf84Rm2P2sLVTlFp9MXnnWMz3wQKPM7dr922koqOfe3CnKotKDQ6ebnQF3Q2D6xJHyD+5Aha
Vu56jk69hvg37N+6NBWKq2kC8vm4FQXYwsqSFjzwdf5slPr8T+loqZx4bCzefwCdHt8BsYekW6n8
2/dTsYBZ+wbouR7l7uAyYIbCc7TalYxkwI/vjeHps8w2BNsdpXtOJIPezIt3mV9e0jhYMUA0Ft73
FJ4hth44XpSIl/+CWXNjp9024dlAJzN8IRWhbZJzXDWmarxZiJpFnZZvd0WqpVS93d1WgAthcXT0
4CN2MyIHxN6GBX9r6dVegYhO+bpfAFCZzckINSQ4MLngcyXlm6CapdKrOrIDVJJjnMB6r+TSM+9o
kHZFWLvfxnWKwuBugGr/tl48Bxv9UGU0zWPj3UmyWZe3itaGK+tBIOPt0X+rAUfBn2ljz5IB3mAy
+5uCuA9ZWSfWd5ubL57OQheRWBagSHESA1as/I8k0WXWm08z8TbgOKbUfM8K2s1lVLSeFeUeDDh7
hkpaeAh11k3OhsqLDJCUWPTTomGjYT84o2uygmRymcIj9ais1e6Ycwj9qaa73Gk09jr1LqMVEVF3
A7kXyUIJoeknMtVrhOsmEW8b6K4fbChoGiYLYXr0tfDiKWRmo0AnfxqzJ2966M39nm5bcbmDxuDn
aa2pH6+kelBNZdJJMY2QgJKgw6m4pEkSh/knWlHkrCLvJuCqif2Z3nrOxeTLy8xPQBCQRWhi/eur
nx5wHqH+ukBsSWKYatjMpywvct8Vcr9AFVBCpWMJAre+P3MY/5EDTJUfydt+sRWoFgExkwWXECF0
68FQAhbWcWtaDWLiS+7kr160FwiD4whrb9x53XmRqoOTtDKPAP+4x+rl3qADeMM68TGfJfhsZHUX
dL3dyAPQDmG0Kic3J7ruL46j7sYFX4wZX87yRF5kLDYcwO/x8pPqLRA09qwe2joVaC0ZDVV3J+++
Jx89FslonA4Gkmsdza2j4e2SlexUt1+6tKQZn0mXGtvmjy6T9HVhKURuwwWp+rM0CwPfnwIxcG4H
nQ91kfNLSgPOBEsrKKHY6I/wor1z/AC1FNrYfiEq8pZ6/k/JM5dg5Swdysde4ewJYZfXO4KaJlEM
0N4KXchB084eZWLD6nlLqQ3vu2BTbjd9G0Fs2zOzruWHh1G8fhVY7fKfB8HBZ8Tf9VVLht/82Ski
KsQX6SpLnOEiuJuhp5aHMoXHL0sFBqg85qOuujOBHuGltl4qEvaX8YnLqJObxW/DrH6wujIPo5W0
eM3cqL6v8C7XoBQIQKFIWZO8ucCupZOi69f4cVDKgNPtclm8N/APJ9GCPWohnZiV/rlRjaT8qKYa
mKwjo2jyX0UWRRWGuHrYlaJyviP+1nYT/OPa5+hGi+JmV6cfCijbu5WKK+PMh/o/TccxHB+Rc13x
TKKtEeomxAzR5nrpVR0TM5dU0ICRCveZcr+tNdNd8xVgr1hVlmWYKlaMVqt9aSBIZ6ED1JGCLmCQ
vu0KJQsN/e/Y4NvHOObjwAnmCqJuXnloxhGfkjf+mAiORsDirvqCrCRE00iGmiB+FRbwPSA8c9OJ
fau7jF2l3gOAk3KI4IL23oy0E70T7OlwYSOBZLvdrf8SyvSHrU2YjM/k/JNp2yFYx+EMw0ZP9kPA
EPcVJRtfbVxxVNqg/ecPfOwpwEW4/Vi95FC7MVWE9WNgc0bhr4nXF7JFFq1HBZQrqb95qKXQolCy
INqJ2uanTXewlN4F/Gzq0xFbf3muSsH4O3FC+wGwbzQLDfvuGtWi4ZCDWKxpWBQsftKZy2EHzPfK
bR6VGBfX7R4ZEpDPwlHdnJsXDRcaIHzPxwwHioRvJqdKUhhlAbnX6zX/XVUlVlFwWP4+TVWq0ZnB
GwqU5dTepZu5d1VOq6DUe+aEn6AV4PFjc4DXJnp7/DIYSdu3B4I6dAwGLHf7g1RsCwYsLtrClH7e
CwV+yaX/sg+s0vhCWwUy+yW3MItl1eKPEO0ZWkRgNaBstLAGzxf8n+BXwDJHQ0IVrTxfdCiAANre
ctzOqtsOJpHP0IKmNVCZiazrYsfNSxLyQqxw00BXSyrBRIGl0u5eo6djOk9KOHjeTW7HucsM0BM6
PKGcXwzURdRrTrQDCN/CD5HR/pAHBARBkIehNiJhzs4ro1Vex8bQhZpkSu3xRwbJfbqv4IzX2aIK
+dKUxc8CPvHWYEvENirXRBFe+ywUQE5F1hohYVpY7MNa6vscDgmLggBAAXK4NbUyD/yUaFlixcib
7uDDv54JS7CjtTrpL/HFg5EaJ9a2k584fS1UiCNe0Is1L4i/Mpcb1RYqRW2EyiHPkObH7Dlg8GSn
CTvHwgx1dtHrr90uS3iIaR0icS4nqhTC2J4Z4iWr4YhuOLFDaU9Mbyd7DNJ0i+aDNxomS6DHpviE
Df3dfy+RW3Mw4vuQR6kNeDGL6xs2XCY/uaMSsnyenPkvuL4+mp4HQ58ZoKDqOEitm2qGNizUM4io
y/GIVYslAC4HO3J+rVApGkSaIqLeUQQz6PcIxC0iy4N5esnfD8xOfyxmKqfE5fdbpdqcsI1EvPw+
MxU3HzUAvq3NTT1IzK5WtNpEObmGmY0gOdWCnpCrNEUqV9X3Rid3h5DTV0JbZUXqYzolP32WokV8
aoxrAqAE93c7VDJFcefonkISMfvNq4ZwrkfgT+ZBsx6zDo5v6HKg2pCjPXGNXLkGIwZ1UTdGthVB
ldnIs52T6XXKyZ5Uy4qQ8GGzlgSa3m3nDOXvhGEnv6yn53DPpzNd+jI5i/a+NZ+Xqg5ZS90wVz4Y
ZaZUNqsSo27ZecXLQuJ+kIrgZ5WKI0Hz8M5w1o87OQ/xpJNDL+dFhIM0dkmTL8p/PFwBeH+qTJYr
NfaTCEwpbKRUXUMooE/ZWYzMTxJBZJ6g/A/8MJw4KT6iqtCyL250v5LIOmvpzkSQ+GcUizTAZoli
mlLu4wExYqgOFnGz0vIdQmwwO5X64gD5urZvpOc8Oq7COl9UjapgmqS7BfKwi+SfGxIAgv3IwYF9
KTHRYMzOwRFdLtzGI6L4ENwkRkviv5ZY3N2uF7T9sMJZu5xn6hoNfm1FojhCtbv55BGspQCp90oo
yQSGHPp8v8hRBxGQ7A+FP5UR2g8Y22i4NFCEBhmzMDw/nmxc2ig6+Q8+SxT3Xp8685P3bS7AYr5u
S/uaQfV9AL+DswMbOi5MfwTgDl7zGs81oFdZgMEynrDTd8FNzgf4AhF5SId3Kiu5RZfZElTOnW0Z
qJ1gcHl8ysjKxMcNURcD+/QuNTKEBGqTQvudSYcW0gqbfF7SS13frlFi066WsaW/IuNlPgRoyfUi
D1b2cPK5EvDtXTlrL7DZ2/Ksj59/Ev+7So5E2wHVjw4OxjuUFamUqmgBdwseg1GRXMy4d6Td0Re1
3igDRwvGWJBEd7eztpvIvKcV9cr3hQSjmwSB20SprZOgySWYjngqDOLnov2v3QwSf1vs3hKkBarK
JRT0egyOYyZ2/jhVc7aKO1KFEYZocNr1RUkMw71Ypg3b1sR2iatq6RBOV2p+LaqlfR02NPoR3m2J
CrdBApyEXWKs98+Gn8yjJir++2xodvbk5h4K2egf00p3z3JN6rqfw219GJt7G5OGV65zRf6Ya9Bo
0iVZ8VSC0aCIJx9SDDJTQD1Un7cqvecBoL2183W8W8vlMHFSpkhXYHxS/1jygznP9L+sKc4ndisL
UHbpblvYXKj5au3OMC+kM7uADVDndJInnJviOr2roGNrxvv1XOb+WdagDIDvAwqVAS4aldtmOHV2
QjMDM2kFWyMzwoPeibOdZw8ufpof0tTMXV0hsvMS+nZXkzTxZSR9mVp8Ze5SW+FMBZAV5kvGd8es
bu1O5Y/iTjS4wp2JuuzZessDVkXvLdleegTHKQuv4OTt24pbQ6KSBqpAqXZhBFhH8k8WkdyRCA+y
lVsE6AGx3hV47PxWfAuOmI3/2an0S/x/2vqa90eMX/yxdcBhQlm7vPedb5xXC6J3ubgY7778O9Fy
v/pDMHsRclM6nJYIw6SxuUN54fe/fRPfzu6zZKpvAjxkNYf5Rc//rTfA3c/MHkdgE/KzIszZIVTy
0eIkSWcmMW07aOeI1OTqvCQtpXqy2OvR3xleDd84HEPFODLuN0v41PJ4UvX5JsVtdXrHu8zrwIIZ
FAlamtl6Shqez6S1A5AP5C7+MuKcHwlwZ5AzFV3WKnQJaiTwSVOwvBzLqDlv+mhDFFUG+cN/F3Ru
rxGISX8ebUXdiLztDLqnfhXae+9+JG2VPhsjzzdrQWhEAr274DFfBHJo6gSv3lCr6CsrpvUVC9Wc
tgtYZh+cIMYd2jir/qiDsZFe7Huei6Y124xOdc1PVAvAyeouzXZFUf2LI8p/ZkEZ+8k/cFFJo9ZV
f1TdUQ1ebuw8m6Y6+A+GS6MZSdIhg4aSaf7E0ark8vok0Etbf83m5q6VdY+D/GhGex0m0SsI6UBP
tRY0BPOy0o+VrqyALBh+JIcH+2r8Qn+H35cnRZPMtXdWXIuFUsuNvg/g9Eele9nRj+k28RNkYwJ+
5OEWHFryu4FlgP+rsQHbhy6VMPOy6mcGQdi97Oggc5JgNChO7uo6Smnal6pz2Fehtpc1jA5QMyVu
hm4beGTSMb4ghJt4FIE2cLqzx/MTNZ65BXtidpbbC91uiKyDggnpJsuvEltwR9/jRwja9yRt5ri7
X9VypEfa1podhGfrpwMRwOSfQFTZ5KltE9z7RQBpnYF47VGTBjX24hhAL6ywZd1EzBhii+1apjIH
Kk/8MjXDSVghFUnHTJCWZwDGz2z17CV5Gqm2FvWwhm2SjqD6/qlhGTEddfCtMgWZ8FLBbMS2kwlj
6UCccG4wWcTn4JPYS4IPVCYksGqPP2ITtVHm/HGtDkZ4zVSN73my9Z/sF4B0ybRgXnnU75zH8ZYG
x2RrCke9cpS1Ywb+J4rORG6pFXiYZvsaeFBf/MazffQbtZ5YTKRgqlrADkv3uEKjw25PKchL5UWU
aogSlLI5fQirS/h/wDQuMeZqVSw3VXsmV8hgfgzJow5FkCrVGxhdONOWP8SOydajyoD8QF0B5hf4
MN9dAfE0bMoCGGLM3TDaLWarth56LgK06/OdRvKLUFMDF3sjLzdrlOS7gJ3Tagi1DAfPEpxtn0Ye
BKwfv6ZsRP3DY9MkTm2g4XD4L6SD41ztYHYfAYpGb8vIgc9qX0x4lEltygj2Xpa+yyg9yxAiPWWR
Twt+lUeuTRhk54nH1GG6yiW8JOwvN+9ai1mBpETlAyXtDAtZSxxT+5Qn7kS5AXaJXIlZKqhHE7je
kFR+EL5gNEcp/MsgKNTcuXG71pzZXLXTTX33/Jj5CGVLcaSsQDGqv1a+++EgFF5aMWSjrfHXzSlU
Q1VALyPMbV6PIZ3FL5OXQHd9ROUR7dztX1NUr6+8v69q0RzHutIF6kvXtqLjHnTSMbJRbZmD7Dg2
lOE2YgjS+McphLNYh+ldvfQF6piTk3lgozRpgbkXzeXpagVYcPTQD0VHnW0CiX7slcLz71BTl7QT
4olFPR3PNASMajFlC65G87G+HNl8msGiBazoA4isCHU0bP8/YwFREBVSA4Dqx9yWzz5NZpAXQqCZ
RnHrrbhn1EK/JI8XV77Y+oNnep5yQlIe8OO6SliWuVpIjG/Bs9HyypHJOnIrHAMfhcw5sPrf+rPH
OhyEZxS6bn7Rn6olUar0NJwvP6lWry0HhY4CsR/gXDgqjTawYnk5db9rLQ+hZMfEJ8XKfmt7HzJr
xFuZiAaQEkcyjlDp+mGuw5GVMq+SIsTivNhO+I45cEE+RKWPDBqZ6oIJNRDuDDKKCGljyeAWnNaR
K4I6Zm0EfUeZwa9+PcrZWKVI2UjC8hgaUErLll5zGxlU/XsDrTmsdW9GEFKhJ8OYC/cWuXrDnTPb
OHlO4CbYpxlSdJ0T3P/j8MMjxGT7HCEJ7A1+cVRj9BJUJJlUy9isdXZRkshPDVKKbROcrgUB35IV
S0JBdlsxdJUHibv5yIFRhFg175xqv/tv5OCmqyG4XurFNYt35+sI9SMa2qN4SNNO8jbKtWZdXcmC
sZ4FqMvDPSHBaE/HC1TOaNuNH9fTWMrhxLvTcqy/L2gpPTs99Z6KAQvIIhWPixT+WqxifE6x0UQS
epfdLW32j63OqBYd9ZxR/ySjrgvwe+L3fxVvPxsGfo9raAR4hAvs0eSNcNym5CKP8LhNt0+GmZX/
fFBXgJ6tyyOf/2JnDxNhNXZQSjI8vcXfncKl+3z0GiupGBKkX6DPTw4JyYb0Rzgp4qfKqVTbFhOT
r4rzoO3x/0bP+HNokV5qvZJvIFoQQwdYnGJv32EAI6CciVQ9oRRbgbydc1KLgar9CjGUxunmJuu7
6hW6awtiTbDqEFH9+cfpHv66DgG7IqwxRh6ESmauNvnwNR+0hG9HNASWXdrjPEPB/oXAKN+idCLY
atzNQngX6RjUX2TfDdJQCkHPa1kNaB6Da4Vslkr8oACb7rOLjsWV+cDF6TXQuNXh35kElEhjVjgz
Fmco8rGcQQfpMGAtDLJodv1uT758jqlGzXQGIlypLjTMkDp6AndzaP3XFv+Cknlcp8ArTmUl/LAS
oaSJlYv7RxbbWyE6as4LDEQZBYrtarw11GWXq3ihbxtvv/ayokSAKKtHSOkyUXeXkUBJl+UsioXo
9/7Du+s+lfu7if3gXDrlFxUHbJ/qeJ8d7cvZgTBrqOL73YktD47hN7fDrPIFhP16uBHtP4nCHKx8
O/n9JuMDHZfB9dPYDXXpYqQpJxLhrfYbq9yQH2N5x9LQxFUwWV4s93wX8L77bcYs7fXpiEE6IZvR
DuweobgnnGBSiKJCkjBdsoOUfYOnufzXeipTYTSSOLCZ+kwHrDiPawbVNTI4iLP4gNWLAAzGUmhh
TdgXxW5tUWFr0Lac4DlDMNUxGfIgqD8jr2O4XRy/ifqx7w4hRlI3w9fxPhlUnuE41PRo8zS37SWG
KTQw2seUNKcXni24gLj0eX2o1KuHtuTxANDkuDKQUgUZSM7IZn9vu01/5gNCR1/xeIGDq2/6gNoG
63fpuTJ24xNltHE1sPtGolILSJh+9faZ4Irez0AvOzOt3YzlU3RQ88GeNxUB63EaJf5Azs/nf8un
KoHvePyMCtJf1zEkD880JR51QWhKY3I0MnAC/+7Xyvshs5Iu+ffYxLBGjo0kGwUeEO4YwAYdKY4t
JSNJbSYRxqa5RgXVGMzBum9vlj37pCkdS+E/wwG95/AEHVH7e8PmVJyNeI1+N3WC9EUP/Wlg3717
fuz1u8QZa3h5wQzT0332U76NTXAprkZmsKZ6M75sthF985wX1feRQK9nB+7gfdmW+hVBNR1hrSjH
LvPE/1JJJuUuMtk0GSYOFxNkopzkd08P/zTTXWfFhWYaJ6jpzOsubATBbTAC9nQ6UGPRIETHkQiB
jJLDG5xxCzNlX3gKp7RsSGjXiKJ/h8Mr4p1Sl5hRPL2l84hq+fySQfVPOZ4wkO9mkz9VnPfP3MfB
DL/yQJi7uthGyMUTh6GvqgddzR6RAsOoFE5C/txalctbh8K/G0Ccbk/dfqGM4S18o3mPRuNVNfbW
RZ/+2J++CGH9cfpn4B73TM2C7DG6YQ6r448opLia4SkMlpZZ8HTK43SLFb/Lg8c4RPV4MK+fEDsZ
KjCupxdh2sVhfbOgXbtgf+h7jM6DyIlNQ0b6zCGjgtsc7iUX9rtsOhEDYB2LN8EI32g+7v/K+2cy
vTbEydTlz2CIhsJrPHfKeaG3Fzh/4hz/DUqjtOplDob8Nsk3hmhJSU8d5uZP6zQFMxP42jopQnqw
Nvz8x6UvU3BjlUFZEscBvNOlpshyM6Il7czzvNsUP7V3jSFGhOblLS3annEQVJnfxt+BwODFkH+J
E10b5H2w4t2Bl6T1LXYc3Fpou1AYRYM3hfVdwUudiRUpAzzqS+xL0msVb7sFhtJn6agKxfD3SnJn
3dSPsOHfFDs9M+hzqxZcArZvbZhSxxupEMXGw8lw/tixiDhIn0GJYk5fBOey20TGi/3s1oi4gPOo
wtS2teFBDtX8ggCrh4kkin+9A/ENqE2H2CuLOexjZCe8hoC9kCLARVLLxVli5QVLT+BbbfRc3tPq
fO/URH2HzH/l0DiNWEkWbzebT4wsdklwPJpXHNeaUkly8uf9hasg5xgD7n8gXns9W2aLOF7lqtoA
Hhl7tgZCl7CCnABFoJafoWbsEKT9qThl0Q8Xg2+x+pcwlSUpqFZrsWBXxGQZUNA9TFz5Dl9atQgH
Kt79x6vRc2w30ccZsxccK+JGB9J/YerGZ64fBekWSAv2RYbIcxhc5RjKngpM64oVErAmD9q+POd3
UqVT0z7d3HqUQH3KiKjasVD+tKqjGnkl5htHONgMnACkSuiG66mm1Bhg0rcapCwmJFwXLRmqszvw
ZvecIN+mwvt5yn1KMUxFXX1/fhwieK5o/ALyzr56R8yQaD97Ycrh5s9YIp5xSLljCnbl1pKJJlyJ
Zgakm44DK2QCpnQXSv2u3Tr920650kKLm+f3NJPAJPQa3DIKuy+KKB+FOJpGKKj8K+zEdnt94NXP
nqrsFp1VuIPJhgjhxxQAtK3hvMMbwlNDNuzf1oLdHc80CDKXsIwgyMZVHHpM/dGpIQU3U6ECoxnJ
12YjwryN/i4L7a8CeueElWkL3q2ZnUvp90OHl6253PBdvF+nqIPBx+Ze2QOVYqgFGwl+GCQYzcDh
rBHprmaPPe6c0Z6Ht7AwwcrlpvnKDWoSEuDYecUTzH5Li2/CgJ+9UWEmeHW1gaEzZ7XkrceqytRm
62ljsD8a8JZU4lQ360NkEJnEnL507F8GxdtmgTB0V8IB8kS6q3v3KfyAJ4XLP3xYVzBQDNVnEB6F
9A7GPuLso0UfuPGT5kE/KjTZgWmz5JkZZXtwkIl2fHchv9HVsVRJJpE1iwFOuEweDktb/rHIHJXB
fMdX+26CT0XVBkHk136dIlOZD53R5PGHkbmuU39UUxLfExGiOUN5prLmus/ibT0uzOC8TUgjCaKc
c7PG/RkKMH7QFaeJAND5/kM56/DqZx1mRTVLUMpHpafILhOTaYZIPCxknN9SDy8aAenwurYe5AQl
D8m0fg0qYdzBAAOLrle1Tg3UlWh97SJWBlNSei/aPC6ZgbaeN1+tg6eFuZcrh3fbQVmapKZOlFtG
4CnRS/4NKEESZUuh9JHA1RnG9OLCA7UICLoJAok874LfAJaVnbtpJtPmpk6HNT4RWRNHT06pgQwx
2IasOshYfSASXFjDgGqtFK6A4cGhixFmlV1PL3g/9wiDw/QRPT8aha8n1k22E5Iv1OXUAcqFG+dq
vqJbXV1cOOrpVRNzBo4+Fj0vHzsyJAsbMBIePxxFYLSu80x2h4ojDPCYx0LGI40gRuncPNKN8eOX
3UQAZbfSmENfU5Oo3sS5ZLIIM879JHLvLAWRzuKda8dFBIQdNdC8xSBdrmyG6QMxfpOu4sZ7vV9J
6Cslu6ZaVmlULikZ9wrxTKqxQLBfkps427SpAIlB+78d7kYYd/zpF+YckJharsnS1aCz1POFFKN1
Xzk6A1gZqUSzasujxKruaUsYTjim5Wmq/vww8CkueRCSOz+NIElsV8xyo9MidcEooG5rcKMe/H4p
aukjHLQWsmubZ9w9jUsSxZExFR1gVmU1zderJ0Jl7D3h6PjllFY5KDC7l6HBQlECUyc+y8vr5FX2
Znxmn816/ObezzkS+4ShO9QvCPl9B9X7fEM3RlvcbJ+bXVfvIHzrk0mF5NBAmCpQ8SVOdbnCq93l
nbSmJSalFNtnewliiV+YGrSdfxll55ltZQjC32O7owJmwcOKk/elfb+NUqsEuKxZoDw+3YrHlQPg
6TLjcdCg09rkCHLr+ogRmacgxQ4BCKS/ONYyTdXR9rfDanuOtAGL+ftiUEkcKt37yNAPQrQrIL+R
ageEXfwQCL1tgC9Ef0tqB1gzB3WgMES1xGyOr8TjlYZhcujh4sTcorCq+zyGfalfq7mjKJTu3qJJ
7McqgQGHWEhXunOsFQ7J5mW3WLe5SvqTq9IKvyyF1tFqC11J4FbikIMTSeNF26Ex3U0nWtowVc6Z
mQ5CiANzy9OYndCYnzP+t4bItubSAxfZCQadZLPb32UIyDqr3mhJr48eii3NIT0cGQgyqyuidNeZ
zDCIjnzOpwNcRzefIfF52BLICYJzMZOq8BgNxulbQ/tyFxnSPINoc4W2WGKviXZ7NuhIVs9VqEDl
vBQyytanQHdAkkFLxYLeZD1LenPUMBTvGSGeVoEoW6rCPeB0Ufkx04Jsk4GJBdMW+V8JOMS1lupK
uPvOIOxgo6NMHndJcLvUCauF76UFhLjEK74PcYjUjl7KETxRUspXTreG1jEz4g/iMEG5/CqeU37O
K1dwGBoMBZX8eC6ao/Z7Ti2wmKe9CtIphROKqWF7PI5ABKNQXt9WHQwnhIITUVjYjQNANzqp69rN
wfTGlfN1owTSW8KTsL2JC7vQ7CZpz4Vy/ZSDTDoSvAguVlLz4qj+zjY3mNfnbwC/dZqx6MGrVgO0
AIohbuNMj3V7qdoFNPM5bsZulT6/JlZXaMTc/ms40r5N4W5c3+30jYEk3fs5k1jGdswtF5pEzhjF
0+IfmIGXt+4hyEWybx3S+8QUYOJ2LQdr28KTtNf3H7YiCHHct49lmDnmcWUSs/XWXU0DGZgCTRxx
gIDR1pUQcnYX7df0WNoagMbgtE69z1/zZjtLMNeYAcDJpXcfuiQKNBI5hS4OqWd28RcWA2aSfS51
e5FBp9C2D3nfYVqH8M6KFZd+eG53FhxEARBXflzbU9HwCh2sCrQ+LkUhN2EsxHb4Fp9jOl07Rc9s
FZVw/1BvZ+ecQMsOll6GWxp7WL3I4kV6Ytrk1crkpaPpV6Nzqu66xsX19LhmbH+4LLa9mVPQ+NBu
g5zRaVBYRRANfkV/qcPEruWp08PtudrHoXGqvJmmrdtdWCTBFFwWbaZ2YWkK1iArAUomp7kZoLwh
Hzh5gdoPGE+aTBRQq9aoBKbl8XYAOuiG+Hw5aPoBejFsELRxL5rtHDMNvyTsQCC+X3m+nfo5Hd29
fJSq+AwX4oVAxFsoge5YJQJ4YoiJ/6gWQK77kiNnZC4ADPREVAUneLWPqiz9bTKaqPFanoCjkbCH
BOyIoHuPi+Yy8Ncbl8jE/msVaEGpxl+Nut7sQstbrVfdvDTZ0lmM4fUxTxixBJAsSH4bo7Wmmp3S
77leRfIw2jwl5SY9hM6YqK6viMoAEKFFjU4AHiyBzY8W88j9ZankghoxhRbwcpUF5+iYT0Rdyk58
AbCoGR5fpxsfqbRCt5H3IVCXNSHW0vIR+ilP/siDTWK4EdibFoK2MmIbn6a+8JzbKwylTr8Xkr7k
dAYpSVA5NHzt6qFV8X1AwazQrGgzfUPSsXrW8V9gnOLqEdIwj7rgBZ1CUZWPnwoXlwOwossVoqcz
PwdaaPy/JJ2+ctGwrCjnKRPZBupZpa/hk7C8y6gBK9qDMO+13YeXONawXGdd/M3aEbLZdwq+3dpt
jHtf6yA9HAL1eR3kOGOeA8tgac4/joLzQaVuylnpBF4LgQPeV/LXfNkPhDX33JOxW+7F5CUXIgRq
PCDAYYFQfHDb2VmowEo3IPZVHAkiIS86g2QwTmxcWpj9U1vWmNSHRM2RTe2p59rS03RoNQk+JHHa
7MxyNjWf6d+y/2UpeQ2C8loI8Xa8ytLSyftdv+OVMNoMT/s1K2g9el+IwexCY8H+b/ki01yECfnK
eiIwxLk4ZUj6iM5nxDnbculnNrtyEAHTJNwRhMIEHEAXv8ZjKRabICMKXFB8PK8s9VWi5cGeiPMx
IWeLy2ArtCOkSJhF7V1OuqLsw48W5OdkVJ+OF7sWkrcCZWySSMfP2CmOU59+fwjEDl4OWn+wUZl2
PNMAvWi9zBDTauKdjgTGaJ6Llr/51yyLAR1G8AJzdQ0bOmZITz4S2E8+4oKsvaqqmE/VdQwNXHRW
rCkYep4lnre8r4fVwmX32NjpD+FQ3kFD7UfjVWjHjBF+XAeQfQvSNN7YRIruJg0dMHLOy4P3u2BL
wtxw7zVRFkXSq3enNFNwUwDtFrtSOuNNdiNJCgfIO8wnhMfS46GHBIkc4jjxUkYUNVQGRfMzZjF6
QQbDTRm5WrcJDhK+C8fH4Yt8Jdn2wPJfDPNS1P0kPtEoKRC2IZJfTme0gNkPY0wsRBF3x8Ue44jo
PjD3R+AyXOyV/4K+CnWleofOKVZ2gtqgnfKHILto8wBQIfbhCdS3yzhfD/8DdseCgkpYZZpIbEqi
fFgph/iDneolKYoCx/2cQYvOuhkpQtLBZiqyi6j89NPhqB7PGW4s+nDBwysyUeCLic+Slv4bSYA1
tTdgPGFrfIj7UIxDDafx9R9K9o6dpHrbiNYraytJmJzQkL+ki5OqFAHwCO6vm7HhXjVaRRtG7tED
qvGxZj9uw4zaRzb1fL/p3sB5g4G2BHH9DPa7qwGAJg8p8vOnkMCQral1wim8tRa+gSU58miSAAJt
JZ1YjMu8ShO72sV1Usc++Umk2DkJGFNIzqv0cfw2UlLBfuaWjjaKOsIvT0ltG3IusInXI6LSAx+/
tKSjnTIheZ+Kx+YgJFI5/H097Txj+zG+GaAHnZOsS7rnlMw6z5u196Xd44nLZRT2LUaruw6G0M8c
/qQ50HQ3j2H+udS5r6z8byaVtONYWy7ldVGqEkz0es/1lk5iAfcd9JqfLJU5QQhwV5K5C9AEtwTZ
vpFVFvgVBlnZcoNQZXVDe5nJGEfymHK4F3Sf3UPhTUEZaSd46ZgLLOV1W0ZQpEaiojtjd+vamJV1
Cu0G4u+RbwVne6gJImNUS0+2r8aAyD7PjcRd3I3xw9TOuRcpkoKol0ECfmCAj+ixXn2f1rpjuJA3
zmODaXQa5aVyMPEdZA7jJ6IzsbqJCHJBeXKCKFKLm2GrpXXa5Dtw6bSobNJ0mYqEXTxx2j0Bk+U3
gIn5Md9seKk7MtOnXSK5gk2znWXdsg55gjYeTVCePRV15vxV6qRV5SLPMVNtnQIbXOMEk2pYRCGl
p5+yM2JDxaZnbPTVOD9G4RwMqvnACi7Ig9/aoZueHe1EK/Enqr0+o0ElxutOOYjZJfGFBG4M92ai
45xyxHTstSzF/vd6pzF3E5JVw7t+BAALfebjQFCnYV99f+3PVu8lvdB6RuFe6G1AMZ3MrZF5XXu4
WQO1b+c2VzyfLrewyJE71HZ500pduWM0LKe2r03uANh35YMbpEV88Zb/rMmHHMqfqV/p2rvaEwAg
80nyPOWTqxrUZmiAGb+yR4P0KJFbfpX/gZTHswxkHgallj8AdOP3sTkNo0kTdBeIczaWUFCRlyUT
/eBB28mB9Zj6kkOu7aFfPTeDjRYJlDN5GLtmueCZ9QbAlhkvyN2Dr8WXBsx2OOi/6SvkmZ8/COBL
a06d5gp+n5Yj3BLqSRIdwpWwK/nv7/aXIsp1+WO1OkuiF5an/jMhldFb19JuK6wEUzfNQj3uMKpP
WBDWJhnpxpc5gIS5+bRGlPQ1EpdtGKxGCimGk/ELe87FHLN6vQpYK2bYd5buZjO003G5qWLd21bB
G6NmcQRJva0VncJwarDJJHSnHKNZEdkTglu6y4A+y0KGdP3GYx0/8I9GtXAB1b2vffq7TCE/mjq1
VHx7SC7I7wzOwANTZNpg8amb5zLFgcUqajO04ElRC7cN5/gTBKfzOeSsqfAi+iXNK529L9MyWrmY
2kr0YUOKEpH4ciaiRwZcXIzdhfU3c3TPNr3nunlFCc3XX8LBYv5vFqz8Rpv6TC+1onR1NQThHMtH
cOWsvbIsIIKBUguQ/oDr4UQLxxZXkXpJBk/6qHInhD6v2gRCYN4+yDKTAbNG51PCRcIZB04xfJWI
2etYRk7UFuNsFN07m/BqSPPQUsC3WHpXDkVVxHlpPtNeN6OGxHIUNWKcOyHIEpRWPjqP7N3ta76u
/3S1bG720nu8bpgkPKgsg6QK1hIKbuTfVKvqkJ1MDUL5dLbDFWDGWDRFCR1RQlbQWb0+4r1JSNHJ
SNUDxpML5ZBR4tIe8tYufYKziLKhxvLBC+C3YJC2WGJ/Vws1+91HpOLca8cLjvKuawcQRGaXV/ol
oEVuESK4G/HQ9i6bcm4CYQ54IZyjI6P9Kko8gY3ygsgUan5uOBmGxV1ISNmzPFCC+naK9vn0/H7O
VVBouE/93xqnueGCrSy7xOY+2UfK3bbTQVVLTbd0jDbRmIRnS5fZKxU6LzXDJ1l8Jlk8TExY/koJ
34tui6//PqNRA9SwmRD+HKGGTE3TrMc5DaBl3NabGVlbvGitynTt60qdzJAw/iukgWSpTi1YrbRM
huIPjdeNpLxg7bK5SWzBeZhkn4bgrEoTOB2VrjSHKNT7rD81tw+2l0M1J+Y/RWm6zxUa2yr4IUIf
RkS5IP8Cu4fFW9UuxH+5rddCa/6wFAiiIOSBs4/bFmj4AwDhVgZWv2zkGOqPY0W1UtVfhbF5rOzt
Vjc/wIYCtOb/6w/Z5l62+njS5bMpNH/cykOz1GthSHsAH3i7VNXiR3BCi3AL8QwOEVXNj8KXkST6
ED0lP+QjiCHcHp3R760henpn1w7e6f4TMhkI+BbOiwvDO2oyhyq5EtA2ux4eaabvN3acrNIzSIQz
zjjNUSwlDy2eZLy+RD2bC+XQHJwY5cJyMV+P/fVAJR3omT+sGe76UO0hNzf1xcKnF8mENKzeZs08
AHQVfaZztdpg+Q8o5YoIny0oVSDiiwC//89RQKpesGLVLQMo2ruW8kgMtAC9dpL3zZGSwxB2CBvP
a8UJQMDRnvMcMf76Nyvfu5y1Ly0QxUWKwt01YFPzI3R8lGRvCRbEut3rDrshyRI9WmeIIzhUtB+r
O2HGrKk0iKBmgTmrSSC3XEUq0WQ1uaWpIo2CQVrVzyhVSVLnzYW4FkAJUxVBgc+bh03V6wnw9JVY
oN2ZV1k4IJaDTWWnTfp80y8AeerxqqTKuq9tC82gS/1aM7QcW/7zPaqSHwJec1XDh0crXOcwzX4X
olxVR6LCon9ZLoNls0oamL6WBtQ1oS3F3qNulXWR6QwPsKvUd025k+B4ZMjroYELPCdWTLgj+Q8c
jaIoo/jBxUnw04X3gtEPNIG7oIpanvQ5R4BGgt4Q2dejXQpLXrXt/PU2ReBUgE9Qs2Z/g7H+I6dm
gOxsox4RA3PqkCzaSerkj0vQCzoFu1iV3jwlm1JMWQP2MGrYI3gB19s8xZr/p3gtXi5WT14TfeJL
215zX2yWdlCJXCgcR9Q9nuPuOYJyGo+ZqeRFyMqHyhhZBzyKhcJpGSACf4HXK16X2IA1Vmh2Ltx5
ytRm/2hxX6n6H9JedPeE9+Siau6IMdEL/xVWA7sTelUN0vWPI3wFuE4ycC4VKMR+GTnXR7WphV+b
bBHQ8DTzooMv17ONd8H+l92C8P8GdChBqjBzJy9c5YK3jmtajs45oYGYLLbX4w5c+40Z8UCQ23Ni
gSwq/XNersRPsouyggNiqAUOygPULviwHYe8m2Wa7qAvOXqco6ECkPbq9uylbn5ZtJHoTem8W4PR
iwxYQCUvQn0Z3SZysT2Az0zN/lMXriNu+saxr8+lprrQ2I8i95Z3AKbaSI1T8+1Djf+ZRN6CrEUg
jn9zKjiXtRq6966YUZu+zvzIzXFBHi08+yWspo+9/zjT4nUaNrDm6Bxf1YMrqCLT3ZcFun16AYn+
+PlrFpeGVHMfFnvungkxP0j8jQz2f19W+u2XnkGuZF0B29sILyhAtrbWiZqt+shvLJKjVvDc8DG+
bLO2nk5H4B7BhZIBt0BX7qA4omnYgz0f00poSkjRpVuU+LVniPYa1tm9SHlmBVnAP96OCpk2f8NO
D5DnVbuHw6FKej/PUuQoZbjWzoUMjZ9VIsVKJjzEucYrlUGaHakvkN+T6iUcJL3f7m1PRB7ClFIV
gXaUC0dIYg00MQjEO54wqK2VzOeS0okW76MmxqHonSqJad7VMAR4O1uo/7T9/FqqX38HlQH6UJIs
aMbBf4r7oJ0yjxJ3Q9qu+GGH8L28ZfpwVvV33PrNZxpmWB/Lvkr3jm7XNrGMvwSJgnnIklq+9iqi
6peWAb4EuYld28FSWtBq06b22hspeOLOBpSv5QX8CxGVIr2QxsmNCtFEVA2qZCBm1WaqedRVK9sO
oLx9WK74z5Mnc4XMcQHaAa7RrBidxdM2KYIigujfKc3SlldqQP5RCpQFYk9OheIM0tFzYiMeDKYE
+UKEb1kvl/D0zhfhOQbvRdsyi+NhR3lRALEIGZBgBjece2SjXvs7hgDPJ5cZ8iESdZzaTbSfgpHl
/5JMi9xen3JQK/2G59oE4a6R8lkBd/48iBKKz6sk99cqcr1anW5cNH9cHfoHXS7OKHyK5/IZFREp
wTBhuT8sucsmwph+X0bIroPsmUbjs2aenQr6QIFzmb2m2KRCxzmmfG0wRs7t6wESeO8R4PL5hY45
X/TE77D8mKk0FQ4FrrqXAlyeX/vfwG/Wz5ttRa6pJi84qO2kkBoVANpUejNU5RdeagsRqDZ74LSd
Xos/RJGec0uZx8FiYXYTsR16CBEBlybtwMkoGpkfkbt5wSMzm1szm1P/YCCKfY6oXxSgOVOc6EvI
t5ULm/WiWHjGHKBo8+qu4fkj3wSi9IrPyDL37+rOuz4APAQu6lp+d1xAeltH8qZNXSmz8BavE16E
lV1sDXMB9vkIkr18wxnF5Uu7gSZzFqthBRMhIIKdaNI+6RxeasWDxuQetFQqMZISWIDeegA7oTEK
aIbBy9oyyp0sT8dh4c+WNk3HLUtm1XKpfEc4LukfED2PMoyxqnKpsTR9QHitojxDYCriT6x4csuj
0i9LyV5H/AjphPXzW/osvR4dyQ6Va+lRQLMuzRL/e6WGBJyCYuCdaz3iL+XUDvbG6P61tUUYXKmm
KV6XktN7sUk45lSj//1XTVjSOwKTRoQuFfDQUav7PcYoigZg7Csv1DzDv03KV3LF/8KU7gGlXLbp
uHfUsCN86EHyhL2XS2GBCe5fLHDO1NDvksEO02Zjegz8n1yB9DMLJKbRUJjGETd64kq/cnYt+1jQ
tShWPDIUPVFQaXET037G9F+fKJQ/VEsKTXD9Vls9cvitAHWanBHcgCKTfapxLKBk25zM5ufvEaV8
8kLdKRJUleXNYmwwsGjPjnT/ipd/iuI0kOG1Dsk4FW0+l0wPqfrrVGLKzZTmE4Au7CyG/IkxHM+b
myljWcfsw5AQx4mNEWGkX6ywrdTSxr9FspUpoNup16Nt5XS0aMC4bZwMgbd2/oNTQWgB+y2RKOWR
bSodV3X9ydBNirFqJQCKUOjoIrxtzvVaVOUByzVGcsxrGORC8IItf/fXxi8xW06KKECWgL3KNSQN
b48d947rdVu8zLOIaqez0mVro36due58P4IhbMESpURR4VfXOAeKIdmukDvp9REX6Zhrkbm2KU5z
C+0G4mS9uKQ10L3lar0Gm3xPOOiwlHLBu2em5SPJ+wlXsQWbmLP5M47mM91WYXJInxlRYMKVQXxJ
fPyOfd6GdwF93jf3egn/SXYcWYk3Ht0wThbHciLgp2Ia/4R5ttc8+jh3PsN6R1CLbuEJennRKPqJ
/EpyokN+T5KVpnaEYqz4IpuEYxYqWtxyBiXWpD6lsO5Xxsme8qjbhfqZeTxSQhZiEbptsNTdONCt
IrZN0FACjVUCK2606S5pmNop5MzxHIHP/SUw4JSrAqyl83qzr1yyaR7ZmgmtldNfR/EPxsehnrzj
LBPi6tTCh0Z3v+aYOKgxBeJEyuI2mowd4PSsmzURqxD0vvG1f3wfie/z3KMdAyguxZjRXFdFjimS
ckqzTD9losQz/5BX535vIDyh7OlZhbZgL42TARWiLT7d6hsilGJmoNXTYmFwfetC9QK5URmc+U2c
+sahQU3BLlP+EXqLig6XxkRbiUpSm4Zh2JUzhWs/KOzijEdOATUYr7Y8bdbBU9jUPOGCGI9vZsaC
AuDTvUWmTnwbicosj1v211DmUVs6f/Iq85PhEGsvGvyd6bp9GKjLfJYeQXHuy7IQ5h1VwpaTAqGU
YotJusaAcGKm/ysD4f+hgUiMtqikv+eiBmw/eXq4imJaMiGK24zVHtu3GJNTo1EdDZ3/IOHAUG/s
jsQDMZUWBQXAcOcmA7zkkdpcN05W+CuUEaLKEdU0JDK+TUt6uUEkDign8w2rXYH0zdCrWvDweSdS
jpxOk0firFi6U4jHClKfA3wj+IOwo15U8A6jU8aXLKK5Im5LztLwCgRH/XTKkEKntwIoGJ/ycl8v
2c32aOai9Niv+2kt2qVmvdMvviMC8dkc16f/yijbeFw18NdxLNMppYh0xXfVqYKmT4lU8cBRoN9P
nGEsjAVhPvy7zpRdtXqq+pII8NCqIPMV6Fvpo/ruculzdrsRXyxQOfWA5CZFuS8wvu5quIxls3Au
CTSS4udE/b8wildGDIaeQNUfC4Xf3t9oZdxSHiMjbUpkK/Q+pqixvdgBnWuBym5+GE7bUD5jHjMM
W6TNjLgMbZhNhbYpBQzbw+EgE+7drrmh5TTEzKDREbMMMyMk6wjmIjcfdu1O/ROGk/mL72AeEGsm
zZyJmHxZ4lcK2t20TF6jpT43hxADv8uTXmXKOFV2k7Zy3Prn64kbZLl2IRdJBDcSCPXThlgdvi2P
HkMCdPZkr2bqGOHXaVdptOzO6u8H3YsfTd3Www7vnWAGi4guCNTEltvI41HRj5oGc5P34JVnPjPd
5ZjiLklwL2VyHZQ10xdUxjdK25KImNPymJjhPXRrKQITs4A2i96icruOvEGXcEskOFUdcRtSj9XE
f3qQ2//T0k9Yz++LoL0kwfhAvrE8mCKw8f7mWIpqNHtdVvGLl/qDysQQaexKrzUNBG9n21GjqPNy
LARINhzbGRuK66uxPYhLCKvdgXpeVhI/0EjqJGExhuv1EnDYOnm/FFFGcoUtYfpy48ZA+cxkaRJP
zV5XhWY9Q6/lTx3nug+FsnpS2aWHDdUuOAvfc/UwVH9/fM2QX+x8diIofzEBDKetLYA8gyOWccP3
EEd+FE/l6DNmQanmyEYtgwxB7/OjxWG8WxMLbmzCQ/6mpgbTdJTrfkNMF9nBieZ9AGyVRh0mo9F2
a+f0OnQIzFdcp6BuMZja+dSm6RAweqmSlS0yv8HtV1swQyAeH1NXGrtvhw8O+t7162E7fFGyu2oy
fh38hteYD87YHXXG+CHaHL9+Io5EH8z6/bS9ZhVP8NnPtz+gu8CRfyd6VUC8I2g8HKbdt22owKe7
s3nz7QQPLZfliQmmHwz8CF3P/wU5VX5r2d4mDxlUwDC9IOe3r45mfkQ4nj7R7CYBXl43nx2IRklS
VbEghiTueA234GLSuI2BnSRHrmvLq8a0UZjyoNc7qGHiA1u/gHQr0czKYIhUAp9ywAvvXc2ubnnC
ZlpABO92TlptRgE7gXQE9cmAi0xc9gd52+/0vaubUE/v+gO/U6tXwdDbHKLYol34dXd5YE/Dlvl8
aKWlKT6ksv5nystcdU9W6wlwWM0PfIefYaOPAuxTHZKECx2vA4jBIrNBeUZI3TfUMeIwuZ6+bstp
60PNKTwh9e5XTnl0OnYsTzSJ9zOxH5/SS+6exXFAXnbSdVdfYYGevnOkLedpLhNFIbpUdnokBfdM
Mg/cgysXyKzXS5nF199Q0f7PfEUyoJa4GSCJkcSUlNWQhayZt5xZUgM3eX6tYS/qhxhTz06vv2fJ
ViNzgiogB2A1ikvpVp3TcHz7ysxgLyzhXRpJQNtiDlZyCwAzx8nfwUZVRvzxtGtOpYqGIOpzvfS1
BQc2a1UYhbr9LugL49Xfi7rvo1gJs8DFbLE+zq9rt0MeKu82NAiieZwJ+2npkaEpkGyguU0Il6CC
iTPnby71X69Vk+5vPxHgAgvAJcYaT3z5BGRZ11ZUXPRoTrjk4DBEHg5CGGBK01rT6U1rlogF/qSr
QGfIeerqodKiKwC9Gg3r5XGkywaJvfX0sKhVPXmpr3hOahCZxR9QlB41XrPJSlTTWxFQZj0RSKwB
e8/0iHqSznqs4SKCNQNM5w/li4544wABnpwyEqkXZwQVND1oP6pG2G2S43pcGIUlW2oHKS3iQhc7
aNpu11S8mVVCl7lZQzVpLiTj2P5+R1o2t/N7HskgEuMKCXh8+G6vUzkQtVtramHcSHVQLX2a3vc1
anroL9pEDcY82SlgLTQjXXy7WlmeekbnUO6jfBY94WES3RtHqD2QWtiOOGvSIoaBRuaTdiLR1+M3
SpnoImz+pk2r+HslJIbWm4Nc4Yv/tHEDU/K56FqfDzcuTwIBKwTDg0oVKTQXMvL37aLzZ3+PCFBm
AO9RdSofLgbOKBQ76ZcSalkv9D63zOtCun9p/DcgsBV73V67kEU6J2JgWrkx+e12LUyoQumfdMD3
6Kwp26PjKDTXzhBAOuegjw4sO6Z0wWvWzslP+LSxVZJYnCtV8YxX8YEIhuj0k1Trf50x4FuCurJy
UIOEwYjVkw0y4vNcCTNvRt+rLtWG3ChFXFaNd37k9vlnq2Lo+0c6/0EHWXbn8WPSfk1li8wUknuG
7GOsO5yXX46fVMhsr1GlvXjK+8AsxmzrotlkD6nDotzvfDqsq/BNmsoEQgbdgF8z0i1fG2Vxn7IB
YRF9wXc+X0gu+YwEkqTQBW+DFg741HCgd81ECNg0a6Ixf++SfDMwkHRT+LL49GTmmhp0Cm3by7Kl
mRhJi/D3cW8JR7G6vzxC4VZCDoYOKuvT2QvDJMbL9cTg7tvqFRPTt1Q3sNO5KeyqCu1QEAArilwu
bcsmrCTeartQGKl49OnjCLtPPwCukgTaQXVSghDSfPZSaDL3UQaVsT2HOwfBOgjrnoZdiqXMLpJp
dUvzmNYUQVZO1fzsaLrwdK26k9GwhB+vx+A1rzM1BESro1uWgb98E6vHFu5QKLE5T7B0uFP4o8kY
B3p1kVlsbmo3+a/d9qn2bkHkhwfll/ANsE0GUTvKPaHZKPQK6zefIulmizZ5pA+JyZQa18gUO+Oc
8DGG/MTFKrnQlPqS80ZmpCtxaRG3Nj/duAc3ExA5NzHIyC9dKHquzDvfmj6vwPmE33AJtAxpKFD/
P2Hs1nqzfoKj8Q+2sPVab+BFPM0OeSBgO4BOHX3l7WKTD5dToqXa7NGcaWM/GfMj2O/HQBDx/xbf
thuFcpwEb5x8NDy0ZHO13BeDsx6nmB/qqwaoiDPdLwsOYRcrb0XemIPWFnovy3SDxMr6Ri6uHyAs
igX7zVrWPVBNLRnEnUlPgg0IN6InN+P+6LcYiSiW8OkU5uoGQlbaaXcJgGW4mhANnpc0BBqJOpwt
wMI37CiPXI80IkvLvbHy71X33AYikW/ZKippkesoGZ7OY9zk6fAGdj8bvBfxUUne4Vw7/rs3PC8R
hdFU+tv/XaHggCsEPPMzxIN/DHFNFR1tKT2b147z5fdTsrJHgjdRZBdhSrpJHj4p6CSnsP/+iJlH
m3zDxAM/tPW2zT7zt+hwJYwqoy8pwxqHxI4EQBqEi2V8FS1PzxR5CKhn0JWBwEhToztVVyVJjC62
H1sVYmEutJjA5PqSdIzCZu1wDgwDppCZ6k7pixnAhjsq0YNbuGi1g74hGLW5dlU3Rm4O6tgv9X1a
uXF9UveBqlUL49MH44GKjJF8E/Vds+5AwKnUurUhipdxXJ1O3njTC3x9KF0yZKjMxTHc4jwCyuK+
BZqt1k5q5whX9nvXUDW/TsXfl0RzG3cl46L97u3GVoJahzErwxef3fSKYmBKJ+83xzqDp4Skb0yL
ClmHiWf47cTnxMTaew+qYRkXjZEwXdO4FDgsc7IcAwJKmN0NrzirT5emCzDvYZEwcwKzSslNn5xP
/59Cf8wwJQk6eLoh1RCU0xVjg+5UJIc3r+Y+HQ7EXFa3Q4lctgtq7CEWLNy6b0hT7/S6ph3hhdcc
VZDR6pX5PFlRXxwsMgoZJX4S+2i8r/7HhJOLloePaR6dvQN3FjJa1liYcQ9lG7YA9MVl6oQBSXNq
3N7lj9b7UEOrRjMQ40ksoBuniyK2bafSBtnn+nJMZiKcxjG8LWjuVNQcYVNTt8FAA2WDHcovuY6c
3pXD75F/ZP5Md8v92koAiZKvKV6JvOCGCyEZ9PA9c0lhQwyznhH++WrorCrJI9SD28TYBBOKxFwv
IxdE+sHhQ60zWTVZO56/bKpNPn9ukAR96qxbZfqjGR3ZuCQRcKP/8rkX/iE/wetI1OXvQ6Pmww6a
DbUp23KIsSRnPsalFftgamfBUsKTzi91o7/BRn0qjVKktmXqLmNQSguXPcm2tgq0iJZsLxPSK6VJ
5P1lndk0OubEiJqdCnzSWMyI1AbNR8O3a+86ZbQKVClQSjNKAP+WEvJ6anucI3bUAe1XBVgUTlST
GUjSQC7W6q+w2TEBpfgBzdfsIHl64AtesmSdhNTXuNoncNWoBM/4BjkV+bZjDOsPkiYdMzgkqT3X
JZeQQKVqZIZCdq5eRl+DLNRqaX6ID2VyZLtcB+GYPMp6g8uAFZ1BTatVhu5mJjs4ZfsNgJpBqKp4
YYQy1g1kKy+lye9re+x0wEtJ4ECLyXf6a5BraIo9+gs7n723GSZNizR64Y+VZwcHHNzl/txEPEeb
eP2OlgKgmVD4sHcsG3CVzDZfeHoUtWBqsb/mZAhlbBNfhe55kCXCmOiHeVQBkApGd0UGjix1qMTO
M2cHplS6Zj5CmkZNUkq6D18IV5Ii3t4133GK4VC2K0n0z8J73REO8Ul+vROlFQL2tPBsdZvCbjcT
SeXyjaxYqEWCure3CB6DR4URnkk22YVVA00gy9iQ5Z2kmCIQH4PgKljuDmadAlGPxoYZDYJbuzA2
DcE27mhCize6XboIJ6AflAli5ZeiuOkvi2ODFXJrS3phSa3VfnVGt3KJOIYqJZw80EzMPCVqyDKW
BLq1+FH+UI3R4KEbLPoVplJ9QXZn7FfoV1lfKtjZvFWdgCV/9H7sm/BKTUUclf7ODNw5x4T3Qmox
KS695aQjZ9vj64pAZqHBUzTti8RprO9u8DlQCgsNUjZ3JUOR1fb0UqroUHCw9WgtJYq4lnpo7xLG
8M7jvQpPjmR8AExbFSPni+/6BvQaYif8dgvbNE0Ayd4uCU4DMyxMffSayox7Jys4/s0UAAaNRhRS
K4n7aoHErmeSdSQJnoCB8yg/mynRzF7WihcxBKt5tIVlxSms62znUqZ4E2DKi96zO2BQVBdqOBCq
ZxxNsXQjn20oxhlXr/afElglj8HsVPkkZ4uIPVRGxt3AVJrwg7PkkhPXkhOiArRGKchYtJ7+ObYx
cSeqUItqaKk9touSDF1EM3/w0EPSWMwj1LosomAA8MzUG+l4jATLqpGTqcSUySp4vl9KGgI1CuZD
B4DZOj3lFKSw9fwT2a1Zz0q8udZBg5xe2A67/RJa7FLGcckNKsvCKF5NM0bzWE7E4nKeVgLJk8yo
lzzsC5l/JL4p/6S5BgCjpXGqvIgrzl2qXnSsKJYavFTYcWjNPQy6pfbjPopZmvYTlnWDmQTdCCiR
/6SiFQM70NrmMvfZ1E9pUWVGAiflw0u5CFGEjiQ2+ubMdOH5fYMZMy8OAtdcJK7lVFnbhBh0xEGy
1Ycb6i0JXKqdP+aLIJha35bplMA5x/Ue+BveG11/MByrMbdYHvle8u1C70KxjBX/kNwJDLCeIMY3
pyw5V+S8+SgScF5E5pk0eAS09xn37LK5F53YsVpr2qEbBQNvlotgJPtflEBzBIPk/6K9cWD5+d7A
gT90pwBXxNObCa6/A9U5lD7sUP1fXHHmfYjULl3ltt47YNqruvoY9YS4ltlUkD+7e63FHBbkGB23
ut5wqh9Yk6hC/sv5PIMh18AJFFY3GYh1QQvAKzzP23zmKzekmwFeR81q7Ne+nvUhGN5Zwj0n2Xoj
BQgWY3YqjaUPXBJfuW+cPC7NwKpmMmS0ywawSj2Ky1vlfwL+Y2aC6RExDPN0KDOO3P4eJf+31720
nUhxaPuiyNSFfpAr3rV+zF8R7Z1COJEi62j+uFC7bVxNWj8nux5aNigdhFtOJMJ/ioTe4HkSGRWk
5cKaF3pxTo7q8R7SGqkxeO/Gij2FGoA3Vp4Vy0TE+gL3Sq6JRHk069MI3qeNZlF4ZEUYEpaYVU1P
nthL2m+ELdyk+FKLR7ETR8WH6PMfWVI4bNpVrXISSy6kyPXxCXpnFBpLTXsVkZdO7layxWwJHSqp
6dzwq45x+E1NtkmfR8tGMR6f+0ICXZW+AF+k5IT/MG5XCJs5Jn5TW0QbSQOci8F3qILI0o3i0VLd
jxBjyba9gN1dTp3gqd9N95LqMFfhFejWQVL4NWM8jxbPYh29dPIpiO6xUH+FizBcyqy7p4tYIdFZ
Jodi1zAbRjIUEjCIz/+WAVlQYE0hy4SlEPU0NM2dHdlatnZApuKU5Yzx64l5GB3DC8ITbIuZnrTm
TzBE95YynqPSTEKdUlOX7d0N01Qmv6p29JLtWVGYezzV0dgcW1py6/yjpCfMHF3obNBGG12gcotd
dNqY2DHjpeL5Us/QCTuX3O9WpS0egnAZHU6OHKBa3Pkj38AG3eTYNR3vJom8VdjNlWsS8hzp+tA4
4xCH/6Vzwj7ejSyFk2AyUbS00lGxI3tZdGt52yZByksWyyqkCQxkRVTLxg2hFNneHJPuPu0kSwvR
GO4yikkUKyoweg23P3NaTm23PYzujN70Ao2ZSvjwJ+m0BXaatSLwgHcsgqBGy+Na82miPJX7/p1n
22q7OLBsgVXdu+ne1PMC0MKyKpFH+5It81u/b47MVgghLJ1lAZdRZB4NyEzMnA09z/x1Mb1It9Hx
FVhuON/KU5B6WsWI50MXc8aFHupxavVKjDRfZoviAPQqcgXSJy+OvEhoJiq7IMcpZVjZ5yLzT5ZF
y79pFoiFAMCbWpWoiqQE4kifQdApl6vxdV4bx+zBOpE2bAb3777ejXSwv35B8Zrm+y/Yp5Kb+VIA
/lMZMmtBsOLgyRWH6wp+YmTPKXWjByWKImFwoXFRcouh6vZ4YEGTeFgG92gqfu0w+poKf7ZeczSn
KQ2N2j0lXkL9VuR54xgDjlKEMiSDyuGUcpNWI18M9x3/B+z/6WUxmhmQ5gM3xiatmdbEm7b2w8BN
lKHqcpM+HZ7Ogu0zqfYtcRa+MW+0vjnt+TyM3OpnK/ELvklhopIgmQ9S2aU6QKwOXylyXNIFrAzS
mu8xl4MEu091kMU5+SNisDO5HND5cBbGmWvXuBpydXVYPJoIeOY0hE0J2qIfuLGyWtfhOwereeCp
cnpbpT/PgrKXEyMOITysrp9erqg4pmOwxyo59k1iTXay/b9SofwB8fBSK3ZOEvGvfNx2bq1YFgTm
KqcNnsBTr1ZEPbaSpRag1xGQlWfUfZAJkr8EprsJyqqNqCTNBRF3TK34omWVsEuwXgkScBv+KKqM
bjOWXeTZMGtjLhCERmHl67a+tYLIpgGhApSvF6Xf9dWc7o/dnCh0GoMKm+/YsC75tTvoq9u0W7pJ
ajG2I7GcLJEkZuOivSh5Qj60hl1OqE2KXORzzE3MANlOMKZEmKUVmvdCb1zgJlaf7V7aRfWe5gfx
DbZ13Cn4jbIpG1INqTqE7LHLff8lZkRaO5Fo9Rx4/15ZUcr5JAcqIfD2GYJbwOaewxsXZ51uxc1g
/4ixInpgsJ3KP7ybri3xAXCK3F4Wyk13ce2J4oykxMwsk7gY7oX0q5/UV7g8AjMo++AH412ef1WY
H6lSnZ4D33hbmC0PachHE0bmr5S0uP/k3P92trsmCumrY1q32L4GqawBcj/tkKXk7bEEHLXxLClT
iM4gYHK61122bcUFVP6tlbbJy8MA8LrKCsqRXpo5Szw/8vMK3gilpnrhaODuyMfS1rAQPodffDdl
wKOswFM5nJYfgyUO2lZQzCgO17y/Pt9s9jjpv1rtnARdZccALOj8/cjL5FOp4DBzYhAVAqtP+KJ1
QjhmZWGx1MXeT+xj9un3Rvd14Fewa4NjhFVvsCDtXE/4Jv9qdTwoboUtgysl3xGuJ9K5zTrqD/4X
B/+tAInHUBZHYuKVtr7AL2Tt5+bEverzImfFQL8SJ4VEHixf4TcHUVndMVpUN9jubjAH9lhh1OMe
5kQiFPjOds2EgTYl80XKr86TerbWzfXp/VzELaCKE9fUXBZH1IgicqQ2Wg5DaTTw8VWJPlaILoC7
0Dn8ekQ/+t2j1wyn9VrcWDyX+xKZ8lbCc0c/QOF++RvUygLZCglIdJIsIiN+IUZK7s2bbmpXz2U4
ye/QkNqj9Br0tbbtQRr9n89g7QtXAhVERNE4QiarX2H8NZuy7r1Z5J0vyh6so8sHaeot04vLaLiK
PdLler/GOeGimwKs/DM2Ujl7GtZLydKB19UKywKRm5GmzMB6/v+l88aFffxGAyDX1HsdsdC8cGj+
OMUMyTPhF76QA0UD9NDYmjfu7uvsTFCvnxdEk5BkZFGOaNNLW5EPHHUvG86xR79+TZrK3FymMsIm
0jUv6GUUk2eJTRdxAKms+453I3W1ddqIXcr3CC8uaoRTRiiwien8MWfWVvsDXqWJV83QiAHw1Ddm
MtyDJIUk9/1dnY0/HTg/vCGvEEFtWIx1lLToqbLB5vL8W1MjEPk70/YGN3Z2eUxkkRZnAInBQa+j
T9u6x4/bEtT3Rl2Qvxip3HP0pJ2RIchThDEK2EzLc6fMtnhbgJ5T/VVYiTCw4ZqHp1HvVGyolAdC
mTozVue6cLJy1NVHTwbV3r86NmHGek3SCz9UdO162MG2UPcei+VAJ4FiXaoWzSk29Iuvz4qztVvx
rLftidJvIX4QUZKPrHDPn4s2iouoeur/tSrJJ5kceuw7W35cfLoPSZ2aRfC4hpYVlRUdV/6vzez+
3FuqgB9C0T3aUzpAQ5ImsPQRf/lQLoRbogeQx+y9XRGlqJpbV74Hr6nzJIB84E0EOU2QBYKKms5C
I/cxCPpJbnQdsmpgcc5qAN9xHStODSrc+SWFRI2fWfJOkirgFBcPfcuSMDO89HEt2iiRHmtG2uvc
itBwaGA8AP+jWXNIJjY9RWk4pF8e+0kQXmfTgtl/vVGJl4wbTW2tGQ2CuMPuSt9BsTni7ko4xy7v
baeJEulTYF3qZ7GXOTcThXoEe1aYap0uY+ZV70XX+W0e96LVuc2PZTGqBU5bj6iA8nwzP0SC6EDy
5+hkpe+18wOoQdCKGuPDNKjpMsE+p0wTAIOguXlMRh7F1kUOkKaqkC30GmrLWYWViDFZ6x+4UzUi
OoWBdCu2YpgoeWU5FSObE8sqeUJcW1V+q1LyvgOVyYZTklze/TK+kAnCCNLKfoQRhtNPPMdd/2ur
AbLjU/JVbLNPvzy2rAMqNT4RlMZPWkWaLN8+SqH0KmDzKDIxgsBVn9+S81SXJPOB7e+K4yM5LFim
dqtnz8x1ZVpz2vq3wyveKTcCOK/z0zhYvW5Lce74n6jXxHnAXETJnt8zC2Ew8qo7wqz1hg98t6L+
X8GQMMCoXAp5T09t16M7UW2NWqMPOE43jeuxxJeSMG4ZOPL1hyq/66ZRvDvzj33kJpRX0Y905pef
HHRBu+GkFxglgINM4gg9R/ncqEVSpZBaL3FfNjSzxbYyzUAh0ks1cB3dkM7QH7hCkmDDHyhIwQvl
Dvf/GUkP4uF54EdAQJ243n7paLrCO1DCTQbiGLoTa5WDlCIpW2hqEaTobPHmV3VZJHiSa9n+LJPY
Mz1Qy9xwb37YsX3DkXamSIojuyIdOnH4WMUgy2At7Qbjm2buLv+NR17rM2eIMfaB9ZDN7M/RjuKe
k/QCSO4OFHKn2yIn0wzC5yt+cer/wKJHFuP9NftIREifBgYdZhqH9VB84gtUFe76jwXXXZpM0Cjr
jt6g686Xt33uFrbt77w1R7aSXoaNIgswL493RQglm0UrqPgm5QvM/4sNGqzLjUo61FiPIvwEchyT
Ogmh2JvAc8Z9YbxVOPRaqaE5klhPRgP6O/n6XIISd+cq0w/YRjekn68oITJZ/5U0jldh90BjiBhg
6OqwOg2uENZ8m4zhipPQx9RXo7cxA9JigKBFbCpNj7NtGwWUITkiFHSPNr/PbhJkj/vaMPU43E2i
pySMIor3Uv1lF0bNoE3tI9bp7i6SCUS/+aXnRztRHNsFMZ/4cXcI22G41QO0bM9SQ/XmFLGjDDTW
3l4Fboj5/SyJcdDKuyXy+iN6WeYQUqh+8xofkC5DAo8MjPWe8PoGnQPjB47gI3KcFSRHAcyu6KcP
AXAarWz5gbmwy8D9yaLQoE3lk4FKsDMfpbcpZXoYDHzPN2srloYpqC0VJaIp5JAKW22ZcSai6a9m
camqzeIkr0smkYGsBBtPn8B8n4zZ8hxf++RXWXHOIj50UuBor3yvbkJFwIgqpjgwFs/v3n4PnNQ+
ny5NIqH6vGrcS4vD7JG5FJ6IGR9/qiMOmQl6zrZg2negbUWvB8z1Opve+j2kvoV/64oyF3XgghH+
donyyJkQAVS87owF2grRJLNmlqlx6HRNxMUjwWi7RlHo71pj3uYh6YUbXm06Xdz9z9wE9y9or+t/
xHNHwT2DaKeULsESmnv7nyKbEGV4HcW/KSX1MFtpo8iuC/aTT5+2AW+qRjPRO2Zm4I/CHuSrFxhg
UWeQ40tcuZq40P5+y7MVMGSHSR9IXrSIYa0Z56iBQwh2iMulPOO3XfnWqfuL4qv3MLQPZ0FZNk43
5jR31QVQf6OD3QYKQslMXFQJ8iuyDr9ZL244Dr5e482fP9IXaHaXdDt7AnF/oQmWtt+XCwkpPGWb
pBOrWz906/5UFu/FZLH9ot+iJveLYqJqGgL1Aw4YA3zz4PUDqF/0EPEsLfw8pE3SbzsYVYHHXt/k
XBazQZXGU0X1ZRHwh/2+dEqrGmRj3spG1nMymzPNZC9jxjS8pGKyuCdi7A/tCqOcezUA491HpM4h
EAh60ykfyq9B0eapq3fJFlyC3yBPNvFRhf+HHVa1fK7licxgycFCF4b56EmWODiFwfLoBmdV2VtX
Hiqr16JTPTEh7ezyi1VeDj86IBGXK34CRq+qgUwqNpwAkUh7SfXlLdT0GCO3NvHA1pBjBru9yMkC
Ri5NVHqNgnHJs03aCSBLVYMOD5M3OVoKhWbR1C68dOgKlQevLPM+Gyb6PwJeBuo330OStVw22iW2
UwE/V2qWowwi3j8dNIw832fFfNJbu2sXBmsWImPEO3ORUl8qUxPB0KDgyyEEo9AY81a8RM5cL3/j
IOJdHOM8/7MaiGxzR7HwRJ9fiAVt3g1V7NAm8wk5CQdqAia1Bu36o1Aor1wx54B09MbJr0xu7MRn
lzlzMvTQJOwm1dV/7/ZgwpLkWGmlin1lcPiIHu7igleTv7zuRrzpYmNTMdU3f7/nvu5/1q5xBmAO
HBCNY8RcENKCXlRUZQoTF5J6s1iaCURyTWeWSED9oipjYF+BFvxELZ8NYXTBPw3dDJb8f2q0McZK
1SZxH8ELQFSJCbjgAYPPxwDgqtW0HaQ6GXCmXNKmTVuBtiugVmSMzMSX+foFFPouWU/Y5cSJYXiT
1nflbv71BzfUdjB8fXiPG93EqhSUh52zOSngE2IHAV39fWppn5P0yG6HOsgW0D6jhD6HHcIFsL2K
bSm/0hcQ78cmfhuQYhiOkouHvGJhKggwa8pGEskvNp8pl8o7clWhaiVSE6EMDo8zQ2LUcSxo+elg
GgLeSXk0mA8W8v1vevyN8MhZTl2uZ9Lsk9xMEa8h6R/qQgoy4iXxJZeJtK6b5kg3A54SlUOc07C8
R0JAEpaAPlTPSUiz/XUGp29YL5Enabqk8B7IRHOjpPVT0Mlk+0PJmCdwMlZj5rm30D2u/u+a77na
iDL3PU8xzGDCY/1BFxeQUDHHDs9G5MXj6gcBLEtyhN1+FavvWkEEzCTnk1ApuNsxaLz7jDXXw2zI
E6cYb9nk+vU7HZjQL09WMUdzn1K23d0OXUPt0SZW39p6f9eeq1W+vjufAkN9UGir138l3TAZt+/E
ehQEJ1ps4WWulvRjWqzwJIaJECVKMG6UY7VeG2952zEN1UOgmxD9DkdDmaTLVEp8mlcweBx74ZIz
NPBeTayWdBvyPCxgqpm4FDzdZI5WvtE3uMZ5+o7uvxoIzlgeHH40AvQ8ebVmHVrJXW2fV+m7YDW8
NoR3JIlOBlElALzlwn/w8CqG2koS5CwPmkeoPEJmhQ6WC4ZNcMN1J2TFZNuyvAreb2Rqlq4goLWb
BrbT0TvkeiPzGz4ZSe1TtVuMAKLG6GK0MHOiIbTv8+ABmTZKtPZsotpTfe+cQNKWSoc42War/sL+
V9fXEcP/ChWAxNiuF4yhZHQCE3V41ZAsgY6XsTKP4o8bEhhipuKRzgQMz4xLgG08dU3ippyR8xaL
OAFsqVd23AdSc+bIYqxhnNAco0OYE+hLK4C00fGLkRn0mOcbvsCqwK+wnh7dPNkf/hB9Z9ArAn2Y
ElzpoZzAGMDjvdKUkdMtUoIVXBE0ThE6ptvO1UOlHbgQcqrr5ZKtl+XbYoF8LSptTSXC9uI9mpu5
1E/KVjDLmY5/zpb8nxZxpmm41R6DvtihXwtTEERJNodgq7pp6S1hCFLpF0v9+MQ9QxHPhpIG4HrZ
1X4pJqiWaCEMnVS7+svnlRlsF0RZw7qyHqF0sRY/o/n1qeTjiJHlCsnIwwMT2pp9sZI9VCjfzxrf
N7VvCpLaj7W0W9gnrym6dJ0pT/tMvgTz2A4JfUJwMr+p7HWHUdPXlweBotQVBbPgQz3RyPGqljXl
lzBY9Cfj68RZC4VtmulZealLWA7ycJkxl6HEFX7dThKhrO67REnU8oOidPm+fteTOxuv/x0mjxVl
yuylQUBdAic+wz25xx6IiKG3TtY/NkRrfMMyvYJiI3k5dYvnKqOwdmKfeoTA5bxB9gJzaT6Lfmr/
B09L2jIU+mxhNAbUntL224/Hui2olw77LDda0/lW1yPIwAnaxYOdDf9dnD0oO0cZ1W28vwL8dhxP
534jPSJJol5hvTrzTMpsOXiI+z+Gi6vtrLMVkKnoxi6nBGUoisV+OoX40oFz0yMGZn0vLeZDZ4FZ
itV5QiuFT6DA0jcYVERazi1lFcKpuCsFW+ZzMRjXMqMMsCLG1hqJvTNULjUz0TURRja1vgwnB5td
R3AswLtcMeLSL4At74uwCOGmtN/DSLjPY4RzyN2xdQEbP1oseLUH3GWht3v1Uj3IEG2jAVHNXQSu
AO9eaPir3iLfFEZy07/5NRYGzW5xjhSVmiw9wcKGpW2MPp0zIfW4q+MHNQfMEsYzTyja/VOm6e8o
xnACScCyx0vM6r1s+Vi30j60xxp3/lryeM3oGPY0euz74QWG7a6Mx4ND8DNXqdta9/XI1wUBVefX
RC+QlDxj9WRSc/4ldIAksUiFD0F1OoA3aSlGdqL3GdIrZfZxv3FJnyNOJTWGe5vFiu90vwb1HD1l
C23dJM5L5nNFb8/7HG1aarX1nrBMCHL0fMS3DiiuIWPEPMjJbSbYYErQ26RfjBadYecgLuy70K/0
7kaX+hONP5/XZ5dW6UXrouUFU8yyKYQgPF7P3Gt1JLSF+mzjJpGbsVSxlvgUMghvZe/1PncRCtji
gBCtZu7cU2nZGcWHuDil3W0aBYAS/oCS/0L3ZlnjRijHNHh0WwhHSOjqo5fLTrGVPolj+7aZuFZ/
d8Zpll1b5aforXKIHq2Cm5+9OD6E1WrLWREdLqsViUvurB9sv/+Xe6vqJlAiia2Pjf8nydQyvFa1
UA6Z50bz8XlYwH3re2RuS+K0BP6gsfbadbagEM0VA+TOK6n9LGaHZC86yOObMO07/RXKrW4fwEge
iiTE5LGi35TkUveh/Wd00aKWvCJz5w52mcm3JXv3yLPk5j2P2EGGzkq6nRbd79hc3fVNK/VXPK13
hqlxa+Wq8Od80VKk1xuH52Wi4q27R5uh3DFZ/ZXMEVmC7lClIUsgRXguETtLxqBo2BGJM36mBpbL
BtbKpHbvM8NGGLjiaepuzEe/OU/WenL9DsYok+eqOVvQSVvQIvfqYBcIpsVW0Pqrn0DsT/xiHJx/
cKztI7T6TNLRu/ZjfD35iGyzS763KmaMeqUrPRuVyuM+3voqxxB4Vv8KgZSKIr8Qt8GwyKhxqJwb
KujCQbZDLpMwGIQB5RVhlPmAnOWfJ82AAn7lvB9aSMzkxwJqR2I+ejYqAg0j/+RxwIMYfOjpnr2g
Mj4/KzgW55Vk7uGGHnf+oW81i3gaonq8kGQIFgHc6FFyJqUOyG/5fZz6i2zu1EpCLxqykWs/7TEP
8kZo2VsF6NaMHSpR5ov9AE+qNUCKz120yU/clsBLQiYcnkORPoVtJRcciS/jj/i07CRjbzj+JXgD
F4Yc2zoN1f75miYTm6BE2pg3s+aJAcSRSEIChdXBEcx6vUo5kGkHuNe0mYALvFcTa/bHnXJFDnKM
Yqr6MKxFvPWdo9RqBfBzSrZeoLPUo0HbcF5XZ3u97ZnQz+pq4L7faMZkSIu/Elw80KfXUU2f16FY
YdWW5xTzMuLhpLavrZVTIxIwyVtuId5TtSdxy6b0neg2FKgRXuLQjO7L0vFrKidreSABB6vzra98
DapUEpVYC9XdHZd83CV6sEUmc9ItxbnAHyAeUlDRLkt93KaKAZQlIswD1uEfgGmB4fyt1j1MzAvF
WSZbn7K9h5QsuwGrRYg52SJIq2e6B+2hJUH9Xx9RJy9+v4zuZzw2m0vCWT0hrfiJidHhUB1H660w
ySF8nL+yrOvnE54I3G/9jwi+zhqsSiYtPAgCYzscC8a03yXtCs7xPtavkwslacxCOhu3/EoJEwAn
IHK+QAvCrQbaBx5FOg724yoJs10A995x9mFceJYQaXD7hpReyoRM/j6YooXUoOAKiMcB7M97m/1g
PZMNepnXSNj/XVRRfQ9Eghf/3Rim5MFMhdXzjcJnFDzaQ/4QCneTq09Lxxutiz7QnieistqMmFSM
rt8Pi4yXo81q/oIjnE8TkmPEZM2NTnqCgtnG0btBB7rpeuM9mv7ETLE24CoaAovgrfMy6+18Q5D5
euiLytf8pa19/NMwgO1VGA/uZpq6+H5knlbmaOITVDqUdtPfK366WDpzWSGWNmiLSrYq64gEvTpc
0ZulVZtIrYFOgAM9VkoTkHlHtC5X6gIrxqKvf1iYcgWgChIscHw7v2Z0QIM/Tzl7/RH9D8OkhSbU
w1iU3gMGP2lt0LlHAY+5iStQm41tOLpicYWXRvx1Vc+uaXcqqtJn6+td7/m9/Bj/feu4JpqgJY56
A+rcAV0rsW3QCL9K3mTZGD/q7uUgNpWH0wR7zp0ase15kdGqXPMd1ZVPlMiUwNu0raFDSKvRm/ey
c0eT2t7T2SUNMkcF3zbYRMW4okE3/ZD3WPgnH8FYq5hBraEGcahJqkafRXWzJrYANekMxDwpN374
/pLILQV8bELPROWlZtnbi58UqNh89KQ3WLWFEC3NvGkjF2FJize4Qm3CnvPRq4yf0kGHf751PnYR
gkSugAHYlI95pm/gSErtuANESV9Dl38TXKTLBO7Qv/HMLF/hRMLIpaFjpCyB2rlVxye8JX2tDQhc
uD8ZVQA0PI58dX+HnS7qOdz0PZGONXCRON7b0DT0qExBKBlWxQJqs4qjdbX177GtJwUCqeLCR95s
h2ErKBlCPEE3HjXH+OUvH5D3XVF3OMYFUnnmW3UNJ0KOieMGHPFy0aVomfSBXARZz4PmnWyDbZDh
e3TadPGb1BrK1p7UpYmLg7gdwJ+w3depOPeM7/KsCpnmXhG7SmXUNWstAEMwf+juYs3LcajjPwyW
obBdr2aCLUl17F6ySsaUij145MV+Rlifggv3qqisIbOpMW31j0OdqiZv6915spRSG5ujr6Cwv97j
PT+c9jnOn/WngteEhBPbnYXg1iPBmW/W03GKrexFBEfAIpfpnsnIfSOSCKmP9VJmGv6woJpbJLmU
I2Vx6JENIR8PQRSLVp8Bo2Pp1D1TLhZgdVfr5/J0Ct5kZiC6kvQKWnjc0xoiwel5FgcAbtXkUDCR
s0kgXONpLcUm54VGntv1TMxuKNEcLf+iMCKA5kiNmLBySpaML/d+C0yi3zigH8psUsuwvL3JulPF
8zsvJDZxSeYUoJsT3HcxypUksPKXyqCHVChCL3R+b+JxgAQCF4LLCHGaKQkmlOo/vpRGIdOhTW64
0xQ7cRTeypmZgYTQLm+ZKsXgcgugucGNF9mm8To2mGvRKcmaJY1cF/Yhxz3AGSXnPoRsuq3HVmOn
3fiCqY0XWTa+75Fmv+mKceyOG+6XD5i4Tux1yADSMM3yNW2+9pVPa931BsUKKiw+I0w78sDj4lAP
9gE0aUPUFqndru7Su8RbuiGOi/PmWwlhQ7o755uXjmeJldiLiPye6kN2R95MKxLtsPowWHNGU615
DArPZx/L62q3qw0ercuzK5lEF4cbm0AigxeyWf4DdVsCL4L0a8IhlM07FXd085Ldj4Q6HxghQuKV
59OeSytH6NKalkI3JzZu2tyvvTC0yhhwfYNwmxKEqlsUVUXSYfkWUS1h/18QKJ0bmRVHNx9qRZAw
KEHD3j2O/sKVSenXfsr2FxN8MKH/i52rP4+uVaVeR8bRJWCnn84DvMNUO6M0ONVldMUWJmeOHhuW
2bqkSIdlhNtTF+mbONucH5eeB0dpXhl+t9fUGodS2g6LS86XrtqcIhh+fRPH0mLhkzFcl5oWVXAn
vdFjIj7iM28CxG/zXjPqiFTwYCz6sNYsFOvtTsMzjoljla0w3RLLsiRc6s6Eq/FoCVSqOPuedWr3
ptoY+wOfsQaX/yVJMdg0YhG7q06ylF1bcqLj5nTXxfdfgmzON99LkC64SEGC2B+nGzP6XBMcWiQb
D2K5xiicv3HH79O0EgvgNsenALhMsl7qJzus/LvM5zxxxWF7TFWJePK4vc1Z8MMn6LE20ci9Maes
mZFe1zZQTb10q1XhYKjarUFgo4nFJbrVhkzM6jdhGeh1gMKLqr0pp4g2N0M8EdvFFEOdFuMJgWgC
GCOfW4b6v3ROCgx9kFAyu3rnhk2tztHroudBLjzOpfGlzCFDe28+Z6O0RR1OQmf9ZrYpegArD3Vv
06R77jrPOe9OuNLY8uTpPMXgM2bMltKBBTn6Fomt02GuRc32Yr54LnZd2YGcLLCck3QAznqRcouT
PF//YdGbbqEUSYOBEzcFdkSHh0TtIDxymL+D1MZdcMd6bjEIwDOxTg7QUFvC8bL5Gdr75cDU/33j
byPmKuMk8xAoMnYfQ5Fw6XdQt0hiCLFeFr3a1CSecM6ZNzPCwGEXqvCInaA7Ek0hgu5Ssf4w5gKZ
Hu9lM4t+UYlLfyOJwzLlHJjA8Nm178FCIpxGwEsDXrvx3ofKTPa9OBjhBRfRgaH3KsOc6DPnuMup
Q/QfgtOfOpgf9UhBxJZUxqIr+Ghvc9v15XN1rZiELJfOcZ4eIEzfdPLanlMqfdV3DrD3nYCCjizF
+7XIY5SlCNN2bfBrwluwlheMmxds7T+PaCmHxQr1GOpZEa0VomKSzH6R1ObEUASoIszACIGT54My
GvahrDKdTvZ3HGX/u0H3BS3NOGoQWkm1Jo2jJEc5FUU4KsAIV/fl/W5X9w5H83c8H0pTY0OFFplj
V+9+W1gHlz2bo/+Sc6dL0haEsJOTCQ+LZ0hFgI4T2oWq12PH4X2yV864q37niJB0xtthQxjz1XU9
oFeR0UGXBDNkz0Uj71mnHof4unVz+1/ONY45VqkPXSBUFf7CuDh47V3E0sFSGKIprYaO1VxGlFZN
iepU4drJmoCdIrAa3kbN3eq1yugGL5madqIQzNlZS3ULtdwPsnHB9a3cssOs8froYfcuCM9OfAfM
E8Qdd0spA5p/PcjqEQcmhrrMmCYldgR6pif4etE5TgzktERJc35E2xYLpmq0cVtjuNo6m8jD3YSh
uk+MQqkxwCteQdcVoE3v4IRNApEE0M/DNqJr5ju9dkT+0De2cXTqombaKlVrDWg4vRh8ES5v3YIU
mB/8xFjPu+7HENAT+aT0i8uGQOfmCWE33fgtDDX6bq+51/MYe47lOA6iiLroygHVBkKY3lXRNp4B
CiRF/ulOpJtX3bcwV4rixz4AW9FzySC8QrpjRZKhZbonC8UqyvAaqMFhfhu5UuZg1hbiSm/z1CJO
DO0eXIMuTkmMOcoFguAt3VINw2HKtjirXUlBwEdGw3VLFhG2M+0EFdMV6xBJyIZvHmLD3zByKhND
kmNYq98BNDQaUB5f2LaSGOkTl82/iLYQkRUlzD9gDY9aGThC653vXJfrm4fg35NM2SddY3lXK0p6
CBfZEMMerLaQAONf0/GT7Hbjp6ReuLJhRZfJ/2c5aoAWlyYuttv4VstW9aN+dYLJZ7NYZm1bbq/a
F9x7mzx4D8/SUzfDhXD/HG9FwhJZ55olmuKoF0hYyr8tvX5vzqU+9etxx8uj8t8yA8oRS+SYC6/X
DW/4cDwuLUh3zCD6WDSt6oPLrJmwYUg9H9u7Fsv12eGQ8NycWVIUFSb3FtJGvMntBMWsq/Zr/w98
gpy5xIPzzl9sB5Cu0n9fcVh0zsqbR4GaaP47J/CqmoG5npUhByEt11Y7wrHpPTT/3liToD7O3QRb
Ha4UwK3Uf3iFVfz5Eb715qWlLInwstucM5/NGFgxxFBYyMmfPDIe8JeNV25cROEvOEuflfDjwDEZ
LY2YollbE4xpyDtWcbcLj90fW5zbQXqVjYH9tdPvYMtbSKcL6Mj0M8BZJ0QSsT1Sp/+RGZQW/Fqj
jF16P2ayQWC9OA4zTZREYLL/khg1LYfBv9K0eBkTuICmm7mFXLustOsSqgOwWUSd5Nki6iXRdQnY
eXXqVEi+N4199K3KRJKoMfYRY0pLZpN9efwnCpUuMKei1/Drjbe7nsIZiHUbspXea2r7hIKO6qcv
N99AJWxMepvBdz+RF4a3cPegLUMR5iX1j0d9K5zfXKB68ITSktD/OzGLecXGLZly4raUygJx7l1i
q2oX+q+lLoWcPAkeKUbMkpCD1q/Y0VTSDGPKMIX93N+TQ5FuMlGOuSzvngJaovnbLMyC64pGuINY
cz9B4kh3t789kkYAZgrug4JSLcciX0yZERqsafnd+bnE8Qqh5snOg7/wAVWnExLId5MuVZl/0SI6
D1TyBbWDoIf8glyxlCBo/y0FaZcrDbOM0VyFrzKIDbkDIBXLlWiEnwN0KswJenidqN1qngHqEE7W
VrQNWmZb8tZsOZgsl21BRPGz8cEmB1CWdUBZjK6zzbJu6IMZFCJiv5a8cYm4jHMJ7Xvh2HRRExEE
anR9NjV+Q0YmXC5RfojJMrGpx3KfBknUXYQ4/3xCtOZRn+kHEBdn8ljSi+XHQ6LG3P6EDUNdvtdi
HMuxWP1y7EwEmMK9CnCCbzKT3Rj5E2IoEWBcSKgbK8Gaugf5QM/Mysrq9OOk6Qfa/+Z/rQB8Kqfa
j0Ttf/jfTiWg0eS09U+FVJdgmu+sP4/uzMj74NST/1BU6TqVmneleSRlUYmCd4g5ru4qFJ87F/kz
K8jPO+YhVtG1Ct6PlRsjFeZ+J+ZnUqgy6T4s02+J7JAPampKrjlUNwNUmFg6p+TpUX2hIiFjEPDZ
3yjGd5Y8X7cu85fxRVL85VEVbhVWWg24D89AKsXlPVeq40kEbl7jaI3x0QCwc49b7nolv/drE6Rj
TA2+IKoAcdlxaYyGWLIMNovg+dIaAs4mjgE1jVcykshbUopca+Yw8514GuBnhw8MEHdCc2iVSYDt
iVesQuZz0+RYE3YQk9fYK6Z94z4eiYJ1AzlX1PXZ4mJ3kyhXNBkMJ8BgI9WAmxBOn/pVB34uvJZv
vjso54CndXDoGta2cNEgEDZZgYoekonAea545OptVu9C0XwSF4OFVLjxLY8b+4rivSVZsQmqGuJ5
HIYAh1F5DEpic5fzlqguBf68FTAAMFMS3bNZU9FqRYeEHfCM9QwXl6VFTPlhYPjHkeV+PL3Toy5b
C6VhNEowdXHB3njz6iqviBQc+P8MSACq1qbcCLUCPTyO0fy8hHEc47O11E//UKwcfbbtX22QYD3T
ONtK2MYK/gZA/HFIHShbfgJ6DLhOHOFAj+mxXgZH7v4PQH7mgTY5e3agBbi2lk64mbJuR1gXRzuF
Wf1bjGJ4t2fmfKWOSfgT6GbX+oLeZoDBeV4JPWGV2MK2y7aKFL9HMviS9O8WaBnt4shaVzHTpUrU
Was7NRaWnNi9pz4t7IFABMCr1DwEFV6cOnYK8MRzNfq1LMJh6TCVtqvm+WGyw9CSSbXf85EDlWpj
JMgQjqZzOnN4lKpkBQy275Ba4iOIvZWzLT/2A21xkg5cpyGW4nRew/pwzXGep/WXeKN9ZjtMzQp8
XffpCm6HLkmC5FtjcOElzXR0W4pI0WbUMEARahKlASNohgXe57FFUUJOTasYmpPaavbnk8Hxt4El
wP9HHSW3SwlaSc5pn1M8pBDpBCjQzX5v+zNE0idyn+L8LGZx5TWuqfnl6TgtBTUTK9sarhw7z0hI
P3hd3QflKuw1RMOqHYjdwnDP2WKOY6OJVfRKoEQgE6gMSPkQ9SCn76MmaWwKePyA29DBA6QgMXsX
MZVlkVGOtXnoevkVTzDW6CGsIqHd/d2XpBq2LLiNM/5WmNjNK7XLzEBMy9l/NOklOfWoAYZCFM4J
co4pyHfaJXpxCDaOifeLkJ3+9ERU1UHCGPFbn2pz990LsLoZ/c5vLjBHL2o6hzHtwfcWN3Fm8s91
kMqX1WI3QZ/WWz2Qm4hbgHnO0cu2MToSEEBFxboOlwQ4KxViLs0i9CUhN0mJ81sRs3krpraV5k1i
v9bq0fC/oB6QSIVffMwV9VCY87G33EXMcJbl4ezzJeCZ8z9AWx6KflZ/HL0E0eA1XCfaQpVthVNv
nN5UhQ4oOQY9T7jr+3zToJMJnCjsBvySqXFnFyIG017JsayFg3gYpz5g0k3lTKLDJUTfgTs0MQx0
C2+armLBeEiveMJz0eeA/OMK37HAb5Y+76zWzs8/Ob2zhQFJAN/cclhczVO4vmdE1nq1Wsnr4IhD
KRkqG4YXyOA33xYT/35Imqpwj2r5lSB2fow89gVgwIYpYsRVoUfpKZhOjoqW2bM4/Xfcp3TuR0bf
87mPuwBuODn9dpvQ9maeIOhPZWdRngJYvRhgGbgw0MdpWIqLPVWgYR/lhY63eNnR0WtDufBEjrY/
GjchWuzewDLbbJI/tD4RIH92Pz9Gm63ppt8n+jO08cw+OJka8k8ri9cP90glgN6z261pcpDOYW0P
5Ahu+kmJYIsQT7FxufX4//7Mm/yDCS24OR0nVR68xgY6Z2lw1eJw4oNP9fqQW6JPJ5t2e3DNdubv
ozsL+yYoJak1KHt57Ys5diWhQsDBAxaQDDQxoQc5TOojHngF9qMbudH/QIJqPEwDJ2MWQ6CIBg9U
WRSYwIfcxF8LyunpDQFBPmwZFbTz2wDOgm3VxbOx2OgRMM+HKY9+qLFMQElYkYTXIKrK9SvctgQz
/79+9J01c1EwdvuA093jvZy3qGKTzr7TNrg/uw1cg3gIag0ezP1pa+7IhdjAyJf7wUjmRHL6Rw7d
GW/yMkZe0Agqr9t8fC+ijqMz6ag3+VIGt8xcU7gnALr/L9Fojy5D01wowtfoN+q0hcHL1VbSlpCy
glahmUk3ur2d45+N1O0H5FbfGFa5gsB1r+t26Bm3KkGR6+sc69ViLweitmvakIl+Wj7eoO9ko/ky
lAocsed/ZerIPQ1JQiMCHVh/F88tLX3lo9Pn9Tb8fwx0kqiW5fdCvgk+n3ORJ5rl++aDoyOkx2iJ
Yu+4zOZRIYnaqAMYVKXn9GXcwq8M8pipzxoUuGR7Fd92uzeESmmfIDV6+9F1y0pBxhYj4kmP/m0F
bpazatDkG/5OkrLIiwQDBx5b5MdwU/sjZIgamOwwOHGq8TxYJFZGPyAs8qJf2DqJe0/1sU5r1P2x
yEGac0j6nJj6FKU+K2Qwv6qo3qTkQ5sONq59DE58/MA4x0hxLlljdD0YK1RWFiEgGqXz0Q9CMW5X
yVE5Tu/3EoNWLwJF9QXnoV6Tv60mG98vR2B5wnJzHRngbEqIORq/Pl4AD1JnSthvcsAmSoyTHLcJ
KElpUpI/ONKm75nfzw78Qkjw4KUQFSNbTSqfKwAKgX5Z815Ygv91D2UTHPAbwBSlBoyONm7e/sF2
SaFUDci+q0+6RMJq9d5VUIeXuJ4+ZTnMud+BqDm6AWNeKp0ejGpdm2DHC05mHZ8LfvHRopLcpjRo
4mXQBmAXyhOtYvTCjb90NiykG6AgOcHEwnhja19RZ6aJHaBN1ARllu6bT6v7I/HW61j8gwlotCWM
6SWGXImdL1JRbZ/0/KV3JUxuaoB3PXbaoJZ6ODLfweQ0Y3nGDAWMd3Pj2bvOZ9cu3UW8IpFJWPs0
HV2Cb5PS9C9CXRgcJjDfzOqairK+t+aEGmrG9ofYAVSoKn5AucoXs+tGvcXrfbo4gT+9lvT1ObaL
gwsqP2ruMYyyZvlpnA1rdByCgmD20Ms9cPtsb3xH7d+vlTCGXv9cieYSf8/aPoHKgmsA9kZ5XHry
kowTI7pBCBLZ7qdbdVib74sa736G7Lur1mjhWNFZ8vIxVSvv64A8t3qRQIlekFk69MI1irP/y0yt
gz62EfZna49G5uMIqBrmZcY0Far6FzdCaG3y4td55g96zcUEEdE+Bf4enIfofiOidIoSk/N9oFR0
1waSxeOzcBtAn/B/dTGHVs1BKcR5BC0STdmLz3YrzyxSlOgQkuAvFHpl7QDP+7Ktu+YL5G1BKBOX
Eo0eLEXPzS5UT/J+Rd8E4SaXG9xo+0N7ebgGVDArECaNxbEZN9IBwGiSn0rYA6Ys7gf/eGuphUNP
vQxTyGDGQm2GjH+HAokSi5IYPu1vuiWeuOD/tyUUe/eb4KcdKL6RyBouqxhi4VoAUFON/L38h2hR
Ag+UH7sgU8wnFkY3FgNUY9JTZgdH1Npy3bDtXGeosMxJKRVT3iNNKD10wam/PGUJ1XkLm0+Ttdvc
CBMOw3ON2pcy5p/3l+iiAmgoDMRgK1Xyv7MlHo8bxsSvu1kXoYQLtoe8aaluWfPU1spnMDkhRdfX
0IVl8ztuygFtjh2pnMcz0IIhlIZQYmsZyzxHSeULOp7wfWBKHax6eR3GyI95yI0wUvG2kqd4lOM9
jyn4pnrfALOai5uGQexf+X28Xu7RVKfGBf1vBtFbFqBRHSHZPWqzWKVzGdERB8IwKKRS3KZp3RvN
/tBMRAvrdD8+cllmZFxKfCG0oJS4fqdVrYMpRCf3YiGTAMkUl2heY6tRReWG21cvfQ8WqBC+yHIe
B/tROmXEkR5qhGaWlcDg1x6NMyo/GLp9ylJrThCvWOrNkIcAd3gem+AHZJHi1wQ1Vwa5cO9dlcGK
ja3l2CgmnusjqoPLwgD7HS4sDRF4YgOu+wVu6xOD3PphQbWlHHTs1axvfch261I0gP4j1HACfwta
IgYSsYw/BzZm0/VYLA7d1d6r8Q55rQ1qpPT8r8vpO2dQ16SR110KZepTGdFsS1diIRAdbhvjrj2v
C16RNPiYox1xoFcjE/pMOshyp5yzhnRaMKheWSCkW8rL27XaqX7EbGFER3otW6mVphTVcUked8kt
+RLNgpDBG7V9JJZQfzNDmzaPQ0LUOB0PYXDOxJbr3Td6NTfQiLrxwymariNejxfh9fuB2OTkiUfu
ApnSovUEMddWBlvagqCxXSbZH5wP3pZUKJ6EgOnOfgJULMVEodi4pVoicbCfXZdRlyB2nzkfouQD
S1sePDR7bNeusgwkB4mjouE82aHXALtCB/bOcpChWX7nWPfTxwYadt5LE8XImq7OAoBrCDO93yb3
/N1li/dxCQCBFUTRhfR9uCy7539+Zk5HMOx6jN/j7/dhPTif+9YAhxLwNjT/MzuPf5zu+os5AIpo
zQf467jHMgqEdJk2Vi0C2EO6HRyIvoUMPLu/95uAJgV27F4nFSsuewzaFIvQciH/V3ylo5dqwY21
SNYTGyDOtP/ga8kowA6xrwumWnZudK7F416OsTgDlRn1sqv9wHEjvRrd7j+/EhdkBqFqtxPU/4/N
HTbPzgyhTCaNiCcIrwBRCUfn8UItilCwTBKi12Eu2j2aNFKALM7Lhd+F2gzNk0ajdZ/enVudcD1u
vFbNgkAYKADIgjkfcyd6Ud5UFhvw5Xx7QfmZ0++hhpAtXyytVhqec+dLuiDtQTZHL6R5+PXS1pU9
ZQMWHcDX/4pN3URNOz69eRkJO2Xn01pqzjGMsmZMPZ/pIqhihdEYNZc6QvvbUGD663TR4mAhJoz/
P2RhWlkZ+3M5fA2JvAV1zWFkL+fEtxvaSR1+dz8Z32mP51zKA37ILbfRAxu0OZjV+vpRBxo4/KIb
I0JDja8rFipohvBZ0C5+CDU8h1lssqUUGs1zWZJrwTeRRGWfPqHNwuPDVID+d7/tZ8TIxA45hQEz
xERQ59SMfP47GIZtgATjN8H5bUO7S5o5MCqAk12xHiBaYfUC1reXm1fMhv/mlgUk2Ts0sZw/gJgX
gs7Ryibxl+q9bJbG400PK1dVHOm55LZkaISZQey45Je8ucF9fMrYxKco1W2GxlajZRGCK4z2OIOW
w2/yCz90t7DVTh0QppFHEHEmjUTH2Rj9SwUe/hG4v+WfGq6SgQ8KHscxe8qY+YBVj98MzB2HIo9V
USqsRpFFaLByz/ZGYD7ABhUkhBGenxk1gbKGzm7yJkNxgADF1Uv22eKLxXU75tuiX2Erp6VI7RBV
WqQ8VgnzbHHGsyvw/5NMUpGwG2JXtC1FBi/NnvFEDAjfCycxPPUEporIZyFRVpPOBFtKr0HIbqe7
oKaDGrGMM2CvSxcXWqrY1ys9uBbzFSTqmW8QN2fsYldxjlBwelde3YQHKc0e69J7Wi3ynSuv8Ykh
u+KB1lMkCEt1iju4Lt6Xch/wuLVQhaCO8iZ2MDTfhGWyzHDdi8yBvpG8VZS3GosrO7PC+m38G3VM
SJBr6ib9B6zBbfNYwSQ8vDOPubjPfksyQIiKi4rh39ejKuN31bj7YCTs+EvU1LnC9AhRoRIMQ0l0
k3IKSIAOzX5VY6o15G80kzsAMQHO4ctlLmhS0LkUlmmFJBim9kWxE0zjxZMl6QHoAyAYsvYYPzX1
jnuAnMcHtJLIGb2eqdVeWy8j86Ipl4W+NNvWT0KCTlIyKkqk3WpzaUZ2xoqT20N3E1+KasBsuXOH
dsq85eMxLIUkH/86pcqmlC2tUZwCSDwyDYY7/hn3aj1pfolm0KGOcQBJnl5LHrno3rNxXbyvqdT9
90GT1QMon6kHhYNjDXMh0mYTu7K8eRboTayxNvmeeQ5TfLm4+LsH6r3iwkChcAbYgiVUcbxz7miW
OWCVz4G7zC/0xWqGFV7trZWn/OneadgqNlcdTSRVPcm331yhtHPfOVeuXEbCYErjuRrCZTVd7f4I
/ys8R2995s9wMzRY2PC/fhoUoogd+rfDhmP1O9SVzSc4qBljsByirphSlLykSJ4X7kNUizy84kkh
uYIS9Ls3bC7CYQF07Rz89N0aji3Jouv/mgt8k3nsHgLDVZBYW9FQyafymWPfswTM0reuCzpmVkIE
adJ8heu0XtDuUcFx8NgvOSowwis+7vX55X+QmH3vCw1QD/+ZBOTJEcyLAOpLahgkAuc9Sfgr3b9V
1Z+wj1TOH2JA2Qo4ruVgWGNRDmWNRJ9JrcQIFHjJ5bBdfzftrteG/mRKZiP/tq77lsehYJHl6x/s
iuCI0fCTnl/heOYjmVyJ7PRZjls8oR5viybMbRFLw4dx/Cua7vpVHnpGmh0q81LHGoIHSdFJUXee
HaGDYeqf82PlfpROIJaWqcPHe8xBWzrIRpc4Q93L5w2kKODONc0d1yJpku3pwEB+nZo68h/bLjNV
Wh2ef/wnMTDgAkI/yJ399lM7UJJJsOJu1KXvn1DPaAMTrQBstRUi8lsN2HLOq2ww2WTNo4NGHqb9
sflcoc8qEOfxmZrZMjDu0ylzClrXhJEXfREA453uzdFM6OYo+ONitf44ukH5EWfPF0QySAr6v6N9
fW3r65gkn0gyl0hD/x0Fz5JopKLdWSAQku8tzDQMoe0g+5eqJ7/MEuBxK33QgLd4HbqqOBsPp7T+
k5Si2smQ4zX1kHsBgcV0jLppge+WhLszO3nwvyee+Hw2xdviD1/I4uQXwCr18AcAWzu4xB+Suku1
5XLWtHfEtX7RmDUrlR29ehAaJQlt3Jq5QIBMwlDQlx06tgzZfhCS2+zsbOb2PDnUo84pi9fHeE3i
dhg8BrPxPcymTBsI6ejRZIonVOeMzlemZWs7ifEYPgN491e+Z4D7CYpuMW9dSxdMaBDFxfgx1xro
2tFSsATrrM6qkcXpVpXZSVXd1vkJqECDu4FxdISit1HxkOfmLSr2xC+RCtzbGU1dyLaV91ywpNy8
Xs/Wc5Sb9gj0ySDInGADJctDO3d3tSB+yBsPCP66D/ER61JCq1RLu/9sAY0qJVxYGWmIGwWwFFMl
Ne++RwKgm/npTb/bWd7o8ive52A6MqksX+TCyRT1Mq/FhCOzIc2HJ5iOWYobbjtKQYxkhgpu/KnM
QR44v4J8I7znQ6M4wIDAMkbpet5MMhCren/S6abTz5mfh4DxOcYnV4ei3sN8jVl6oJKx+IpX4GLF
UCIW6qSqwtP1HFqsVh5stn79TAzt7E58OwNFWwXKxZ7qb9mzFCRIaKAU/KGrPabB+ma4YmQYdHvK
russSk6VDn8u/vNOzdxILIL+IYCwJ/HN9j54C5nHcuPRUryYE+Czzr+ZKDaGax1HTHOmCN3RlqPE
xEBhMHl6/qBqvQzsd576F/6g0R0n8ot9/WvPNv1NKoPWOpHn1868ozLtAeTikk3rio5tx1aLAc7T
eeZU/vvPLrV4HXW1kB5QIN3kbBluClUfUd36Q6DNUDszO3d3d/7SnVgZqVh62tAlXWBIQi9VZ1vn
6WxbpAjcr+BLf5Oz7oVmuM184xFbzXUzLQ9vRCcakU91p/Xoinc1QzGdwYKiVWcWzN7s3A2oZgyc
2W4HCchxfxrhMuh/bpHu6G+P8RRkMSVpshRdaClu6W94gha9OeyZIT9C7mJL2sItXnd1X0S4cI+c
peJAlFp8iBVUv5mC/Ope+mMmG3Oo/OvMuwp/8oGvHAYT5+oVotgMcBDv6HsMQieZtGglfM6zxP6F
ouNHSlYREpubKf66x7V8lZ2pleDskFYBgswAVzCtdRwUOIcdAVTSMhVWvAsj8fQlRcWkFji/j3p5
DCc95BYK3NJxHbWBTq4eidx4YVKTYDVPQa3vJyIj58xO1h7c60JE6mPf71ZbWdy3GU7aWEo6XSj1
v7cZbBvvADg1mpaoLN+Ra+9JpGxJQP89b5K9LEgIMEYwolMdWJO8x174Qfd11vEj0nIjM7sz8W7i
aiTg1CFExmARNT15EaJy6wwlclI6h0ZM5hey47WmTVWECB/tLG7/HDZ7xUpHjKUv/VemfP4Y6XJR
kbam645F+FCX6hCg7b3OigWD0MZIfU/fPFRLt33RJMmHAspqnWY6olEFHAIOaLN/rzTPeoSMatm0
VA9dczwYQT+EoZNFqXwFlpCjfuLo/9i2aPiHYLvaz19889AQ+pPYvVUpbbu4JM/+i+NE1vHEyyn3
xaB1eZz8jmPBpwmD8ji8ofpDG3X7PmDO8/036iTwl5ayY5vz+BCK9p/gKKiQgJIEXIlYHghhY78K
yatPiScZTEa+oF/f588XmH4C9Bm4oiyRm8qt3Wnt9NuPxMYnfj9ISUUVT25Ao16g7OVJKcJplWjL
eTQEu4x86EoF6FYXfI2KrVMxll06pq1IwCEBC3GpKvzb3nGVLoH8/KWbb3TrqBcvOiSfl5D0bKh5
Fn7HDcZnHqeaDTOnQG1oXbYQbg/Tl988jiDlSyCksFPeUnY559r3DxeUNvMBxC3PHU+1Mq0HLEHE
/QcqVKLfLmpE6BszdDoi36ltH7hjd59e+nNmsLa9KfnS2CQlMfCvGTkCeAOYkd/jizR3Z3X/L8Ga
eYsKt0V5JqXtWDz4fuqu2ujmvfJMuKQgkyr8PJDpY8M+Mz+uDYFAnLFtKwGM4G29VpdRRTREyfE0
tAecKffJRiBqCQs1iTvOCB1n5W5TXHkrS+OLXmEnikI9wEeMzTI50vGoysBmqCGgy4hdSxi35htF
t023rpr35s8T4NL+RBWpkov6RqPyK5rPclOe2FOvj+80pd0GYw4EVHqoDrrCxWLpVDmpyPF8oYS1
WVjZIhpfCAbO4t+RSYMgXWJ+7u31rFr8kiG9Nnp8NwdoTfJI8FAk+rfiog4AXMxbzdu/pvEzI0NU
T60KiQ8OzNEJ8f3baN5geWSdHS1pUyikEH4TmOS0OcfH+m+474ph170UQzfPOYoP3+xUMfSsTK42
Lmh5c0QtVhTyWS0wIpu5b7o1CRt2ngKuV6N4txIK0s5xdX+Qz9Gg4GnFN0g3eYxkxgeScqXpbAIM
S22OHAOaw+JyRsu6KMHbBLRXzeThgyH9GytSMTYimaGaav+uEG8aiGMm+KJtWODk6lri+Pv9gd7+
zKgUIAVByQ2uTl3BZl9UOswjPRUnMpQGNPx9aiZqPHTAk2YBN/mwdHftsxSXWjqruTRjKhw2EE6P
7RlXq7zTtn2+LBSPScggqRdjstoiLWm5glRRbP+c+kNNt5z/gBExTPiseLQOWxF7bk9c8xC4RNeJ
iidw5NKCs7+N1frWEAMJJ6pATaCOxCCKZYTRbHaFzgitKFZdXQgKj7PIGc9w3fqqZ1hLdITcNZRw
C0v4wE4ULepHdgkbARRgB/8Gz7VQ21H8NTTfabouyEx/dBW4yEHVNLFGcubwcR638hQkIKaCpnhU
r3ysPlPBE4zxNC3hnNUdcZ7+YH84bYAJNUFb0wWUH16io4kLk3SwGeihMCHSpg6+epF0zfO89vpQ
BBTxc7wdaF4VU9hpmTogI1a/IYlCBWrqUI5vEs5jpX8zRF6VR+CN3gRDnVDmrMMZPMHpL3AGsf9c
dqX4ZwrJf/Ksd4yNhsmdZGqMCbt47Js/gR4zCaSHeuh4tbZflwRY6HRamRQil6YWvtxLthiBv+mD
3ZU34Z0dWIq3p3RtRSSSJt1rBLMQBSaKROWr0MbDkHJyylPdAt0qaG7V2inuGnvjXrHqPZGFn81c
JX7/ElErqhMNSvbraHvVrtU2N933L/7fjpLr7kBPRekiffOvj/2gagz7ls3DSGvimwcg8YkOX+Ab
+VYWsdBoe3A3Z56qJigsA4ZZk5pxCBfjEPFxl0osHEm2W/NZyplNWkN6t68l7kBoATmy0GHn0+kf
KzHPUXzS2Bq5CJnCJKPBnWoWtBfHIDz8/K5fLEBg1azPRNtUTi2gRaPQOh07hI3Ft9FoWvD3ps22
nu7lyQyeBDitGkYKPIipGHyufYtXdoGagZcg7NF+REgcYA7K5WmOgeaasZvXUhjV++0SGlqBh9Lc
MiCJhTpmYkmPeesRyOsx0zTFj0qG0lymmSuD61ftfOGw7gLn71g+F2xAMNfZ/S3nfXHTxDsNUuv9
gOCC7p1tpx5jbFsSzMedbyiJGnbdKDkHqGDUMVm7xkHVpxyZf8OhCaGwhmkble26oE0jT8GRfKvi
0hp7mnERVTRBMyzPnZ3hgYPvX/hQoX/I4gOzyOtHz2D0PnvsvruzV2FB+bCRByytIQu6Tz9yjlNY
b3lfkjYYBPZt64ZhpovjU2nG35hNM6Pga3ahT1b0mDXnSNAmiTKy97fMOBouYLq7a0lZFAdmfcdl
ZGphyvunQQ6VaEijIx6pQ4T6EV0lMpUqaeI//nRfXvjZ0+2+de8khX636sUYHB7cDB8nRE91yNzV
7DoKrpF7DhWjrbJgcp2otHfxvrCjxcNgk9sKiJYdcsgIr+xzx9JQQDin2ot2RFl6EaFg6Ej/2AnV
+ria06AHZu1Wm3VjkOWnvN17DH1HHZNdBi+FbbG4uTQqo0b+9i5OaVyU3IaukVYs8Swlnflrfh2A
wZTuuJT0wz2ijUo6kYU0XoC2qOMD5jXvHFQF56OSEO1cGXMm9joDBeV1Ybe6QOZT6nJhqJKLIgom
k5otnwTvkMWzEu6y1rmbKKjlAnFsGNHYVwboc+r73+8cfFG1p4IgkoBX+CAvnsObTd3Tvvkf77Fw
Ga3vIEWwLaFbVp2qIsa5/iJKdXSKPscSi3ruu71mOv11uN1HSV8IfNB3CbjZGj7GT1bJ4izXd+NJ
mweNzCqLPWobZWdwiegyfF/e8FUfyLtwnP79twe1RKY0VKa/ctuCZfT+xR4LEfrKU+XYG1RUJqEi
ZN2EGafiBduTCfk8OgYVgXW+KSRvGGTkkqwTy8uU7e8ilU65Vv0d69L6Xs4q45eDqxm5UqClbSGg
oz0oK1HAVIPxRtFX0h9Sv+nmqcFUZNV67z0IB1tz+CDBx6Sn00vI8uo2W+rHZSZ/fjS9StpTBdbc
SjSt0pgjwoZU0/1B6kD8FxHZP8WW886YxJKK5ZK+Jh5A6SD76HOIbKLR1Eb/D1dalaOOm1ZcqxcI
cPVg5f9JOEFd3UJsIA4j45evdeHQnIAlz4MXfo/MlIqyKMncdGMOjMN14MkZiG2Hy6fu/MJPkMx0
Sg3hXHh6rDYC8NgT/TiMSBzECS/dv+eIGWPpY1wveLt9JWAnjQ0pMA8h4fpBNPS21Y6In96jmEzd
464/6Usf7SqLWQVaU8tUjF+ToKYx7mrpvOCopmQc9RKb+WLptAoo8BUj9XZ96uXRbVnhxKquYOj1
CK9FXPbSG91y4X6jcRuy/JjEiyHmSx7XKMGz26/ey071qAoYVINoVyusMm9+HPEGUrZ3IyGHORIC
IZBRDCBmjWJ9Syg61onvccAC7/d+6m9Pi/eWtEP6aRzSgeuu0VXXEzhFcNWdiJj1TtbJEcIoH9vy
LNAmh7ylAVB1WLINv9Zoa5RtdP5sl9HYFFEDtAIB4XDIx1w/R2gUVP0PeWrX8VwGbF4QFrTY/do8
zwnne8Oee5hhxyYYVouAsyC1tqPRp3tytroTkJqmBnLCrs5Ei3IsYC7Jj2K3hLLP8IgTb6RPqfGp
uIUTocGEYA/JlSTZn/jOB/3/m+M0L0P4JOVTc/rMomWvnYRS0xInanVenMFOJxRQFV2BdSQnt93g
9+0jjteqF3PZx6cKozsLoWqLDD1OaC3aXbnazJfWCP3IhcSqBGbYiED79EiTNXUqXjTgspxA4pcO
/0wzuz6PUceguk/CYGGNN8Bdk7py6Aw7IaHYpLrW0P49ipM2S42XVNB3CMUD3ps85EXy5jxO8vX1
T/RS4KG5kCikOjVzYa+FhfdYTGC3Q+Keyfl4ITohJQqtEBDEDeJvPw61lY77LdYkb69/cqJAGjls
omdF9qL48YMDL9SzWF590zuXuvEnVifcVvfx0iMJ91eyzmOuHO0S2xdxI4nb1C/BSlPJ9C8haYxU
kfmoX3c6hgixS0MNQJsMKIZjZFp4hbl0ixjafRUsHw0HxGrFiEnWpK/ajEaPtZ+mOJO8WIo8EXTL
nwj+ppaIthck63hi2RSodA6EooURE2YAcFAHiAcl/7AmxgvsfOqZuwogNEJuTYc57gsztYku8ssv
tYMrHKvpKZ71/3F26DHsQaaNoeq8IQ7f2t1G7Mx/iCpifZEGQmXpqAOxhdScMX85VN7pN9PRzQTo
D/q9x8jvlawKQujkdDA2misalv7/uOF5ZPcLweywP8kv3fVeOtqu5HOaivCwOXVq3w56NBNnILOf
lKwFNlyhvby2T6qD4iOR02IpwWCrKHs0JfaQ+3vqCVmq6v6sMmP8ZYHehj4H3pGNz/zrDfeAeFEv
H8oY4d6nAeX0qOkLVqX3eQ8PW191ZrEzGXRw4ri0BiyYP4npOqe7IAbZVbHJJEZze960X1ANLgVO
5mV9bu5PlhKoMxrZw/aVg38X+CnGYOn+z4EAzGolbML+YAhps8XPu1SSeGi07SxhKWZYkjL9uq2U
n0nrT+7dx2OgpAQ6ygqw/9WkIwn3chrHYK8pZuhg0hVa3LHqhUIhtsoi/krYWChCkyzEUWit/6Km
XGHB6p+JhDlATbBBccC2hI+Lhx00Bvr7/yU8X0/JHjHIyR4pquhl16+a4pOV+crXH6LToKCWS1YJ
4xEfv5J6ocLU7sl/9+8z2Ebo3cxgtngdZvF9CvDYY17j0m/XNT/0cLS0YpWCNEs5i05bueGfbJ+V
P9D+8WHMOww33RqnSv+r8r6wKxmH+gmcfz0RKfpnKeHL/a9fYOqSF82CdbwVuDX6OiHdJyn3r8Pj
Gcdu3WEAqt5y1RHF2/fKD38oib3bo4vJXL1pu+2BAlpOl2TzYaQmy8/Fd7VyrVjk3thYQXxlvzDG
M2kiPJtVsTffiXDB5W4Chmzjf22WWGwoYx1IJ4uIB7VTdokO5bwUW8uy9u0F4Bq7gt0UUxIrUqQP
MqJxIKqyx85bYFmU7PhyUlNI35goXZXuXihzAm1FD1jaBdlDaQRODS/7fDYSll0nQzFBGDO3ohpL
9WLVOhmRGIs3KSZmVjCRv9qNlJqIwrw48LEkeJ3B0JeKivUWa4hhJtAqpeOBD6qciotNfRGuD/NM
iF1NkPozZCWxPbUpq0Y15wSJle967ktPjGI5fwxWFNfv/lM1EsB97osmbcQKRuQY2oUlzKxUbMLd
dGkTbEeijo2ZCNtxusuoV4p/Urdrr86Q+zlIlk23w7fPYgISZ2JyNqU/Vf0BqOuYg/M6xR/rGROl
YiX6GPK9gsfuCvk6F1F6D7IEXsDDmvzlCf5Kiduhd0oO5ZsRRhjSiLuPztBXdfFGtutWF9yjYLxd
E0nPre43ivDqqcVm2XU3zhC6wcaxxsjub7p9voX7vTA5SGNDkwAvyjl8qYDl7WOGTNHwWmsXH2PD
eMRfgPpj7xyZ0qABLLKqXP8ZgCk4YUN/pioDVYpnca21vRFVS50XKyeed8BnO7W/AJ/DpU+NXMWF
Hm1dpWak90l7kuziCGxTh7lzrSSGRW/MD1HRcKAYg/1Eo5XtazmUSCV/fKC89mMf+jcQIHo5YtND
ZRc/Rr9tdtdldIdH2zGNbteuFzveVCEiWDS55v/+IQBCRFmVwvU9h8EpEi1CzI5ysxyt53ec3yZq
0Y0p/+xBuEe0in4Zqm2gODutp+bSt7FAaQHHip44cRP3YBtwu+CtD1PHlh7/ItK7rROkI43ne02A
/NXM5iKwtpybnEJrhycloU8Ifzs8bCPAiqvytYxr6unnsOPFqE7fh1ixTI4nQY86HePBa3EIrhyl
GU5FnohKg4QEcrAYqhZqVkRyZN/X1Ea0ZkvLpy9OT0I+Ad0HPqpSYg03ohXDBGMIikxhMnjF2VN5
H+oVsQbOf0zTwh3UFDVEsYQ69yxT8BgxzPj91Igcqc/Qc13SvkcOy5mCMJ0MXFwyec33gRy9yFnm
PqCxnoT3c3IeEd85nh64ffnGbnTXL1gO5tThq6/SusNUMwHxhpcg1hR6KBBQAheqSIE9V+rnUOTg
Yxoi5sLbysttTXaRs0yPSGsN/L0ATcytvMqmVsewSbt9r1yDEh8KsaM2zrUiihC2z5FdocBK1MTY
3vd6JVlGSiHt1YrXJRTeIaY0UIdmwxDxZWUt0YXwJywZswFVzjpsuSpU2D/KnzpVWRnI/5KNM5Io
LIFPFSYaZOxSkSbi3dg45H0YjcBSC0iCzZo601EjLiIN2vMeTvpNxgvARAj3YEe9baWlfuC45/qY
xpsB/Q4vIVv4LBxF6Rg6CTCOnYDwIVVzuw8oWXg0eUtQIwopWjuIIkTZP7+R2NOAE88eUBWp/S4V
MWkynogebuJ0WM5EVsw1Pg+mRgu1XlgthiID36MVO4N6+kk+zi5IW4fdtlUmnXOQscIf94xjRq6j
c/n8vQwSgGHk66zjKvfUkgsVyUS6KcMtzpoIlmt+FKaqDQOhcugRpzAkaRjKVm/XBwLYt/yuVRY2
dOS9WXwZCr9tgrF8uTSkoAFqjysFnOectb1BgkxHY4OjU+At4oToYd6ExXhIlIcaHh6j0bkFQHsK
UxrjcB/b3iPulG3qFnwHl8Vw8JV9mGTeAp1Ah9pXh/ltD6F5Stbr3So25WUNMr3vJtNHmA9FmaD2
ClOa/y6mgEh18QboavQf6o+Uj3EGoBdMoB0IjAFRcdNyDOFb46Y4zv+dqCbCkGdUbH7tNSsJJNMm
sEZeGgLM1zjqNpWKLxa159uTK75NK4zyp2hgdZWYqFwI+DWm28qEUJhnqgIYkMzqMXBmxZhY8+xH
fNYKR6gppuYMEUIUJYvhUbW2E90VDb6nAfj6/LrBMEazC1Ek/gUHHIlDo1/VlOwG7Yz8byahZxSB
lLuagG1MlbiavLtv92YZ2UIE+74Iey9ByCGjKJ5BeuttOEtTXLUUmwzb5NswRoM6CNUV9VYQXGJm
oNKcD3XYwIDfDEFVJ/xLUM8owz6FZPVVcPbqG1N7w3EACrgpFGIUmNTteCaULnMD1MXke7gtF+50
LJkwCGnrDjOROPk+Dg0hCyMlFivtyx4J7icRHoFYa/RgsyagZrPFiGUHEeE2vIfP7PN5KO/HykF4
EOM+4lpqcImU9crJKwJvQiHNU+vGqjGtiiUEOIlIIi14gT+3qwUuszgDE7BCQUSnPy98PjRwxyXu
jgaFHB/yL1xK9TAAV8reSFQpoghhFy4l8nJMwugUaDhm/EuboEfa0c7anrVsn1rV90XTYwnImyAw
ShHlZHYIEEnPXd8heqyj92+SZOqtiaP6RnKZN4j6/TAilgs2bOKVd1yhaVYSX0mxc9vhOr9VtBPW
4qpNtuz6DcnlaNPeb2xenpoZ+dIRRL6AYWwNQ3rkmTBLdJSxXOCt040Kp+7gwUPc++HMpRRGixSG
z46ADUO92hgehml3B7AsB6rDj//NGS4mYOZqhMQSlLdQlgcGZV8J1wrz8PtW/fUnqC5ytRZUVmbZ
rpvXuP9M2PYJmHlqReMzFLNLJU4eSC6bxj5DcRpNPA1Ts9eeNj27wwVI074rKYVPbQg4OE7TK+om
3fpNSkOTUME/Aq9dHARg1DNMwChd3ooh+HsyC7BDPyYoEuHQzTlXNtaLrTDmKzQ/ENtiBhySivDq
y4EMTc5BXs4fyLbD5EGnma9+5bkdrWKya8vrJ2LR75/RokFaTUazlyaYQiZMXAJS4uf/jXxyqv6m
YprE5K0PvJdjiEWB0ygHc+Q40+agTh+aaFMxbdaqhVVJ5bNdERrwfNZ32LhQUlxGuFxtCjDo+wT4
8tQEa5aInHsM7s9dDajiEdzHLih94jCxpvYVeGshzq1Py1mQmxTr9ZOsEpub1tX8teaF2wDDS37u
H0RbZkuNH5hXfb5VPoP1OBvE0xqh6SrsVFtJMZlzOC85FZcatoevm6Pqm4AVpMgOmSLpascmuxdH
6HuVOxCoxFCgfdKE7UKOP2TyihyClIMBKLf8f9TI+gxCQpyWO/PwX3YYR1U8oY3teYycbQQPVPva
h0l0x9dRsMScoHVMYJ7Lb+yxDzXP0vgxCvCOZMHn1zbiseHI1G0JyKo7ojzo9OzHxHgXN5FX+6gm
cURinZm5UnuDqD1WzOFotMSQBF12Zyg9Qw5KUjzVtXQETx/Pk/1ZUorKikaZBBgWH2oIHMGzmzMC
rq23OgVOtj7YTmsfhdb1/kqNn6OAX3xOcFwEB+oWWSsu0cugzRCBaXb+14+qb3KesNqBUlivxp06
kaFfkUSGUdog1OqvPtbDGYrsA1n/gEORf/ePkCR1zPpnB9DLrrsHWrNU/6181WRWmuhn6LbZQRfI
pnqIezRsh9DaHvPUxXy899/P5S7ABemF83SbErsmo1/+SARUiPeBhJjoVklcPL+8Ln2rHlIcK9Cw
TvQjLI+5EsbJM5i6qFqis1K4d03xGNhTEx7KbLUGd30w/afF5BQm1oqC361vZ5c/L7s0j0QWPXT9
0UPbt3KNSf0+0jHEnceQyHvQo3Sfz/FeZJFRO/rneridXB8yDuuedAolYualUPE+qlFkgNObFZu8
AQWsAcA9VaI7ic2LdhDaWD+Whga3OozJpsjtidUXOQGCoVgd7x2JO/tNNRDrUi6GMzTptotDVAhe
MdlSUlc9svg3wBkaQwUR492ZKew3EwTFNl1eEsOzC6RuCuX3l8d2GS1QfsQ5znH2VbrPS3CdMIum
MtSWF8ihxl6eQyB1+DLWTv/Y4VKyjVPuOmVFgJH3hBxxWBeyiLgPMYzm/fWYK53MUvOcehj0F6kT
4/d8uwNK/QsbvA1TV9mB2dOhsWzkGoILsqMkye0x9poHiyK5GuIIs9Fr6VFB0oTW1zfu/ZblGLv0
AqOitN6GvVfvD4hN0EiB2uQWjRO45+TCTojASF/TAz0rCzup+LSmeEffnM74j+84qcl2uCiJZjIw
xyUNiqX4vrovigV8BSEOa23Sa7vIm78mJhzwdLWWpu2ZXmcAz8EkOzdtnIZL24XUGNf5y+J44Hqp
laDbiHAE0A1eZwso6AXrE+kdGkj8pfyU+ptZjw2a56DongTosB1aSnfualODyHGJCsnsrYVaRsXL
A5wBPDTsq5AqKE6hnKHR+1ktMZH8sDu0EHZp9qrgIocynvIvWWqngX3lLNLKRPy101VA3RUzhrUG
8CNXQ45puQCAsd0UQAqhhptd38cy/9JpVDk3ahjSEL66ehoCAS1xV3D8jrt11KRmAr85r2pfjqlm
PlzAPDxiUMB8zZTGtn0aW6ewzgXGfpl7UC4Q+PmbsneG8vDjuxVCGsjFLwXDk9LiIYuc39ZoOwJ8
Vq2sySUg1pygBcxls6dXwahE3TNaIj0CBALvOdk21KgseT+JNvfptXlrEvyWltA9LD3fX1qfaTgU
Jfbu59bBS3+tXvLNGI/PYmMMaNw7t5rG1Q7i6PnmvvyIdVPAf5Q/Qi/SvJf2WqtIFfdhNA/ZY5s/
pdXT+4C7epuEAk8vhGj/Tkw79JoFXmpk25CMdhjbSm5fqHl7zFji9ozW6pLbDB8eHpBYjN1NqMmp
IoTe+3Vmxyt77w/eOZLyRGzVTX01BK2TIeRluDScvNAkke++cj+BZC4ReUno9VVhL2rE9Xhcidlb
5WfK5tq9scIm772GPaAtJs39u0x6TUGnnFiPCw4eajeNB9O+gTX/8v2L9ZFRGbycRqdiUhRRMg3l
SB79Q0n701JZgLOwT2zO3nBG1oF44wnjqkQcqnzjVXf6RsdMFGPHsXeoYNVqEDETxz3t4bFblZ8E
c/coMGLCA5FtvcGHxM4Eke/idA+ZGO8EgxExX/gogfE7d0IUPRlV7qWtneTtDStLKt9HkuUAPbtG
CNStROpV+hIc3PdUGM88Os8TO5N/qtmRTVvGU798S4AUytYBKMoiKKgfebX83aykvKHya8OfQUPe
k/TtjFgoFGE08r0dhWa3zEROaY/DJ4Zv/OThZAwWHog8xBAKxY+ywmCzFhe3s1iYEXaKNL/Qsqfr
1JTzwI4DQHn6mwf9u4u4JPIeFIrrjnj9bTbxi4kG689tJuDSdv5AQknLzn4D+VjeJvg6raYtHNQw
TpjsM3HwBHjq2XE2JJeO+ECRxE10MZAvMsbsTRBmmGos1lMJL14vaERRypqRq7EseAUtKKPNypZA
Wh1GmbqSTn/bUQXsZd7mFPXjovtQagDfIGECZfCJjQcgRClBon14GOOFcxOlic+SKF5N+IZkz+fJ
bfE9U0qDX8jD2E7cY3o99o9AUuQKjQJCUiUBI0dW3w4A2AIpmWKfHjcguw7G5zQaWiVy3Ev8azNM
I00c6PT1X0099DSIo0nRpPfajWCwJCwBh13Xo0tbXpxcOZ9PUbDyMG9Ai9XADi5ehx72E9PLpUpO
9PMLLtPbKOm0N+o8QSSQuiqHZ3PCgerckY1YBD6K1QCRsbNnuMjdrP1O7OyHmu4AoBX6mrvhvXGj
wmhtoo9312EBwq0js9+uZTvzWypVf0rriYOtG2YbBvhR3FDYWk0p/A+U66aKb6b8Htg5WJqUI77o
W0KBVfchpCm5AyhqcrxVNZh6xmiCgXyNPcbVC+cHvx/U/Vn10X2u5YlS3LnLixem/ae1vn6sL0mt
bAe/V83e/r1T8I1CGcKWbw//tzWc7xcjUSfG9nRszuDc38gSO3NMPK4GiQd865wROxspfaw7D6ko
jTDhLyUIR3QuRndBVCZ1kd8v8IwY78XAmr5oNjMgbNojWxlcv9BQ4LxBxD7Ix+huUKZmblUBJx3K
/CyiQmCuayylyjQGW8AYdSYTjAfzQomtOtnRColClk9Mk6gggemdWERD6lDv06lX+v+k2LRFVOCk
oUK0rCb6ZREAUzU5gIZszvdgxvQL5ccFjN9ftN19MzpvhmfpCdg1kfp8r+Tvha+1W9lleLH78OXs
sG7BIw+cQPjrN6qg9m56FvAm9cCfhZzFhpMeHE3Gk83gbZj8U1eDt2MAlAQSsmtc/Hb929txVvDO
ssKO9ov7TMPam1UaYOnc4Uoa8S3hWFvMz1wX2h+GHapLylFhaAom+HNYtrYMaYVLCeDMR0wxtVrA
mx0A0cYaY7Nqgxk8inikwAv1eYdSTLDOlWs/Nz2icvP77TEYbU9dRK9SujfQN2lF8zRv89jFPT4m
7u/3AlwXLpvyH28nuykbG0TmPbOV7rvqDRJXgceZy80janWQaw2pf14WPTvFusrRMUxhnmiw3D8F
+9Lc1zaM+vlD63A0FA3Pu90chmupDxkE4ua3R9s4SoL/soKiXIZUkG3IZAsO84mgsAwBdCAYCYTI
LcjPHbuwfvFCsTt9ud15pDBG/coOa4AtQuIlBA1WDczjin5g+ZGwZcGT8keyXqbr/UIFW+3jlapS
2CwdsGzdf2tc2pHV4iFypDSB8sgwR6WXRj16rnWlh6TKb5V6QPL84hFThkdXgTyh291fDK8B9a7K
3dkym1kVDLhn8ddoB8PCaxF9EQp85nH4X716qrbEC66wBmZjs3dqJrrEcgblXdRqWjxDG5FONzEY
QjRcr29H2Ud9ugTxv9U/GkHBTUvDoZz5+pGlmZ5/KFDKAb5PDexO71bER0KPeN40XM87GMtyv8dL
oxYt7RLk8ruBsPfpls3YfGzp1Le0MegqIJwCGQKPpsvlFRH5Qkc6YWNldhlrW5rvch9bemgYGWJF
ElO/Fa5gdSGx35He26UtItdclokn0qD44t3mGfG0c0fdgoyB/Pgr/Bzm5vMK9RtVxHpyQc4hRswQ
0eaiMv2UiOa6gH2DO3GTar1tqqbwOi7vXwRFSUoM5rxQ3NUqdUap7ArL0e768kYU2cW0NlzkiXtO
yISz/hW7391B1uD/qlvo/XahWLu9wjft2J/wWjmqoGmarn9XKWqnbq7w3J5MvTJBE+4YfIvWtT9o
PcndpT1MxWRfbkKSn3hgGzRDqcv01iaPIp2cm6279aWd3LhiVQrAVgRm2dwahwmY/QzAn78z5px2
XORxjMLPENl36HI+P/b5kPzUfa+j73FKlf2jGKZOtO6UsWt+Xz5LdhLr3IoVAPx1yHvfVvf1xMs4
AMOFKHuLEDd1Z5uVN68Ok9iOsz3ndxOdyoOW4+g4/1PC9CxDW1eCSZtxHs0sirQcCExDM14rIxEc
0rLYj2WMvyaoBW8sOq4lxjt9TTJPnBt0dg3HJmBite9K0RUBPPyb/mq6P2UhyRkl3kFFLhTBS383
qFzsa45nliMMFbQbsrn5W3GThe/SCoX6UMR9o7tKk6wTMekx3hPcPyUs1ngdetmWa93Lts68yXo5
pxFH3XcOzceS076P2G+0u8BiMgxpATvrgBigrKDYmk9qXsmm7DWeJIND0wCVqDTIdlutHXZNPijm
PGVIhykWnK45xUX0CkQyZJH9sQysZp8Et2QOYXg0FsweYLmQSSY2Y5NoUxoMgnUherlH1LL5Fx3T
V9WWs2Pvn3ku+uK+SCD06MAGFb+0lI2HOmMBziRr5yHNGSl49Dkyvv5a3zdtgEGymBXYAsW8Thq9
ddPrtjucR0B9jcOTcw5r/gCGeCPgjPuBN2Jd8GgAVojZ0skEnBJO/344RM5Ge/SmGsZlLG0KVW41
MyDh7ARnzUeKojYqDaWA+HEOTeoGpX3g+jYsecp2Y2jRhfYVhsPkdk2m833kxEMrXVUIiZDJtmjh
w+EvNOnAc9mooBIj7jmCE0gr6lpHqFmibWu53nYHzkiU8kcRdGOvBGs7cxwnS5zSgAoP5D8ZXPYM
9YJrg0kUwkql81mAG+UyVrDTaYodE54XZczOZw3hZ+0Gyc3o6sQzj4QtuvXGlv/ruMr0hVV/2Fjc
PfqruJ1bnYg+y7amSiRSRFMOB4DfeVZuxvMI2nvicXYzKgkcFlHYKjuhEc6k2X4njo1+USunLcIX
KH3KjB9B9X/oqid7wscI8HyfI5LxjqIQJmkHRIybKsmL5iLnudSaZnkAGUTXr713g099ODMbBE50
E9yR4cjMrq6XgFRoNKk5cJCL1cv3MWOW3zvJNcdBojBGgq+hGYrLPCA6Gso3eXhX6AtgLvds0e8o
DmSqAUognLFRoA5CqaEOJ/DI6d5P01OnmLOiThQiBeZ6Zc5kncAEKg1FPqTLU4AJO/Tmz84/bmtL
FXXYryE4w3R5EZ8Cv4Yco/rirtKT6DERtKqqAaXrPesHZbADJ2zA0fJnVvc4ggF+fsJwDnG5xKpu
fiiK5sGMcIwjAX7d6YCPrf6onCEJH8sV/94rqVomZocVgWfI4KkKeqPrt5nWI62CQa8g8Nx3mUNE
zTEzaFQrWHiNJYb+SVyz3CZ5oyFwsa98D257xbTJE3JjoYfg04D0Af95tUyBrjjbo/euypMuSktu
wpjE1Q3dr2h4in2C7T1OoC2wPXdO54VHvXl3TLpvP7ppXm4axU66Vy4VmMMC9H8VfOTzEuImhAoR
U/P0WrSCVYQz6jdHuiyALXfvMaclbiMv5FBvjCn0SVgwFhWD2ZgfMMKzDqB4jFcgdQWnRAzfrCiq
pOncMe4NrdFWZI0Ma/CZlNQFlYA6pvCq0ZFkxUP3msjaIyn9pkiseYqRlkEqbcwKsDYn/ndxTsk9
IsJ0lxc1XHvdDi+BqFXc6kMAerH1iezC/aC21Y68g25G28anO7cgQHk0pvCIp2htek+QdH0FUf/U
S6HVWyYTcA5ALxx/ErGEecMVS+1oV6asRvRuUHGlUSWc1b18IjbRs0pDAFFKdAZH+JEL5yOdZESR
jUVilYk2ONOuVl8Rx+/K9SWfwfqy9GokuCrxbgcf6lJLAatTjjW6fgiqim9gC52Flph1WmrJIx+M
KSPyQ0ZsUy8Makxi2nroPtdBtMAsBPxhxO5RXGRu9aMmbmO3Mn26/JV1ruJdGvrmLTu6SY4w4F4J
s1es5YGgOHgdfg/5Ts0hlwyxLCUr9R/ZZHqb8my7zHwzoJym9dHVkI3uHpCdUwTUYvaahmUqUMJ7
OIt8S59yBdnSipo+fPcOllwWV67Wf7l2/dnYFRzIg1D3Rb0j7kbtsqIcwz1nwFxTX12weQSyei7/
mPpJcjoWLwXhOFZFqFbA9ZBEuCPPu7XSyp9kn1e+iUwIjTeL06A2ZR00ql3sMNT21aa2SPMRy8VI
H8Fkx2kt9pG3U4T1VLfjtaNjI2daukZ+xFhL86pLykZHNfnBj3oQwu1laYN0A0uXcEs0qg9uurXx
N7l84aPx8ut/B2jTKrx+rvUkVpBOp8ZsbqVawjZUm9MzrVKGrhgWV/bx9U+UZqzTFEKdJAu3vEwn
kravNn2OssQlmgt5cwkQC3rHkgchTbQbHJeWcGGSEzSe/Hjn41HpfeluEHhZMdKZ4KZNk7dLrq2U
Z9X8jllP/Uem0J1d9UGsfqSEWhfeE/l2/kyWwHUDo53SO2sfEu1uXi+yTj9E7K980WxMPCxOcFdp
sBZ9zi58wqo4WzXC/YLbUDmvMVeTHYc8L3QZFVNPkn0OniFiqxD5EJ427kjEdP1abQaLIZjml+J/
tQm2/BsVlNiaKSIlMi/buGD9uQykMlJs+icOgNSq/2EjCkTIx8KJVyzOPNbmt8rG/HsNYPS/Jv1f
8aD0tXOmUBu7YLHfz6ZnU7LcJcqgIt3DbUqJrZ/OVt+80ITjc7nA8YPuaSRTLG3hVP806KFoTo7e
wVCckK19zbak5fORrcpyiXfkNKRokgG3OSij2p1jxuq+jxQBTTG4RoOJAsrdm3t/0lXqI1DvxhnN
rwNCv8AmrW4u+Qt8ubGxWAbodTVOZmNXMwpiXP7O96OgCN7EYz8JQxJS5fWqmzUITPpd4Lz1VZIj
nIsD7ekKsFikZThZcIGB+8uXe2kg9DktcvFrH8ay9GLTHhckQyzTH8OBSZhTwLHE+SwuvXGR1STQ
E/PG12ALtKuc89Np+jWuylSV5y2gNKKnMq7LWOI78QqcBlWMnBmqhtGmI1ViSPM1L/PMS+p4AlC2
Ii4gHCIMHCJthjZOlgE2bwknbYbTd9yOuhq9ItNSYCJMRckinIiDsLZrwI+lfx+RwjYeAlTeVQTu
Osm8kYfvVRrD5In4cUZhm27N3645vdgb8bKa1OpqJ6iXtHSFty6OSf1NYqQRxgeANrtJz0frGQvC
ugEGYNsCaR3Ez7T6+wuOzAbSFqRpcPnzgjOxYxNqxe+TTnB47VM91scbzGxLviHtzVkJtSMxmeOZ
M8myyZJC455yga2XN+mn/+HDeSOM+gLt5jnnv3hNBYPKVsLkxPKzYYV+9iV9wAYJIvIZ/O6Mf7b6
+fM9DYjSdMPHk8GRQMX0SnEHVofT4QPQwu5aRQ9kuuU0huOqEEbQJh91A9TQft5kdu997d/Br9HP
sr/tBVPPgvOvfezQc2/bpCNAOWWoSuWWNrnXMxFbfIA14CENXksr+UPrxwb4uRy3W3BtrC81WfM/
tevbZyzfjsGYObl8e3ykq+S/XrBjGlSRufehlOyawLM7ShkypWYGQUBgIvtA31nGdJ4r9177ykRN
5R+r92ixET83NH8OsfG3vZWQQiFqHR7OvvSqe/hNKhb3ksa7SExXKHC4yvIOiTjw5OTr+zmem0Dt
01SSIpV5hrs/KWQK5dcUEZqGGkFElHVkfKInhJK92I6Xod2J+cXxXOqM5LFhx3uVZrRmGkt+VDLR
p5YWOUbYKUIoAuC6xZCA/hZ2HD2Z1LOEluG/viHeSfHFrJOW43a/PRdS7AOgBtaBipzuknVqqXAn
4APhYL+2gyaDd/FlRIRhCO6oFUIv7aO4DcxHHJU3QxlsVGEunXibJ91T3ivEyARI3phql+idw5MT
WbS9tYYnLhnlfWwDK8E3vbCKOR+bKW8P05LDrm1WhcydsF+q70jUsV0TL3UPX3cCa5smHPiiCjfX
muhK3l3335nktmQPR3W/4lNi/YcRhDWIUM3Jy8cPymT64GdP27mKGvIAuZcybLJ41fwjq7odXUOJ
6AWYr8kibAHFhUZLPAw8iylonYf3iWV8TnxXrQwISpyrAeXJpT83xa/0IBllIRUHYP6GOYwLBTGF
LbJMqzBXOOCV6XRgp6N8NjjPBOLhto+bI+2dlXwcaZMyPaSDgGX+LfiOa728Qob/xZzvTF0XC+kx
evrCtrLem8+rjEJHghXtx0vhpMrQacxJLysqHRpPe8uxX8OqfJpfiq36OlPvD/R7aB8OCB7JTHcs
CponkhSA4TlBw5A7W4M3bvzbL15Zl1xjGRHLD/RBxZEnqG6SJshOQQjX0OWoQF0Pv4jctXzaN9WE
FdkwQV8utSqXf5T+zypg5toilXSvTPnPkcUau5JDMi1gC9xNXscn2ClTDeIPHUbCuOX6badMe5Jx
StB470A4EKTb1RCDdksfp4TZHOXwmBC+8rOoU7ZV8wcsrfVdEr3NRvdTbk5V4HgMp7XRI4pI2PJT
Gpy2SypoT007P5rCbhmIhtU9BgCwYEnOJcjmoH/65a2WgJQObf0yPztgeq93yGsqJiZvaX/ZQSCU
WlT+6f/xBaEcxdeu+4CgoUqjx6z2Ee1fVa4h9czVs40j6fFKRGNvyXyi5VkeMLSM8/VF+cCTI8DM
8k037lsRq7Rh/m4X0ifu8TFDvYdv3LvAUAUTR5g36lqtUPJ++iECv53Uh6Z4TnZx0wol1bF219bD
GUJhPjDilUIdxSG3k1Xwe8JKHzflKyJGqhUaED7uhBUgcUc/U+y9cfv643k2w9RqnUdZzc7+FO2j
NJx4Cg27DAJEYNpef8z0m2ckqBT6pKj4SxWBfQ/anbpp0f2e4EU9/geGqefQWzg2vefo1K4CZblk
Z5FmMbNF4a6GxqpfgerdpFU3euUZHEz3cSPN1qCd0YkI3xxjaQ8Sp7GCvDuu2jEs55X45S7C1n1U
aiQ8p7vGeX8FDs/Ry5oWDRRg+rYmBKbAEmE3f475jNs3Btjq5TB/dKFI7bmTB3VtQ6DfCdnxkw5V
PIKt4umApzAh1d2/knEm2OT9DSlUV4JZdyIp+RBtbQ669bNzAM6TqbAIhihjHAhSfH2AGq7HSc6K
FBqAY6klTU9fLAHUjDcjvwTz+q14YP5ORZYxubkt+w2+yn+ugwmU1Cfn0k2I2u+Zi7+9Gq+1ZUIb
LXBVTWQ9YRDnOK3QruwVHc/v5mB20UKs5/kdkIeDDtPICJJRzjYoNWAUx7eibjpUGvTSJNk2L0Kl
4AhTtXpJU3ysVICnD3aGx7Cw88qljsZAAy5fHW3RHGKefeZeoKVLQdQK4XLrM1lAVuLA5NfoS/PR
Qvd4WWHX0xzNbIAH4LTOKwSW+3UwloNd1q4HpuKRZAxVxJk2hiVSVJ89VQRUrPYmEybetgIVJ3Pz
/elncI5mvmP7/syf5iAnnH1XywejvOH2W1U2yy4kTLGbo6ajAhM1YBa5LguviM3PaLWeOytqOPt/
SujY+W36G9oCtPdmU8538IYoDiPLdo7gsLmvoSCdM8f4iorUZjPAjdhdT01nnEK6LtbSwLv6lF4U
FaIFEyx55uI6wjkSEOozFNDlgt22SalYvSCM0mFIy5ApShTsY+87m5JFADMqDbifLXsByGn6C//D
cW9m3HHpUMq5zY+88bkRg0EG+obPKKCwXKJP66iqvpiacDmv1QYSCscfT7ZLLYz2VBj3sk7se4bs
WH+nhPHySrYkIrr6IskeWHIzO53DqEPvpCveMEVUCIwyDMpp0t5cPR4pyyUp54Z0oG17ezhpqGxb
Rbls1aUGzQoCW/WsP5bPzpJPszSKg+eN0xLrx0Ufe3YF7FT1hM8rymWY+Sv+sIu1MKYW8bLEfl3s
6EHEkb9o3ItzatpwzEXYDQLyE4PvlOBR0gKXDkwhGscGfLToMOPqsYsOrBZjRoeDJo2XLlxd5E5n
o4qen2Ikn0KfmtNqtnJyFk6hkmpVGWC4q3dqu7tWQlSVaIfNteMB4SgRv0+APIv2XlCA8Dt8VLxd
EaXuyRX5nrCteJSmr7IBgvjnJsDfwb8NgK/7a4HYiYSM7gRGuPnUedb3vHxaeRXKVQL2htZr+HzP
9tfdXMBntzEdNhg7sGL69pG5tvGTpaSqon8NYnA1EU8F27KxHKGjpIIIBNx0EquGFVU7MgSCBK5Q
pTUxuCM06Ary+3cX7clsOvzEWhAecRrsU4brturYtzjM8A7iERa6KySOy07ze7nlzr7Ie/4c0Fd+
jxf/tfZniFyiR3Qc/ZnzBWx0NTKNTxzUiYQRG4OUxD33BDGIpuLXdfHQLMnyyoegunYmDml9SHmn
hX2IgY2VcQZPyI6ap+1DXzMMlvzTson3fi1rMUhB6X2QqzwjTMOIeYXF2ygiiwwq+B1B6/CbK+u+
HRhsKeVAkWBn2l5OVFrquaNj4o7Y0WoPtsIBPpx4+IVDeFdutiUP9Kx5QrYyiqfaXNkZYzOj1tGQ
mjld42xzLqT+4QYbmx9PGeVWOkL9SDPSSdVTGdMASzha61cEoPOoiMvckO9fwihitrqz+nhNk+OB
QjI+hwTvc2Dm8kTzdH9ELOL/+mhLYvBFR+MuL+DcZkj4bGEPym+0TxxVvXnkYezx26Zrod32Amg/
UzmHAKmHUnL/BWbg3JHMzulybinoETW/cfvvuAJ/1IhZ7lampSGAGFrsUqZXpE95DutwOLFGtyv9
SytWP6o1tcV9P8R6wp1F6MC0CEGNFiuX/i+YqNxWc14SG8Yu9sR/gaZsB87+hB0II6W8c8/09vXl
QTLpb+xlIsNGlPROsBcHwNz+cCmNXHJmuQETna6LIDGmXEnyoRrhPEVGQyYs16S3J6X/jVdJ//ps
fM2ADskMSIuZJ1LXkz5prPYfqEalQxy+X+N/4FFkcBA3CT3WQgGfNIN+VP6+8sw9DsNLe7NneVyp
sT04u7ELZugCMfF3DuseQ5gWqGbtVdFjoVyohNrAFoXZ531mAqtRQrOX7hirGCRq6LPYi3QL3D8Z
j2XNpSrh9azdgTk3W5Fw6v9TiAj6zwnroDlsbS2FzHIISF+/OkxJiZZMyq0x5M77kTm6iL6SxETg
/md9lwy9PsMuNB5QTHfAM+vLaCe/BeMbVDeXJ8u1Zwm/uhJnH7EPZ/CCzADX12OLrco1IR7HCUVL
TEA2BUyhQtpU0+QfRcXozPBbDLzElBdC24MqSC/aY4uTdSPUCwLhJE3GyRf+eM8z3nzEUzfhz1en
tR2KOMzdiqDu1L6KHfJC89Y9lfDZMkTSwhbnYk0LP6b9cWX+9nwrHrwpfMkzbEUBTmgBdEAyHR43
uI0Auz9dE4J6fRtScdHNvx0rdSfstIBucu24XRaq5vxJGysXi4aEhcDshXxOa/ufY+uGiZVBCI9Q
i0YLKxdMlOY2/Xf0PHPG2OS8ec3ZWohEvZI5rVahnOfrjvMZRlAiz1m+arjWUSSrE23IGBM3zZXQ
sg1D5Akrk2amTIYWZSVjt3Q2JCe+QgJUxVnsOnjwZJn2k4mFTC/uK+L3gVI0ZE626lJSBUWzs/y4
Fa9tGsD8tWcDvrCAJkOpM0ANc2gCQ3eV0eXlaqwiS4bvzPKA7XbWb71HDp3LmSuaeBo89hfB/sIe
LLoR9NQDpLSxXQMpz4qnD0DoD3Bp2o9/lEwH+RBlzHPtVJLyNznM79KN7/SMqyZp2F4GkHNWEcR0
o08B9ZoxOtXg4glfCMkzC6hKNKCTDuxVZhNVtdoceBPI3hjHMVzP7SM7qFqFzHhgY2zwnYWrd5b5
dDhXTBqfTi2Mri70E76rE7J+DVlYYE7rKbVrMlrjIhI2zfjzayiu2YKIlESucDw4Zb27t1keY6AW
jDqpRRKQV9Yx2ktjKrqqIJTeRXMGFtdMiiLvzYSYoM3fdPgsATEv43pj2nrg3TSZitC+Gr+GaT+s
gkQfh+2w73GXHKT/eqjQTtIPaF+HF5LMVy3IvaPw8QBd0UzLK9nsiSDu0c3NoP3xlLAG3TFnnJpa
j+56w4GQtZzMC6SEE86SIZDsc5DKhaUWdCb0OaSievg11N6s6Sk3EJLBGbKg9D0DavFkCIxM5j7w
wtQuIKwiCTwCt5APHA9SIxaM8XQGxJee5mOCeRjENgwiWcJ9BD6u4Hn9jDtsMtNPEidHeJS+DAef
VF5pTIQJ9pmjbxIh329ckrcamgTaQ5HwokOrUzslHyABX6Elal0o8MmbHBWTm6idtWel4/T5PoPz
dmZP79kg9MTBZwWDZFdvVoEDSrC5qiV+kcXZ5ZOoBUiof4evcMSjwSIeMvuMcfFdIfiQSCe6vOBE
OLyZMrUq8Gb1UghDgLHjlh4jlP96j6yi16uDGarVOw4Gqonatdky20esY1Kt10AXS4dh8LZVGwhA
1JBJjTREdGneKOOi9PLEMSa+m8DLsuqPJfIJJWJQkrZ9OkXz14xcLGQJKD0K6UOU4kbA1dX3ZL7L
0MipF8E6iVMlJOxlFU3x+rJ2286Dj1VzZLkZZ1jV4l9oG07/FAqdkrwrgmoCXCSTqNvuDUVUUaU4
lx1Dn4lCX7iFSGxPkHvvRBm/dZ0TaJVL1iL812BsQ0aQL3KZvvBCoUutLh7r+Iz16GqKWSBdCfuw
WA9adsc/qGNn9QVNw+TVMKodY/R5fMRHJKAPXynAq4/awuRNVtb0y3dkayjUVSwGhXZ3w0NfJHqD
F6yQVlFmyAYNsVL/T736MKInbTTR4L8fHI06c/xjjBmw6C9BZ7Z3+dZK0HGz2QovjuYypONjtKyY
LS06NnSsRBwxdI6B5f7uX+ZBJFybInBb8iW7I1RXKethlc1hc9je8z6G+POIcpWIQmXutx/9v9zU
iecahOatFGVMaqJGeMYh9FunjUwHnRIATddmeIIMjCRz8R45yNIWRb8NGGsTp/bgOfnZb4+qzAyT
UMUyECs7h3h7hXFSoOEkoVucXJhVbjVK1ZyWq6pVw8POKUAja54nb80lncp7FVSK/4CRiimG4Xr8
IIzi+bwO/an2xK/f/aOnOv79ZquUZZf0LMzZavRCCL7t4zB0b+d7QhJW3hmbw8bJFizky94YBUGy
yRCwF7wyt/sduDST6IwpJux5vSpxJ77nqNeOuvS1mgNhSQ7mZmTycb0kjzc9SsnlF+f26BTxROPp
iXAPB3xe8gKBaFVQ6HQKuFwVEeEt2ly9YBM4MfFSLvGDgMum6aCWP9DSq3/c8e0XKBCmYDRgfyHA
Rw5+6Myq2axOZ5kABaWRfJfhcnAXMQCMZjzPkDFbZ6sZv3dvb0fj1tgZMAyZOoDpcuUEhn6C+Gx8
ub1QltRZfOU45Syt7WP9JrHvWjWGdSxZ3JtVH6qxS5GBxfle+wkSTVsSUot4vb5RFJUPMBZLyJbu
QUNi1TsmYmyo47147aN0G1I94X50yttL96CdcACw/J4A+D/pd5KvG+YeWJbYFbOhWkcLXAZNNQo0
frALOCmSbvSH+UkL2ILBJNwzADPo/ymCE6cRdHFnOgbPcwh90hvcNxcYKg2p//OxpD5VUcoh46kb
Rf36W+iH5ALqPBuqVrTbXndAX2hD24KqdF+0cPIDuS1sE9bBuqPTN5k7S+64O3+1pEOSw6fBBgM3
addDnWl34UGyqCwQuuav2/KglNU/LT+yHvV70XbXpagNOghlrJyLvclRy/J178QzfY5DDcTBWxXs
nFopI2AlzKltfkN9h1cFNhEvrMzIAZQOtU93Cz6H7HIMExyHST3t3w9nDvEa3lHL3eOcGyJecDcG
Kc82d+m/5jTJSfZcve2QIoKfxvAjDiri9tOcNW2r68dWXSih72YE0E9xrLU5R+bWxsbNU/fREsHF
ddlAfdczUqheZpEDAdbryj+6mzjZzp3OG55YSNc/rFvEY8xclyvL5BGkGza0hMNRV7qfSBznXZht
Qy4h88BxWExiI4K0tKnniDcHQ3iKKWo4bMWUDY8BxICFU9qbfD3N/zW50LlepDN1rPz79NUBCW5u
OtjmGfLO9jUP5eivfuRgtrvLP7IHC3hciIaE2GWqASSgT05BdR8cnarcA2mA1y/nLdHQ0Rr6TRx2
VfRGadkgTK+PjPUk1K/mHSlxY7DJM9RyF9q0viBwy2AokrZ7TwzwfjAFV1b0Ll+gR6pUHUijWnJQ
K4GJRshjudVz8VvjtQIhWe5RwnwQcSlm5aO0m7bY9sb9Um3ub5f/UEVubtD8zc7dWRXJEiGAskOh
F2oFlmxukv+aofuqiIIQQJ7b3CToVS/p0h7sfq1Cfc80VGRLvA4O3Nr/YwRtpFJrqUH9is7Sf6lV
LqOUeQnMc/gPZwb/4neDViYX5Z2nwAdvvSimrQTg8+b23DHQLcSg3PZUAd389AXxa9Y/PEpioRz5
Po1sdaEHdP/PakVleW409jdBfeNawdNXOb6boBseqc/YchAi0zBrQYLR00shH1nqXFEw+nOvyhb8
MmSIWdSziKCJ3AxRkIRh7ksrtccFDHmC3ZPKsR38QzHeUPtSL5xBb74JEJjTcIbzRR47AOh0otx0
LHwIauJWmSxdqNolAbXkUyQp04i+DLUqz0zCfqiH4vln7Pnrfk363++3Wz81Skyb40QlpVAnBQ3W
PUhdv8fnXEAnBh39HxGvEFcl3MtxwUPYYJ13dMQA98rnsPM5AnZCUw1+/u8lYht+DrNU2RAL+ZlQ
xU89LDMzaIwbUfFvzgWA8BDICIuo0ppCzjoFUOYYufYUDRKA6OjOt3R8yaTi4mL58uCrtHcvyXVN
Z77cpw5AeJMn3q8iBdBlSG8KLw50hqQAU2YhA0fQSq5AjLX6LsRSNTbCl5a1H4g9ZhCMD0nBYkkb
WAJL+ovObJLgmAeljVB19j/2AbcKMdDA2FQZJzkdWevT5oRseVk7cHDjGKKzFhVLwyDW8Aa/xnU1
N4/d0iDxTsNBNtJI9ByjeQ2ztnCBV5i6sSNBltN7Df/aRPHIocR4CNsjMfooIf4H3M5zXA8AgBgA
yCVosWmHOIc2swvUTwaB5ZfK4kw7jQbximpg7HRHq8pGM0bvJDQNs3g3gmYDnbiPKuLNRpDHU0Kx
WqACm6p4fann6IFG1wkkG6YkCwaPVFiz/ZLwztk+G/1da10qHtKyiliQr7WNYyzC/rbyplqLiyuR
vXkTHUm+fpDqYGOKGo+dcShwsj1sGupZ7vnL650WpO3MpfyU7Icy14RqueUCnp20ANWBnT22Pru8
nZcC/92Ex1LNqWIdHiqsuGxydJEUr9GcE87DZT58M0lf/uC9sb0T09LYdV7K6Kno77QKF+CH52O2
ipBE0+fYASwU5Tv1zbBgROTX1kjQlSgZW4pzaYijL79oEtccz4eL/yYMr+LKidu7gpu/0FUy7l0+
NHJRQndH3BnMQUsiCw9RLU4/z8r1exdxK7B/PyD+i2eGNMMa476az/v6/w5uoUffGTIXSgkovU6c
w0evjR4NiI/cU88NKmZWOZntPO4ULlZTHgiXKRE1czWSCInclijOrLRYaTf1UfP9p3tRCtiy7yT4
sApoqZLNUoiIkzUW17E7or4SnibpKtcdKXP5MTV2irXULtKzflnm54g/yE8OAuIhYbem53ktyWD3
pkS8lxqSz8ssH4qmqirLWcgA3xxhCzlf+XVeHYaMyl08dobyO2T70MLgWBNSVShc09Ec2i96OK1b
4wSlalUT8cVgQlGDkZjGVRpiIM9eiy6bFq2lKgzD4vVvvogMkrlrfOv87FiHwtY8cXKpaPJhaYMx
r8rpRZQN4JmJsuPoaLbJahX33Td5lq7Fg6VMVy1UtRTD/luEgidjhQdD6DsdwuXiJMJ/fCyYOot8
1/YSG46keGgsii1Xo1yqt7dxiRps+QWjD6GjC1uktxcIybzgmbmJ4HxVxpOWOmdo8pyOkNv0I+/M
Qk34cZOEwVBBXE9k10JTBo48ZoH8dybLwiJZ3qXt0PGyyl03GmJ2CuflSJThjRNVVr8dllYaXVdr
iN+9pD8xHnSYVibksZcOQKZIq5Oq6gxKARK024cuLQ8NZbIPEPF6UiicJuWUdNR+4UZHw1n5jWpV
86m1GJ7T4JfgKcIoXk7K7t+ppHodgBrsc26gUOedm4nKnJVZLAO8f8Dg8/tBarsxQ80sU7+G+bOH
bVkK7bs9mmwLWyV7gyv+Ji3tyy+/NS1eLcameRzt+4J5ypOgVdx8vUoNKkUpvd+YpyR7csxIqt1A
jhfk4FIJj2n5enGmhnV6c0k2lzEWlgTvTDiu1VAASsIK00pwvQAqKsF43KKoNPUbgjyaKSYu6m1k
EC9vfC2422IeUFE+jUUG80UdvYN3aKdbTe4J6/muKQtxd+7132GOJQ/7/VEXs34I9dBDhGcwvQJk
G//os7Lj/7zs4oMB2nTa/XSpl19QznkvmWFZyF7haaH/IKk3xq9PF7Ypyut0E396Ta2kKoJdXKkH
aP9UorUPMhpR+XhJHGAHmaJ4Wpr1BcYn4Kkq66CTTht2kjzvWlZjoWuCYN0b305anMfJym3XldxN
MhK9Ow8sVsDGREZPQj9z1E4nVf8wT1W2dwByLy033KjTTvZBpCMTkoPDCwPPj44z5I0/i4us1ZKw
gw/huZO8CcwUrXwtI+0BXiUdngsroOBzRPGMpYgrhhPi7O15P9Xr0mKFdngEGAkC0TdunX8ppR9G
aBM56luyAb1FCZbOvvyuo1PA5TVngA1vqJc6MkW381QZOvlH2s5BpbSnMKxFcLV3H420Tr2j5FWK
M1YRSudZCvKNI5uHWG0XRJZBA8uLDcUFfAmP6OkibBbeQxQ3GzPfdc9Vqh8IDwzHmzMHotdU2IvI
KzJcArLxfaPld7aHOL691yeeLX2xI+MI0v1E2SBjbkHvUw0jFNhdYS/skNqN0h1OSQHKqN3R3eh5
vPxTMNLHu3LexgLNZcabe4G+4HhKAe2hY3z/tRIepEbtzCFwEypWVJHn8IFpamuoAq9uNikWHJCD
O1cuP6V86TxZtcR2Zhk4Nkgt6pT7fR2O6omVTLiOPKAXDgLD3Lwme+Z7LOfZSltFvTtfxOyTp8Iz
FbX7/dz6jWAtp0LL+QHZxYS4j/IGTwBoq8QDSzMUdZwb0BA70ennB4AEvF14ogieDbNhd8iHC9WE
Ua6jsTx/KVyK1I1luFFjRQPAoCe8pUjgwjiVoJa476Jm00IH/KKdAsCI9+3obXL+mju668wJdd+L
zgHoTg7H/T+IjU556O7dLeoVqoB4KOnsj1E/4RENAcxUl/beZyounLCfqLHoVd+M0fmIau4NDtnY
7Ro0oz/o4xttoGhNtRUs/urzEK/9odegQmFqT9eXxok0axQOKhefZo3j/A4z5AwcG2nCYNGlI1eS
EggIMglig+bqjHYJuFxQz47nUGmSC3TN4hWFu9IHukPq4XbIa+0MYTIybkILRsr7lOkTlfU+xiuP
i54DSyTXJAVwbvcuF2FVD7fFZA/s8k2hjbbBgteEqNeP2mlo774zTQGmgEJBsuHVv4dh9MwYxSU1
MQN4ffVKpDBiVinQllQrSf+qQp9nvx3OobAwBHAS5bzAnhHLOGw+WppsbheRkYjTOfZJ7akJ7CuM
Oeg++h8FbDkvFBUowe17Jzmf/zkStIdVBAzryXnhdN15LKXleYGyS3w8Sth6FIAiso+6lIqeiB9r
XGYFmV+Y8uh1kCfwQU4wCXDNVoZX0b0dJAVzSuLJsigmt3ogLVLTeBFtqbyoRBqqBxqhipwzrcYO
OPnt2zrxhx0I3EmAtMs0tFiL/eO9J5NGEQyiqetlBjNVuQeC7q1H7Ofe2ugcfP6XuNxHWPyXQT1Y
tOCiLezSD1b65rm3AWFASjJhynPQS5dre7xrO/DXqCYm80UODxoh+amUsYIncMmzuy0iiOf/1Ziz
bDHNjyf6xSw5ulpp5ETTgXJmtY73yvcJMzUjgEMxfCmrwpa3X+cUqPyjcy+lfC7H2JhLbOYOA9dH
HgxwcLq7BTX/6HH/JsWrqRzA9+z3n5AbfY4Lk7f4TTPsK8WG/chMlYon0XPrw0oBNsccmRu0tZMQ
sjREP8HoSePNP5qExFo19+LgcGJ8OzG3BdVZ59twYHUvxweZHaa1HnrA/9tmGAZjoKlU9p4VpJcT
VJ2VfFyFYKUNXj5dvwQoJ1J6Wdeyn2NO0LUBQBSyhrUIvp8AwlJO7kKT7TNsN53a7MKeDeKkUr3o
bn/FfjpkLI1rzE3+ZD78sTx+Fg07EYZ4hDeWefX/Ly5dK43Hfqz7uiyYjznjbQ+tO7jJZgoX/QrS
ZPrsfLvCdShConvqTOvqImL5oUSRx8l+oN918KTdDpsAr77Sa4/2Mc6EDK2MPg1x2aC3zq0POh4p
84I0cYOYbeD3j51AsIzhSZI/LWlvV6HtfSJYk+iQqi+aN8UmgC+IT0K8Nxz2veaMsCFrJo5CdZmT
ySveDO0MqICZ8M/4rmji96QlkfMPd9BxZ1vGzlkFbLdPin72uVSKDq2huVGxu0WuHLmgUo3lEIy5
qJXkYSUi71fv36ZAH1cGEX/vs8EAglS59DR9EvO7XjbT//0U5rSmNiUHC3Y4JN0YmMOrF15Vfv+Q
n0qfBc0nXzlWT2eByhgUMqcYCt5DIxIQhSqGnl1l6c7mwpcGUTZiu2JkGJwB95yqJ6aMpWDm2Sfs
IUZrHUAmvI9x87mKCd7fQN+KFhB4cK55/qURR7MY7cpEYkRWfo/4R2EeF9Nb/qyVruGCIW6ivCKi
xn1j45WaOmFwciLdNfyaBxoN+W2no8bvP/xhA4yZOAS7zosFTN0BL+Qqp8vavWscKF7D3quMRvXl
V8VtuP+hw03RQGBdGkw46HAx6Q1kJ8V2nYF1yRQpayjtf8LIGKlG+D/YFX388rD++ngEhcB1tQJ3
V704pCOyvNGiiJy2K0Px39OajneJFnMWXQHZexMNqzwL82glw/Gm3CZiJv8BeVCPUkjmeIdTwCE+
wDJRns2gPoV3d4DatVUv4rRgwTdKY2KlZIP45imaO8rJXoRGy9WsFki4dAtLUIj4p16PbZ6tHJhn
2LXT7VXftVPYf+dDklGmyxZ29tKHq/S9BwFNkzR+iiqwk8RDaXVQEKtUL1QjeSdWapkqScxlmCy9
MsplsNSvp+tHD0ZbUgVCsaBdmZMbZMotn0Uzo+65J5mi3KtsG1zzyuUPuATDmekKfzzPmq+WPc5R
tlra8Nep6ZR8QILaIHMaSseA+gymsxePW4t1qxFEPPD3d8QZ7K70KHfsHV3OLm/UIvc8lEAPMKTb
2YC+xRbxE8gWoYQGjiKpGHXFm/x5vLnJf2cJDIeJccHHB8VYS91JWWrabtyBdow5e4bJZcwbTqpL
agGIftbPB9cQS4AvGSEMZvcFWuPpCXmJPC74rxUYQ5RyoR8JB+KufH9evPA7RSfnZrv/PlwzpB9F
7v0DVF8iwv0m/s4x5M50G6RnPbF4nQ0zjg5paAFxY/e2nzdYaPfY5idfxfYzF7fAUyF3ASu6874h
S1za1xe0HOXSBBK6TOTp9mEr5WzjAL69sgUOYuCFI3pR4F/X0vVnFfR4oqLwZB6++WSonSxuohDH
olnfwUAFm2gKumt0VcCurSMWVWGLDHDxmEYpMGxYt3TSEkRSILdZBZcQo1tj7UvY0SpczleSdAXO
d2kJVKD/AD0zV/FoxQrnMlTr2WP+Vtww01syd1hDHjLNdkYemAQsX/HyW3ooJtRGpxCQeYJoNmDL
S0CERm9Z5rLH2fPSCzqbMHa6UcWj6FK8SpNsWta6gvJGeT+EHQvhVHNkzHtmZjF+Bye6VsGKP6V9
xl2/AmFyj5/0Yt1tH6d3lslbYbjjRNtk5ZS3XG3kxQ7rX+M7vhSXG7s/goG9Fr03VY1Qql6c3OVx
tvNCmsQiOHzD7eJIbwkumAg1qRrALrCbLn8lw2/k3rvFpU6TIStdjALmUkDZH8DbW1cc4atBk1Cf
FgcaQijgWCJ51WL1W9O6pZ+X3Axe+YlZYRGaOnUY9mAnjorW+Qlie9ZDUVrBuaSuYFg0N0mLSQoJ
DuiOJHHu1wSLWhuLjlZE2boWsGcH7RCJPX/9bp/oLtsa+nMs4BP6AMsLMkuCHMlJO1rGJnCpDiAO
lK/m8goQAtF8HO2iiN0z90fJjbvwAERw3BGO40pPHLPqo22xn/LYphlFZ1HohaZkdeFZ28T9JJXO
C7zBfNPyz7g40yLqEu7NXX/JbXa7HrvYNwc1veTFbyxlsPV0ac4ATS8/92m38B7t3VyA49z9XyiZ
RTlu0w85ZQV6fg17hSLXKh/m/jikiEt0On3WsIpGneyAenRob7gMy0WOs2NOZuMqhMrZFTTyC7AC
J1yg9kRhcyI6H74spAhZLCU2XxvYcpoXEwtb34LvwfGP4P2u1LJJgUNFr1mI3CZYrTUy60duaRas
nzsXDTm7ugL7Y/O8OWOb4eMlqWs+PKSHZrkkHwz2Tps+xMtK7M9pNF/CJzKrt8FjcqsinuC20G2y
Ibt4JzXg94stIloxYGQDG5eRcAYh+HHqk3Fs2oj8qErG5MyHWY2wO9r46ccrRFN/WH9+D8olMlvu
EGxVqNzcjXQT91yh64GtU0cQZdYvAdt1K/4YkmGwQpia6d9TmV7tUMHBi8yl3OQxPgJFCugLJCt3
3SGB2DlCUu637XOopb/ynlQPk6YAu4H/8vPt+VD6LqpNRwNxiPEPqoeW6dqSZbNn2zMeioxsYp6m
nuasiABJPG+JclRpeHPg5JxYsWVTDLogFFVRBoPIPUNgot+UJAUqIWgK5XW1URMiIShrGZtSoFP6
DTrW4FxQ7RqTk28e5wPWj149rlKaj1/Qj+FrPFEOD0Dd/w9SeMjsFIdBY66VDvoPHISZ0+9DJTjh
O7U6gMJ4MwPbs7JbHeupl2AM+yAYzeWAAQdal+cC4/ugU2XKEYC1yzeZE7e7vqUryQMC0ejLZ9SY
QwYzk4AfhMKjhCqFzHGMRZmQPfXjtW+Wv0XEZkbqAqiceGooyt6cDaeZTmA4YGYAf+HS67xcMZ7o
IcvAV/yy9ecxnw9i2946a4IUmrFD1+LYe5P71GSZAKOjgum96zZ9gsRD0P5bqeu0aIGE3m2llTFU
G0viTEn2s8dn952o7XxjC4ixrBicj1gmnXWhM8mEn0Chv0uo558mL/EoT7JGpwPf4s2MAgwWCeZD
7jXhX7CDk0FccQbVySkOLLP8fdce6vw9JUKUJrwI3RsYFLmDmFqL0hxUojsNnusTXTxD+udzcmqb
6P+yjzDjcp/Wfvtm1xXeJ+koxl2+jB9fJ4PYwLYrSRqOUlAJghrubkbo69k0C60/IJlwLvRqRGUK
IHDlicgBZ6AoIbsT0J8ZCcNL3XEE1FkCzCc3apq1+RuSRye44xYCVQYnSxfFCnBWRMyaL415oQGR
bFiuG4bdBjauLaRd5be7oeu/zE8w2QAjVgwohjmuck3+3aput0jHJSJ9SRi/eCaYcF8MLfqZgQPQ
pcm9AqjTtwc5yYGzD4fxVQhks4YpyV5c/VgvWLbCtaGnV/amFv+SPwCgMeeec1vsF7c/rP34I+42
4hvtIQVFwKH+KQczgz5G+MxP842MN2wZbWbBWXSV8h/hAi+I4VVxi/qHGTRze5l04wSju7Shpsjf
5uv1w80U5vuZt8ksGiwZjThDOvF0nX7IS3Hgt63huv7pbyldasP7VqL1hi3XasHTDIsEbPG3Zepg
xoI1BJP//paEqG9XGAXDFSD+ZV5iHjRNw4hocEoHXi50TIFxaf9FEEv0ZTd8bDUJSzsev/v2EPxz
Y9H5kDTUBjHrm88I6ROS2Iep/9BK12xxcDu9j3qR+P3eg/V3S7jArCRguon/5T2OG+u4VIIUkzHC
gh9QbOzgZRf7jmVUcUbVnnTixTWwgXJTnBc2bYcI8MX6N4Sr4bVxbanSSDmVSHjFOD79NYAmMk+M
i6wLyxaa3fcq9OgWwGJCwRQDw73IKQE80aZDUms2+EIaXwEopN1AJMwhFq7vwTbex7nMPtV+yi28
pIoxKi0JUpAT/gy1iLGZyzNIYKzDggeY7IJiTwY1Cw44iKnS+wx+/XKp3UTEMn6IfNTDoFxgTAQC
tdc0mjQpztA3IDZYVbSI8X+h5S4GFR9iYtdcL3G1crARd4M26N7pjJz5GlU/A9GljaC9jPYuGHq6
+qMbaP6h14a1pJsSa8YY7QYNA4N+1U3sap1eKbobko4jezv1DNWhb+7utrvNhnqexwEBUyf7tWdu
lhktGzC8x1hToW6z4LVidFTzgzuKRWya9qxEHdu40Om0KzKqPUYBz0dyAn6GHojc/fMbvmVuJrbL
Mx+NgonVQy8JYQc+a8JgFmF8UoxSqM6LjOvyO7738xKzsSNimqJFDB3rIky4V5SRRA2qlM5OUV1R
syojQki8zuOWjjBuk+kI9aFj5PO+fl+SpWT1GldmAuzvj7ozgZL9zJoMIzPRsdzTZJwS6BBPLEbv
tqZfm8/DXpIcbZe/scfLEPL2I4BrL3DKzg396m2AHGxih62nJLq0dnaJiOdZH6s5ZN0MmZRw1oaa
pQhdLc7oCAf7OMpKvK3i8TF2fq27A5zDbYF71GPF/Kv5owjQ4JDrz4Eou4vQluAFxfi1cg5SShDd
JzBnfRsjbS2FZYr701QURusjtGrbyRlXG4DIgVv34LSLZ1BBy9xrH93Oy3gsTDT7dS3Etqvvj3oo
DMOyypUBBAArwY2Xc/Hx5on675bLDMyRsm4XGW2ecLJDjmmTq99k8Z5g9YwJ22G5jNwQhB+cbsR6
reY5Bmv6Jf+R38Ng/FCUAvsayzyUtvtKjLENsmEzCx0xZTMwmNGEOnrpzwwzfWphrSHYfNmh8fvh
YOpd49uF7/l+d2kd0iGhpeT2/Jx6+J/ZNDlVHPtABbkJ4TDgEY94YfgxmPVvxf/U5QF/sG5jfrrV
LQy41epbnaxLhtlZSQwyezSkgmLtiM/hAQM+uX1WUBpY3d+H3AmqOU+D/eKnmSZIhTl/ZDpb8nZd
tMVRHOG4TT9/1T5gbguw0hjMSmIIf2fZFL1bnh3M1i8DwWyjPPrPygIIV6ppXjJk3hSA5pi8Q1KF
rI9C7LSrIFEgPGaHQVvpQDokMjI6UrMpFA/9iebr0Q+UxMyE2M0fd7REyQSI7XpRYJASEj7CzxDV
ZXq2KrPLGy0MwX5QHMHFfT/WIx64Wo1wW6+DGM7+h14nfTuLwJElafhysv0AELQZG6c9kJZp7Fgt
QXiGnZKI2oXIGg2nHQqaZEmIKw3JfpPeIoLIFJ0reRCxRSdQHQhBNiIqxYRdJGVXrIK+4RGGGweS
7p1Xjk+BhYXRm3J5ZwpTML3MsZ+k3f6HNeJKuNnyMvlAEBh07q2VH5IhJQs6Zgr1rx/T/NVqivBJ
yX8sKXdUf9msHH/To+fW4TC+fRJSpraJW6BhXLklfIEh+x+nAv6Aw8Am0RqKwRlwVUVQer74ch2s
JQVS/BbcynlvYZLD2UhJqqOYMsmxX2fKZkF4mtPjChWwqc1NLsuL8RC+RS54Uzo/fyHR5WO+X4rw
6HLJZl/mDiL9H5LYMFgg18raNh6bcaAsV/A2/y3zfM98NHYUX/4Rc/YDoNo39uo/BmFvzAuGjxaX
DUka8cKI6lITfpClleE8rLd1c9JrZYMw9ja7r+FfJiQ23i12EF9uhJWyHODpPSj1LguTt8ojW0HE
PEOTA/yatlHPETmPK7Ghf8/6aRMXUOImVB+IHkvd2C97dFrbOxTbLnYYH6MTVUcAUsaq20q+JMKS
YSUBXnfTXPIeXpfcLqnUeCcRyCJN4lBe/2xbmjp0Avip/QpH5WoeHxqceSwnuW5/iFUa/WtLpAbU
R3bObvLSxYJuPAVsRsIlArRg9USb92X/w17Hc2x5TAW2guDUCP3Do6ck3Fd0AiMo2PO8M7sBPyT5
6Vk2k3U7mVNtGpftF8ZSvwmLOTnwplv2XljJsTq+l1U8BlYnQa8HvjZHuWyrzPyMJ/LOfjl26xFI
95cxGaKL0DXxWRItwH2cVn6W0djvsujQrOjgH5/5hSk7zdgUves4Z2Qnpqz7yEI5rVQDv8HftE3+
pyOBWhkzWUR8rYuiZQma4RfZ1tkN43/jypQeQaH75pUFyf2Hc7bKAp2HBZ+qvqKngT2zU81CEqmD
4Kl4x+83DQiF4qRUcJL+XD/l8E46gulsy07Ds75pjj/gvgTOZD6zkaSOtPgE/8TLOvnn0AJ+W+JB
6Osv+o4Na+dPivx1mBZWUplHN+1JlfW3cmGBMUpm6RTRB6nNPHxZWmaWL+lRhWX6yywdHQelCeJK
Wv60BIo/C5nuCB8fanOXx6XfGtAxk3p2l6gnzFXQha4uD/kjWAyM5+tM627HHH/zsgk7zFyHz4Uh
KJuVFvPaiUn7jVfutLPpWgfzAE9LSzegpvL4k9oRGlbuf+eNn2y0rvsQr0AEUXG63kw86rkRXgnK
op0azzWDM14lnlo8eVkeAVYznXiaqmy0Ps6FmCHgEmu1A3f4rOHIEQiyjigroZ1bm1q5pjV5rVuL
Ug2qVYqsGPtWORhehCtEcJupAtEXM288c6UH+2Ksz+PEBaVSO1poIKyZ1dUdJ+QIFBHJaB4hF6m5
jOe4bU2BJNNsZChSBPG66w+6GKZj/j5GFt7zHxtfsw21HwZdzV/JQLxGx4f2CSsAcpb/A2MK7PjK
Kj0qKBhn/TVk+Ck+ARE194/vunh4jsD35cpyisy46EY/UQB0jc4F72jwaqRb+sFOIxNYEjoixJes
B+f2eSouPnyucyMS5VDEL2+YUHaoGDAmggLG8yBdFjjyVg7qlhFOx39IuWgzOUkwHtQZL2Ka2BDt
eeCf1fk1yHpf26lUizzbXjjuPbivdRurx75FtgR6ybWJI5p7NMd5cksA2wogJmpJRkqTRu6TkMAT
cNiCY8ppPGDXcY167FsWCvJy3YNGquphLfgcw24rBEbfs106t+6dneLFuxjdRFGlJyVQMj/YXrY/
5rtwcJQBtrLnrYnCbA9fMBCURy2tWgSi8ThpMHJ0nSBGxkAlztpybRBuSr4J/xNuBd4my3dQpYEv
HYZO7emYlky1O8mZhhIwgr4n7+Z454VdIZFAezm8qCAYgwaBGKPjJZ8jNa+VjqGpEdNnkBZEbAsl
1iRbp+zCCf6PwT11zfemHYxqbWlbJQj8dasnxTKadJ4feR1ue3IbXKXA13djofvFsFiX4ptGAKvG
nsgNUeJT2zKHvzH42nkeEPyn/pMScxaV3Va+xOs7W8o5cPOhJNoIkpZoKSMUk/5zd8WpjB+Mf9G0
PKQqrkYj0fi1HhBcKEoJq0ZXz+9OZOTiPGb15WrnUT9BvtRf+3WN4rJt3Lh9sdcqSnilFWpxI7UK
2SZIhjwHqJWC2KR8LtEGq3LFFCwM/vH1nDJvoqzSQNR2LrCPDq1AyAm2/jfSl661jEUL1+Rr+itN
Y2d2bDHi630J9sedjcdTftTvQxRGAO748d51sF8SZ8Y++GxQx0QMWlSVIDxWe5ZlAoNvVFyR1EQ0
t0cPWbGyeKJyNNZ4r/B9wJYcfmuyia4zGAR/7MeH+qARG5XAOiY7HMtM4hCnSElawbhxnsfYL2/w
TYMyi7Qtqb1UePPAhs/DB5ljNwWvv3Zt3VrqVR9bYfQEHwwZZxIBZxAAowKEp3weAw4CTUmdFuV6
gj0BS11+8T9Iop5KGJA4qODxKPvVf2gP49028Qf+SxVIlhsMiZkW76JzoFNa8ORQNsud6IpGgllI
gwaxzYa70h0GrlsDhoNL34/fJkksE9eM8gxKVshzJknmZgDKNmCQECvCdU6kuLpDn7aXJJost3cI
aIF/pcw6QXRk5ZZKe+FAveCI7MOv0fKFT54kIDnU+uZUxUFGUzHA2s8ir3JGbkolkmzKqtx2vT58
PbzuzJL94qOfkWRJJ9GuqgAeQZdN6tOpN81l6uGtOpGLxrwUu9sbZstpquNQ6ZvV9XT997aTpTyc
ZW8Dc84PegZJoxx4Q3ci2oVKgNPhHAwa0oSjtNInq2HRmoFbj6paEB0cB8UCT1B8hcMb00/0zle9
ctwiKjMYc8BbBt7ZEQ87mdi81oiUU0youjLLSwi80qDrl17WLu8RLe9RK06sR4Q9DClFNq8HdszD
crlWIzZX1s7IBE0/68UAlaQhlBPMRSRAtO6kDigfA9V1QcnZAXglhcU9/d9H4G44WCNPeHedbt4R
6dIxOkaCsMLWaBEker4oY6my1jBp/3qnjAkQ/y793GkbYVVX9ukmWw474KMrfbYvBzCnUhxqsRfb
ITqXA7PwPeERBqnG2PtDNHfD0OSQ5BBaonyMhGXZI0s24Q1s3eZr/m4199+vSuMTa9Vfa9NG4/nY
cg+/5aNvi6SG7l8IdVpLA/WHP3kVzJ41v59oH69hf/K6Q/d7DgmmdG3ykroJIptPelALEO1RuRen
fwOYou7yKR2p6ka/4q+60c6bV+Gobe+tysTTCy6zejOq+/i3Nyrsp6w2vnaTa/fkBfKI9Q7L8lEg
TBsS18Jofcaw8Due1dy8Sr2IeYzQ2my5GOmuqEbrehUlVQUKYTOWhVCGT1obTuDz8rotgeXYVogQ
u0Aj+HpQSoYFZTxCd6/gkwK4ZoeRlO8OBcW6Nytamp6aL8XfESn8vHgVef6pmO2+NcOAp3p1a70D
ILqIkGk0czKgTC8nWMDZw7+Glr65+KE2rh+5UUZxM931DTGTKUfkUyAcvKh9oClqvBjVKrOVlM96
NQ4Ge/P/0252KGUZ1lIs+kLr7OEExfxKfmqmUkIh8lhmbFLKTXg1o9zRMe1c3QOCGAV7Jbaqjdld
INtihVuzJUMh8POUYn+uJCqn1gIeeeHRpTpnsluNQ/a0dy1iElDK0YLxzghWlbC8wt3VSbZ/uJKg
1wyOhuXZvzF13zapwFJN8s004lWg4eAfX8hR2VXZrXLx9U6Pvo7iGKmiLesqpIilhd5cbdDda4/e
odYCuEArgryEtmBgg2PUm1ELZPhSt3lsJ7zAW7fv0LgsTwD6DNFyJaFzB9ft/XDH1qNoV5BCRifu
7eOwZcclNR5X3Ll6CI49NDWNDaEDoOoEOlqWN9IQpiBGJXWLgzZOz5EyRIbsgqAepSqjI4Km7Q+O
6eZyH59dnbKls+0lbAwJ/jWhard8ubQDyHsu8YXChJaQTInaGBn4U16u37E+8EcyX3MBFUt/JoL5
aL1cPpiR6pdiZd1inQcEQa22D65kOojjL1tY2nd8nmFlJvCZAoPkft7C9BZKK0ztf2NE5U+mrsGu
YQ1eq5B830DkkrNCnFajldLMX2DKRJhD38FwvZkXJ1ELscmuN/jE/Z8chh9OJSLybvfRNkpXisai
vcpRiIB0y046DMCeIArvuOIs54c7xNkgZzIE8/Fg2bo9BT6tgxMnmdQwHSOdVLT/eDiVZoQj5NQd
kqzLOBF/fwk7/cigZeu7PXf7j1VCGXrBUjMRu7IGUAB6OympfgqAhy690t/BgjK6QM4yMRLf6izD
a9NDc4jBHn65XBXvHSU1OS47t4ooRb1e57lTwsvDZfG4Ej+1eE8obfN8d86d2+cRa/oM48d422sJ
DgpZh/Ysgkstgnv6oElic9MgFe8AVRUrdTe1ENpdsD8B3lksNAzKqq6vUf9Fflk+qCulV6lrA2PE
rxA80UY2WHlAT2EPtCdP+wtFQAYSKoiuj9DXRe0sPaKt9v/hPWRBrn9j2Jgpbn/qojLtyiFN519O
nLtVJ3NwhgLHE+8WS+r/G4RdswkQdaS4C+QTzCbF1AbGEmGXxK6EDOOQaNPfgucCLGwBtnqWGzbO
sK3I9npqF6bS6ltYgZGn9T4kpux8zASJ/kx2PLbK9R5PE3ZbIMH0sktPpv/CdAPJi2NrphT5Mya6
sD/76LFpBYKXwntdDr/E7tr/IzQXYG1C/+gLsC2rBRRZ1DbwjzmCWhT1mkl1UI3u0eQVwEFSgE30
NIxpjQoeep+CBAIVZORtspnTDaYyIuPhybrKci+tRurs2sKo5iy21RMV9MCfXqGfQM69Et+tPNq8
XcuEaFHlWI8XN8wpaVoFG2BEAZYISZYaadZCPA21NCAf8YOGBv1/7nulPXlGSnZsSAALvIQE/emd
NdC/D/5CO+bWdl8KsZziA6DtoLJtnUcjBkfwd/IK5i6gwNzZHgbKBv4Ok/waPYMrmzRZpG8AHmGf
XICiYtOut8AFgGhKO+uJGwyurhSF/NMU76AfjnqKP168nKguDRjDhYJFjH4e2SjZKe0IiCyJc1vZ
Xge44jfhLhsaARS3/OYi96/cDDSCWsZXN494+IrAuvqnSCCr1UKL5QXN7Vqh+Rkd98IWiHdIp7ps
uxXj0tbQdOmkPcxB15J2+ehfwW+mCXY998/fr47A7YCl5+atqr0yp9u2qf/mn8XUG6Pn0pIbzzJk
MsU+qDeKIwh2cu+FA5sC40IkBNtT8dvNCRqpX+b4UHFM3e4cxovl1XgfA1/6tTPZMzklJuTsmPWV
y3ACCmaf77gjYTqWNI1kDT7Ls9NUGQWzq4CMu3nQs/7p3f/m7EFNWz/TJjQY5JDVQUkMeXRHYe2L
l/aoPGJbqjG6N6LFkepwXAyI7K33mIEznPTYBlOi/quG2w9edqNir7LJ00UznWj53vHZxVHhptn2
xzKpQq40g22q7O03f5wwQUfET/RMC6OeAsyIWH9YFdHPwn0/ZLEzINS3nDmbi+z8FNVdzrCpxh9B
AVk8pbRVrk+jJNOF9zjWqGhOY7XzkBXWXc+PbWEWEPW6BlW9AJ8+e0Axm/E7VQDfqQWF8SE6AhFB
Dq0/CfNVcOtmnqP0In4dGPpkscFPSXDPGrxnpveJ4smU4oINyWMzQd0WoZN0MyqSQEhGaUXRWgAs
Q6lDohvvnGvRDfmHWgE0yd22Hly+m9gjCjw3EZZph2r082Cr2uMgf/5D3cDlxrxE2mUauH6xbUwW
fLZYJ0KJwXHnGvvHR23G+yEr/PFG82t3qAc4xtZHvfbVOy5mvtW+fh+lq+qxOYlQhmVh2N+OCpO5
NOJt+VCJm9dfDUK50QlDAz8QFcbJOgfptYPSwti5ojqIsaJbDwjyv62UhpokltINwUofFVxEf8H6
+Fl5Xqd4ejaiMVDjxVt5uAsS49E81/Kk+wMnqlfgBN/1dwH+R17GGPetKBGylKcZS6G1+Rqoau6L
hopzoY67/E1jJuJ2idOrR3/xx0WklS7/Vh2kYNKCOcDBSEq2SA2h7cTnf76i0DsS5rzQ/oKjPpsG
4+wyXIuyux3rrOsT6eOV95l5F9jWhlcFaYjo9G6UaHcwbhTFBg1IVBZd/qtvJRN65784kDiCHrZL
xj2QRPM/r0QlB1yl9X1JRTUhefZNkjSrQ6aUDn4M9ht5e+wU9UtrcQH2+HtQaaXAZxkgjx3wDf6j
ED9KcjiGxOvzSTotxnR/g3Wo3J7qD8NHXtjVOLHwkVNzX3N1PQ0icGPqpasxatHRDwjYmo+2+oxC
vbPBrCxxu7NeWhcPEBYLThiCtNWSOPbxZM2WSyCyRoGKmaNuO5ycLNNeIFDttm7yhnyi34jQLs8z
8UmOEo7+6tlbXkPdK0dyGtzLgBk312YYvBNu+ia57E4UlqQq3BhMRXel/op2UHiQkioybdQJ8/n8
Poz0XFUDiOnjXaw2C0Ngf0V5YHEINM0TDcZL+g656mWdzhU6KZ2bCnwdm/KQxYpK3irMXAGNLFGm
k6fmJRCVRSuvffi/ZAGPPObRB2OKJAgG6sZoYjnaD3UBF0f9782OiRurBjBUCIzwkco+nyTgwhnN
6UJmhznOsOLkP1eaeIR5MCtXEchb9W5spgE07ejGq1B80WlxCKC/oKfqHV3wZBUlnW0s5bdG0qOs
K/6kPVXyQbvyhLI5J2OsaxZwpcPl2aM/+ZptQl/n7CibZ2oZYDkkKJiueejlk0DET/6NdH3CYnlj
JJLq8VzHhDkVil+MtBqtKovlKOI/1KpYE8ncvCgqoKjM5m1r6w64eIez00q6zvlujCjqoTeZHQax
mRNA28hmU9p1/VELML46zGjQd0JSyNKQaZXInf1JNnqZritDRX2pWvFTGo97d98IgH2txEOvcl5d
tD2DXDnXhYcZm9AlI3qOXdpV1Jletpb2OgZ5F3ghdYn09Uw8iDm+MDhMVq0pBpOXsBMzYLBdqrhK
EDnT3fEoiWpJI6VyHG0eIjWd+bj/UdFKebShZadfgrMtOQmhouSMFMMDDJrMg27tQoXtv2UQZdHt
KqLJ+QNUI9zZoaPP8AUx+OYk5NPq/EWnQbhtBttHlZB4x5qTqufZyaHLP7kaWBuhdks4UDnUf425
0gDz0r5pyyi7x1EaVZ6DCH4qX9QZ3E+jicQ7hOTz7HBNQorc412Z4qPxN24KAZAGQ8RGsc5e6ngX
DQvXZldhCRwRuQPrmnnK2xjCzC/0/usea5mMD7l+3sOpLLO0OOrwr/sYdB/Yfm90+ppX0IRBnBJ6
AzkQFNFa4N/bXtzucfqQmQ6Gvx7zXPhgDatkpCN4BUFGgTo0X/A6G85TvuF03HojwZuf7/3r2BvH
/PnZrEQeCvpBFyIHgAEoaDl1yhOa0cdA42qmgozsrYJjJR8OrIR2/42sekeXgc6erpXoe+Y1yZWX
pAnbPgdYg+Yw3MKhSh27q/+85iFWZySCNWqEoTBkwrcW+AuI6+uC/ngUQnn0zsccILfD5auQQxql
WOAqhrmVttsN6GhkhmHfjXeDXzbKXbLKIKtrWq8CYa33/x7Y1ZciHuflmCu+9LO7YOMSO8h6Y+BQ
dWCrgeMhWi3+rOW43RMCH+JlrzONSQ+jequCHCVyy6DDdkW/Tznc0OWj9UCB/rlf7tv4T8vC2VpI
nQedbE/7ex17x2f8hGm7ZqXHhb/5QvgtomwRVLvfdTtwZbJPozpIZ84MPVy46s0B5g0b/Rz0H96H
hKEYpV8rfIN5UkJLQ0Gk0nXKYeucUxkqswoMbP8S3002hUqWxts8pI+eukSvJaJDRd+1U0hUsXI1
oErNd9cCkb8+BXDm3ZKQ2zYHptTxRdzCDfSc7txCx/PPvngxkBC3c+qDuxs3NjA2BENBj3hwlRrk
CY28B/y9/u1mr4ryaeyQS5Gy73otG7CBPuBqIPXBkQFUpe7y4Hza32oqzlgw5sRLj3pVE3BttPo3
sCzy2ELlDZMw+VeBSniC/dbau2m5ODZ7P3AupvarwFqeES+DrZCjApljq4HIHOjUEdgi1FT3VJl/
mJmP6pkEleGG4KS777vYVLWdcsX2UPV/gfW0lTxJfYwY0SuvE7qPS3KkjVgtGCswCR2F4Bt0OYZk
9Hilr2x5+/pMFsUyMNMdYqtKTf1JLOCJp4UnwO1zDOx5p+UyjVNiAfMOnBDbewAIU6S8GZ3n6JaF
zlgwLu0FpKOWbfKZFJAY3TxGmET946OhU+Pa8FSr+jyCtZqD4gMWA3sEt1GeyLKIeN3C6sEVYK0h
sTHTNboDYsuiVsp6P5xXjgKkuOu1hu5Tl9Mr5f651Yih0dIm68VKYxQTZfFe4iZ7+2fuFOt0OgOJ
CykL8VUIcZAl55S9SYYnZ0sbSQxbJwAjO/jE4nwpdseXqGd+amnri0Tp3bx96Ayxj18LvtPo0s0d
C2vFiBUhJ3uqYVZ7Pxn/g8JbNQGjkO1ApPvAU0PBrjJHeEreVtNAPzqseG+r/P0Z4Y8paOcYlplo
FHOs5FgtFBQqe08vEqofXpo5sL4v2NB7nq1ByP0gFCrr6KN4jUAPns+jOuBgQJS5UOxrfMWc2NKo
JilptYG4+IhgT47sCRN1j6wtmzLDcB7XlYI3tlVJ+2NdB5Gs76BaFH1sy4GcxuXlE15GJ2Cpmpon
SX8ioFUJqFdCdp/0v4fWp8budhx/Hr3HaOU/isyD0hhJuguLGMVmxySj3u1GQZak+eqSNMAuGKjJ
xObjlEG47JkPkf4SKGSVtbPJXOKM9cyfN8zGnrIIXuYKOQqaYqxb5iJAUvucuUNyI30lN/jLW5mn
sXSQ9sbmx3V9CT144ob4JcWVBDjTaMP7P+BvoX5pcU2vxye1P5gFdtzTivQMNuAg3DerUOJZb/G/
OgzDC+RmOuXwCAMnMJbIyzjvCRjv2bvxbn2FWJlHm+6W3U/jmPHSTnlCwxfFB1lTGtf/BXpT0NVk
NA2lLqJFijaQh9jlVXm3P8OP1ILBhcQkv+wHpz1U6ftz1wt2aFqhf70V1LKjtFusgaAKD5tlTIVG
3PqrKVq8Ye3bw0t6pYMPdotS9ZgsZQ7Pt681BiGt99zCPBiSeQ5x4x3Sev06XFuh3dE/MjBg5qZJ
ZAZWBaGksRX4s7WRLuRNkGBFgWGQRzrNsPI07PEK6ALLYLcoga/eVerjR+gyM4d9GAjRTlDAsyr+
fZz4TKlEG8DcKcHrI9BuzF61yOWqRGX0jm5pyse9AW3IgACPscWa8HqTyD7B+4L2oAfUrtI1VZyT
c0JwhU/ecS3v7zoIAqf51s5qdMTk2A+Fb4Bu3IDUTbMmCUBw1QbFHyqaLTi8wVkZhbhz+hnKk2Qk
9HpZ56cZFY0JiokWPCjQDhCv+6g2FBWfRsy88hCE6n13OZed1fgnXYDipf9Y3JiRD1dRCGnQakEZ
T51A4aSwOCZe5wMuhT/7MuT/bPtO05dfqeJt67KNLUcOT8QY7eRnGZX5KANyOnUlgSOGo3xQl0Ei
crG2eNJNvp/CMn6hxuRVJExiqKB5YUNL3hUhSnxynKmYtLv7aO5XOfVpuqzHDQcNQMJD9s3KabdO
1ceiiisXfdRg8QSCJe1nuNP9WUNrzFT7ySsuIz0oPBVNE1kFbSAEOq0LTS9BhXTAJw20tXqUjwrS
569yKMnCfRNumIuh4+9ggcEYDO8QPr3bdVBJPkjUKbEvitjE6wwpLoVLuOXdDKVF+YdDyWC2U4y9
FtLVW8PcX0sFSW0OwEJi0Nl8q0T6xq96bIQ5r7ocE7t8K7rM5ADV7F9fRG25xS5aofGf82B7fLi1
tFzmXpOBP6jvIwui6pcN9Yqbj3PzrATLuD6VnIGb2c7yKWwh8shjm66OEbierNlzGd/woT8RDMav
WPGk14xE2IUnx1ihQYcJsn8Oe2darE++hwvV3YIWWB75gCtv/XQuGFE3JYvGHzDXpl4BNS0YJz52
A9wwwQ4KCsX6rDLS5fRHNXeFoFItzN378zFeucOeH49SFxuIBMLUa0wy25YJSHGOngrXcua7yNF2
8uzlqYG26dKj4ZrGysCMj9D+5EdO9caHwdyFgR5gWWphaUC+E5rH9ACpnWj3RogjovtQrtOKdI6q
53KvcC9JdcIvk96aBdYSlxmLV42JZS8uAs4HVkA6RvjeMWTXKFtSnZIM2PrgqU0JOAV2lKjwrrzS
vrjahyO4v1wdHTFaXKUwYkxCyJucncB+40x2bLDgCj4aKCGYtBbWl6g48mPoE28H61GL2Dj7AwNt
Mwfo60zJ+1cuqjZNXW2sLwh6j/z8IF7jTELGz4Kw18WJSxX/vkv9eqWKs1+Dr5VcbCafnUx9h8ic
VcTLl1M0vVbO/fSwTnZ4hHw4VArekilMY7C0U8MvrlLgx0A0T1/q+4C0OrEIEP1Q/7q/ktpD43j0
FUZQlXVDBaWW4DY8Xb0Id+1rCyfeLSUbMlxgqru6AnWwJUqa4bWGxc92VR2Bh/hcSSez4pmUHt2e
MAoSVaI+dD/DgqWmknOI/BQgeqHOEPxE8OMyESV7mZunbtUYbOvn1G5cwUp7sj6RtOeR7teiEtoG
uGB9Cy7E9uBezvVSceIePn4VWL0r1p8jtaIbeC732NX1szPoOlMUIEAzIssS1oHSms4p453t8UQw
+RaqGwTk3rrmo0aVgHntDvBfTmQNAkp/TPmfq9mpkCOq2MqS38TjstyKz0khevg/J59hnJPA2nVg
q7Qi/vOzxrDu6PnVIXl9AHil3ffv5RtIb+2yGU5QiqQq96s+zXtp2SLmog9+ok7w4vy8B47dlvfD
lH6N2v2BBsIHnYksIyP38bJq/fFwzcvDebPiQfuF1R8AU3uCTklrZmlLY2wWO87kEe5PoQ7O+y6q
vy61IZUE/J3Ibxx2dJbg3SOgUEE1POAJb/B2rgIyjY8fxneZfBfmd8ZaMFm08CGbHTfpGWyhc1DK
heQ91u52+m6uLYnYWDRB7jCZnYHUrEJxVlrq3AYDyZuSr44/4xM6eVE/P8JBZYgCDvAuXOqsfI4t
m2c181mCU+NrJUjxLqRt0PmFxhNWH/GsXc4Jj/bgDJlbN7Ol4rwwUXzCBO0z/qBZupAbY/3XK3ZX
uuRBdPhe131u80moWeIDqXDvg81vE6G+99GETtRUhYmFs7FQMpE+CQy+vFAX5Kfm9PtYTx6PYScC
KCtP9h0IzmplEplI84ZobIAF2jmej/PElbgVOrivgaotcuhYLsFIKeIg5jk6ia6sdp3Xx5hUpqoa
m0pe79etRoSZpncAVsf/0UCIJKjlda4YcjIWkZqB/ZgHqs1JXqpkq6aKlXTWHHvnWBF31FqJKoE/
Ga0zOpKCUJSF0tzzQtyfBRnS3vrNBqAhVkvA8iRIrC8pdbW4/LunibUM4tgLpro70qJ6SiE0ixI3
qA4MxUib3JZeqYk+89mNKDFcQLpbkvJqWnVtV0SQHuFdH5nZhWhKZppTRWiOqpyHOwMdooQxx5tA
k6M1YpWN945RkaUNDvqj3HayQ7nr+CNeQmaSpM+FYQVgoshl/FpAsM7558uIENLgDzl/Dyq4hU14
ulkk3TMFO+NaiOTTa+Igpvqjr/Co1MOa6eXQPTzlj5kPt2qDjUGm20cW9KHeP669bHgT8N8YXBcR
dpN4CGeebtKQD2QeAqyquru1bLj6PpFpOFpN+wI+g4rDJIf8lfSVfRcJMUhHfG0oFjUNoWwYNVbJ
100T5qn/ssDhq4QS5qCK8/SJ2qx/dvFC5O64Yn3Kx9VGGZdAMf8S7qJgoYujZE6sL48vPmnpHOnb
6epaemMCO3UaJG4u21sVvv5y1i7oS2PbvJgqQOmDglm9XwLcm0+FHOz+08D/XVTvZBkLymSw28qx
pQ4KrPvS/mSgSKcharJyszN66dNmy0VpLOXCtdXR30iQkGA/IIf3kxwwyIgYFugTkKnomgcpPjoW
mB/fUFG3GvJIq7bzfZdATJENI+7SDZs7wGQGUFucmR48a6Sh8xFqdvGio15XVDbkNyscePv2199S
fTscpo3TBNjAtudf03eOstzu7xDVvzgye+Koo95maTQ+0xTYxlJ3zmOMDvllsLlq5Sm/2tpHXXGD
xOclRbJuBQS3fbKR0UUeoMf7QcQ9sJnAzBtGoK7Le4Mvu++m8mYgxLxi5hBo1RJ1Phs65jZzWLbY
8C/rlYUTkCeKgga98USMOoxHTO04uUz/6DCjR82MDDCLHWOwXLWZHx8zfLbujwgWsL6UGJw1hyFh
gjunqsSB7ZQMzGdPo6+awhQysfp0gsKnxHG3WzMrZcZo4iCG5n1cq4iluP7bFsZSCkxpAKhmydhr
1SiNTeUfiOTEScqmMLpjZc6dJWAypDJ0/PrFZhBtzSwrHvLInKmnpows1y/CZ56+x7mP4I8uEYFi
sIFTBuQnL7LNcwgitIDdiPO+53ahPmKFVANPW+3Vs077r3MEtsx52dJ88vZz8fwPQ9Wcw3EFfawJ
bfiH3bLwYcoogfSMQeiy72r2p9tfjoVk8VxwQuAPPeCTs6QzGdfRFPK/9PvvJrBLgH0uutbVb1IO
5bfOVJ7VhiQycU9z6aQKcPzXTbWbouMQFYLZI3A2I8qr7QoU4WDI8GuSCjCet2CpZXlexOjQ0UzK
VROY3Q9eVopwFyD+0aOgRmu27H88d2ctDu+NDen9Ir+/ezRJHb6EYkM37HhR0DnmFY3XdSU+rgTp
Cg4laHG5bXSHc8fMxrIcF83UNRnLmNr9gFuJzYUFf3M/BI19tCoxmkDxOnxdKEGk7G8cfLleLGFL
eJYd2cj6JnXseQ2BDz8fDEkkbf3W/FZJ+DpSK1KZjsjtSnraQbZVeA5KOHCgjXsEhLXKZnxol+DX
1/NH9GPcyS6E0V1lqCFL/S/VHq+4drhfhtya7OPL33DYoNWIHLZSQM1rc/ELnnHjMhicy+mJmK5G
anOQPip9H41esLANe3O6xNCOZwdVERZ34B0Pm4u6VQ3udZzhXFSEwzXlQlKzumPn/7tgAhyS5Nzh
g8RDrGc7p4oevR0rU6MY0OxqrbchzrrLRMtFZru/DNFfelfOaML/gfReYL/fh93kjKv5SwF0HSNn
nyE3uygx+xM1lIE8UIwdLepBcoo9lUCgfR1+BlwWOisKAswNzB8k6Hah1jlYqvGzSSAJpV/4LFGw
5/VzjZ6XmdZrqkKo7BP4SsPnte1Pnw4MzPE1vfag1yTtzN6jDNGvVNkCmdrR/4PsRED6fCv8QKfo
FVK4xMQM1hVN4v/NHPenWl17rTbHhQrLHd0ks5Mjpv5mLOajWiOm9ikfvfkB4anMSucslLxTkVl9
VveVvj9be9jnmpv2S5FAffMuafwupc2sPmKU6mYFjkkbx8VAe0KtFbevsyygJj3yBIIf47KBEfGd
yFW1j7cPLZWBrKWneeaAsLh5wPfzGBszyCN8zMWhkgZl8lbTU6cMkdVfxO+0E+7kDf3AKa4S8wE+
cIz6s9ysP5zX7e7NL0EzxVxjfI/DuOLing8BAWkAeVovyzVyxC45kIOPXEjWIFb5ZHCZJKiBK7Gk
VBDWh+N7Cf/hWjpDjtHI4pNKBeEU68WdSh4lS/6vgmvFgWiwpJQGn6rV6sw33jL74zYsPu7R8cZk
7VXC/sv8GOACjcexCJWWs4zbHZ+cDAxVx01Iw8rAs4OsMvx46BqK2cqp28PZC0XL6AE/KUO0rrBw
CDTLz6N4aKww3fdqRBvMfcxFc8kogBp7a34tvixv+s58lXmezCR7FkU4SyPnNzklB2nWxzMGHrA2
7Vhr54PXXg4mSOI7wnGi9xSwps7eiqJdrjh152LglTSMn52hlxXEW5oAXMuqavbks8njShtqk9ZH
dXZGSuPrZVNVv/MlubW3H2zpnJhM6JNbrjO9SHDNbYpH2dmeQzyRfRoifT0jQhXP9AdaDTxkorAn
RXhjpr69puUw0RQ4gCpGwC3vBiMlN9gaee4Eo0JEHlMwaTap10d2ITh2grnBIrzsvdiiJrYnC38i
MPeISthpt20+ESzQ/kp3BSFY7qu7f7G7islEAVlJfcTQzUMadHuvVAhy3sk5YhenogYN7Hx3oe2Y
IeAvEZQEpOQVMMHhiOJDSSx7saTzAyllNsxS5Jr4KKPDyAPQGhKzjRlmrY+12droi2eWTyGsjLjj
Yt7a11YiwnvE7kU/i7oy8q5xxbfn5sAQbGX4so0AX+1TfgMWlfMz4tWQpOdillJAs6KAWBlu+lPs
8W05dpLdduXLgaa7ugqItOKKbzY7P5gN3o8dhRoOZuMtcbIi4I5zyUB/Y8QR85ZYi1Obr+edcJAu
lTdA4q3vK2+RRsC6D6Q0z6Psn5KY5IhKrMyGN5IuRvW6DKtsU8u/JKjwqS7cNU8JONIejQX60lkD
yFpt1i7zIsd316EVKKwQtb86RGeDv6/63vnFX7c6GPqo6y08NiR5A/+R6CqTp60VRWG5R6LolEal
Irf1X3waMMc+w1coo3Glti1/OvuceVP5JjEnlNymemFQ8lTkb++NONnF8UwxcJQwZEUoccfQygin
eXSzSGrN4ayyAcY/bXBsM7M5h+CdbVSB34U4yTqUPbOICp29dGCE3s+Fb9L4IbnbBA7OGHu6HLTa
Fh9CC4q47c1B3lsZAKEcKv+6IIHe1xbrAKExWT5cPDINcyyPARE3wkcBaDY6a/XMCO+5Ax+B+CFB
8ahhUodTyLtoLTvTIz+vUpUuPM5HpXdIqLtwYSGLXlMvHoqauBFXjB1gMCnm7sYf55Gyty10LMK/
gtKamaqSSjTsl2icuB0wAJOOEq0m9zMeMaqozKtrw7/7dMw8t9GEiLOcjBFTDgnD3mQKScAQ1kis
Y0kyR1MrvfkDCah0SBBGMtVqM3ygokwlbJcGAg0+Qn2ZL1WUNojcM8V9Bf5P8fxtf5PCGokYbXIf
+g2l9fHeNG9ctkapNzxZHhCJCk8UddKoF5rsDAaFfrqsgnR6utmlMg87IRhN78xdUyVeDfXEPLZb
XY/qJWtKTwrI+im0cMmXvUdC/eZDuiUNxHV51wyXppVPnq8kKgQviFS+Rn6Ggy2g40iVHqJq9wUO
vyDbfgz+uwlyogaHQOv7LticxQnYGSJkx6u9OMch40IorF7BpJNmoCjImm94BTPbxQhG/9+L/BkR
Gwh2er/+QXxsfimUkA50DXcz+5eNBGsnA8aILdXEr6lXEWLUQbutJUo0Qm7N92I5WRGm5FsWam6t
JAcmz713Uso0Dncl5CZbw+GPegEmwXiUMkOJBU5sEsqm5YjapCN+TzXvf5+jj7LADEvHaqWy8pbz
fvL83CVtRWmy2L5oXkzlMMSTEB9x3kBRqXkd8xzmTjLh9PZZJgGok7juWr26jhgH8m9gzr3X638i
5F3UIW+tV0xAkXQjkaq5CMKoqMvZVaXozDKCxWzWL+ZQhyGmbqHZGy7qzUkQ2ANUdzNOW1fOXVLp
lGoQsXwW84mYVtIB+q3RTyb+KQmIy6mihm8Z/Ch8JSZ2Ebq9q/LVPsOlrx0xVcrDN5Q13p/eUjz2
G26cSoWgI5+VWJJpyJHwiwTpGJyxJ9bQvLDe027cvh4/gYEC75LQLs00ke9Xwe/cumffExjSxPH/
uldUqwzG2LI1BpDgJdozr4EXUsTCYAcUM4cMUQSTG7RaW5FuoIraie4jyPDEQjvzNOQ3rpMYv4RY
vf6lQgVe/Q2b/NjMcMbdJsDrRkkRAJPdjeoaSYZTUYOqDHRnC0dNZH65NGCA9ELZWIYdljGJu86M
3GNxnm/eHZlnpUc8Tct4/66VkcmORFqc1FIzpP6IGDGyD3fLt+sfvbHkk5BckTneLD05lOw6SZtg
tkJriZ72T6IZz/If+Rc07s9lY2uiasAp+hyDV0s3qTMUnJ6YjTNFtVUr8pbpoWvAtOkg74u/XDli
pen31sbGu6k6VP1ss3RxZ+4L3RHeZIiDyYsLcml3Wu/0ZP+fg3F5mbHy1uRjYKxsxG5ZLvpH3/nC
W4BmAurfN/3tZhmrqzcGFD/+DR2TSf4MoArqH/Db0mEmOJ0v6/szXju2fj05mlP14M/9rDGPj9kW
fSgDfvQ4eCMTIPKV8QoYX/s3BiUIvGQSgLwc1Ig7ekokoklg4on1HK0i5U4oLxgcoDFOVRXki2r9
FKxNyukA6dXqKYpObNaL0HKZJmE3KaWUycUo+YPsksPJYbnk+gGF5NnGzruoRQnuQJK2ibP5lA/H
gyuzvceRI3yo9DepCLBwVkKiRtgVYqtlG0S9O1Y1EkI7VNA8lxznASfziN+8SEYnjquzefYX2rEt
4LTfJcVGratT7rtWu993HbXj0XUaiZguT+oWiDB9OA29gnbvOm/xs/eEzoWcnYDvmq/m2QBlPUHu
SHEFplMYoNHCZfSk3mIUhDtC/gWpLIoLCTAjFNPleCZCzR1kTLnRZzc9Vx3u5Vj2HPOIYTCtJ9H6
VC49TijcRG3ADiCiCpXOkTKz57dRVj5KBoF9AAJmZN3tJ3jj1Ksoc7dxexIlu/U3UW+RD3MvGz7K
PLi28G5rSdBpby/XO1MRS2XfEIn+rmn/Xs6R1ts59Yo2si/ZfIMY8k+DGYfwgfTD1zJtrkGjrPsd
4QOSRclZKWZZMVhawFpIec5siHZ8SlSlKmo0+YGjgzCtJVakYXfIJz34cpSDQsxAnl7G3jeUyl2E
2LjKfo7SAI07wyM9HHjbs0d6iNw3cHiOxBmrllPuccJaAH7DsCYdkvgdNAq0KgCQdFRjmHfHa4+d
V+lTPTp0xJrTn3KwM8KuBK/vNhjAlYK672aERQJxTMF2lTdN2MSn/YlQ7rX1GJQ6cNVJDgFr2cXG
7dGKNV3G5TyX8Tf0TsJqOd5LdqN27smIsAuAIE9/VFEFDHot/91K8FXrVZRxqqXkeczhAsOpG2L7
Vq23eDiBnigNsN0023Cu2oE2yHN2yjpnD7XctVSNXXL7wqGJMBmIuwI2SY8LaRdZCY22rCzjNWSU
YUFtFfNZa9WU2t6ftGITz3IBEn8Jx92lUPJQoAfG1bZhg7fr9ldW3bnFXHlc+vkw1Y3iM5+13mdA
fIhkP/FbMLNaVATGqZ3huMV51Ct9tduUaFolFoUqjhnEjZOuRKUKTcJ/HQeeF2Gf1k6XLUEe3299
Kkw35Z6vBwLWuhuRMBFjYrjViFcVxwuAkNr0WjWtCTy1sLNIBi1In7J2PdomcbJCiSyOqx0DRIXc
ramHk+stFOpZ/T4unnWStdGDDFhR+ofUcKO4hrg19HS/avW3vnnN24IAwDPVYWji49ejCxFQPTfu
qCGwRnSqhLcHM01BgM2r9iH4RM+6HIufOLti98UziGP02tYDvJFINr9V1Jlep8fjbDLvYMVRzVDO
hB1fvxyVj3yvdX6GEr34fzYWtEMpCg6IRAFcIdHQl4iDZqUbDtGD+GSk9fZisEcoRNXkepC49Iqw
+nSgj1hGHxOFfhF2pYIbA+X3xOLk6hlBz2IbRLVU49Ap3aCnZJ/SxdhrdsQNhlsTNfCUUNJbZtva
cE+6Gjf0TGLzROqheasp4X/UJHoynQv9ACxQb4o2K3dfVmX5kpViNIlbMyhRIgrQUgqw87Ochksm
VNaQ7u4YoIvx/MdqBpH0Mt2Ke1wgm51IrJVW8xk3n3pnKNaXrnV0sE3d37TpVNTU+X5fejem1J8R
p2jtFGc37TDKs/VK9ZotqNURcBX8wCpNovoffD9v2NhFsqhIcJlZkMxFqK+QNUnegDzurLpz+Vxt
FfI6ylMhuB5Y6MX9tzbVYoP7+F/wVunjaDKWQmpd+v8NJ6NS9XZccOelZUuGSaNdfNcAwCI4Bmhp
5ocnU2bV5ASlpsy2wE3wJd8lA5xBn5WtOy8NjIvFSrA4AXXUYUeyG1h0LVNYaNel9TfhvHAB4VGq
OQ6GT3tc7ZiRe39tlDpFPVI4xDUU8kM8f1ChcZQC2ZhNMrq2NBFja+X0tydrDcyNUwTN8PuIaDum
dj3tJDxJNVbIwGBMXA2TQJ/5IHmrfgcCW03slM66NefXDWClBa+NIV8/P3YoU34KqHm5pQ+KM5YF
1dYVhbRDCZ/uqeERsd540tut/C1mKFObOXeD3jAd/n5UKna7/+Il/R2I1wTwpnq/UC2HlFHg24Zw
vrXrOCiqYomfOg+x1fsJv9gTN4AekiVUEmtYnGss7oxAzHXBYrIdqlizI34kePtNaSozOViubrGW
jwr9aHcLylkyVce2L9ogTAWDIHcO9AJj/KcvnA0Y8QjfH2InX12xfbnWmkVhsg/k76jpSqexmMQi
urdFLFlblLEY9FpJ0VDxP0OFDsdpKiKBN0hn+eSCzNw5CAi+t4/I1cNe7SYv1YMjn6HSeQyCyJKt
sgAM6kDh/WpTkYlcL2t/+qDs851ap3n3mg+VBIC34cywPEeqxUqWAwuO0nXxCF+3c8Ujv/A/s128
Vqn8DPJX5A8/tf7GnSAvtDW2M1LchF3wR1e/TTJ5cdbMk/tuhhUkpUdN2QJaJx07h6hAmEwDd4ZH
OyZXtZOt7qFmSUvWIkLGcTmdaUe/Z5M/Vexf9GaaF3VzFK7SYJvuotWrJ/F/zl10FAHsEaGKcJu8
4A7qOpbVJh4GV52sSFBosCf93k87V5o3L19oLzZH7NuRCzrG6THJQVi449HiF9qduXfs/7uhri3o
+37R+Da5ifVDMnVn2wlPbu3s+QozTTSWJ3BvkTtip15hKc4cT8sU44uxM+GxeY/IDtYSAmHaApEg
F789ffisiYEzL3U06BAgM2R/cPxloGTce/35BOa6ei5AVxKNUOYC6kdUve0ZKBwPR7HNpse21EjE
aKrEQnxXETeKa1sK+uneozjie1V563fb4aLSjh/+rBXdhbOSnxUAUwTiWdPz0e0KwlFDsJ5iyiLH
fAnEEEXTS9ZdXpGYuwtkPlCLOzdy57EUnoUPZxJAgimqvHJJDczHWdaQZ2EIgasS86vaTfJQA2/l
uXl0qBsi/zRuf25EjYzmyNaY5H2Yc1GFy3k7BUvLtfb0k4XyqdN3lvop0JONYI/ZvrkY7VwrdxdJ
LcpbmH2YOt9zuVB+zMIZow66+E3qSj3N0y2j6wy2q/vow/5ok3aZGbK6H/WmWBUwgTAAGO9vkSeL
izJubgY82bd+lX9A+1149/FhpwciZwOmqTYNJQXXA3/zw/VZU9whS3sCeYW4/ya8x7y4HPxDA5fT
0+d2/LKZu0O5v1WPc8Q/9Z1Ge8MEJYkIn0FT2DPUSbail9cW2rcAxcLCVyGhWag//FU8FPcSHiXx
9emXd744mBnm+62+7VjLkSUhfktjDbn+DzpX8yGCJss19OvNovHcNUrGtqXjC9UmhSVaA0qjLFqC
utVrIQwjhyTVVps3u1/Lano1/VQ34WNJHrttWIMxG8cKd+hjJZ4rfaHLzHR/cmYIC3LRQCDdG/oH
tZLOcq4iNF0/FU9mZPzxYnTg7SltYwTHE53u1Nfu/oq5gbTq5QyBy+fT72TJ+0zILMugDHNigZKI
8YXC3mE7EzbI9WdUVSCUt6jHE+iIJV+cDu4bsnDvybguZbs+lx7VTCwazDXQIQylhtcJ/KxgRVmP
4cQooZLSQysKtbsffnedfOGEvoAogiUibfha6mx1BeqVD6KmaXVUVB+TRyl7ic+US26dXzsdJIE8
S1OJZ6hhnwTOzM/zMXxqIxg6g2bNc86CKnT27iOQ3XAwb0eN7crfdOkYqZcuspsSoq+kDXanNjcn
8uEspShUVB0tX0j313Z4C0IEtp+yXN/nX4VumdmUCheqsbZ07c+BCLv1ISzJAGWRIoSToXYxy7ch
FQm+2N0Cvir9qJJo37xI6ZpSs9oyFbvWg4QEf6vqh1M4Fl8PyU2BM3NX1yuryjslVYBpiATiT0RF
mXAtKKkvDqKsdy/M+WtbYDqT7ew50MKq3onLlA/xRTQQW4nqV7YTSBNPFBMEOA/Y7IYW7//GXLaw
jnjv0YltyeY7BFHHINoPoyCCDzJvtvJNIcLbhjgeLgwB8DIAyQU47uivCqmUUifxdlnUejwJmKGr
yqb7J09AiOGwP8hZ01+wNh8QC5hSYo3Tu+a4NzzPswOm0Z3LtSnYhD+/5nb16JJ3aa0uEPITD5QF
0ia6jqIo/1CpNVnrFxIyuLx3u4lJ9uB3G7EvvAyJz2GeZdIK8oI8q1M11pGM97mhAzgUJsgZ3nJe
1iSqXMd44cZ0FCbkKsrPCPw/eQLVYXNciEm+BYHAujOittdd0WXtXuLpS7IXvACTEAdpzza7O4Q/
IidlSXgK23+jrh48n3rJ7MvpDPgxH9nw1UKRWx5BH0Pxl2e57LLr61zGCwCYMdc+h//WW0XXFhNp
ffd7X5HM4g69TdIPJJMGdGpwyOVNsZTC0n/tMMO9y/x6XcyZUKbITVmRUTwr8OMepossbSpKvAe3
al+a2rU7y0I8xfMApzBG39pGJmuEHt3dCI6oL5mYoNc9DZyMoMP6/7hyM3TaoNpOTBZ5I9VQuAD2
QJMs/oB9/Vaeg8ZjcOu+MUJCD6pOyO6IUeC3R9h7Xk/VGJ6ZmOSo8ma27u6yXh+OgzgLpjH54ATZ
+PjtY4+BzGYyyvmDbyteH85oHrtZlN7ELT7N6icQ9hcHP3AQU7Ea9OAqWVoUoJkIgKG23FHVL2TD
KF0q3x1kyGFCjBgJbRQFZ91KGS2bBNVFojscwUsmRzgax9hLsNEHFmplLYeWKbr73bQshXOP10Nl
uFysTZfStv8O1SlX4HXIZRXGeuqNf23gmHSIsBNicjVlAfoSZ0aYEEcaWCxkhI+vwGx9A6amkFVf
xlQ2Z9NvAtXPALdLw256y6pMORO0Na7smbBl7KTL39+CoxB5GjxNoxw1/Ju6O6evu1ANSBawqTGG
CADMXzgSGGjoyJfnNf5NX0klVPJbEycCkIftXcJsNydqLokXhfpssJLTjLL5vQv49lsIs0ZjaVU8
aA0lixmGJYHpkKHnbEy7kvJ9ZwYNomZU4RXos7xWMAMLwwAQL8yfKPHyODFCuO8H34dNIAH3WHO2
Q78iRG1xc2xQEQK1GeshcFOqSET2cLYqPWlnBdxSTqYTfeBtmjIPBhZlVpuBpTA93Mjvvtv5MVK0
IH72MriTaK/bFe8+vAs/bWn0NvZcO5lhGWj5eYdvG+DfW7F/Esk5PDp8ciSYq2iHzn/wFMArUDcT
ZyIxq8hErY1f8AgYO+Zv14oOFoVuMfE9rKuCvAEsnuDAwopH9S5RtDAXfc0DsaaECgdCKZ9fRYEB
Ht8hCSQF1y7nzjvdeLFOTO+2s3MqIm1ye1m/JIUOQRuWEExVFV9Uq8PWwgav68NJiLNybBvQBc2A
Y//3M7evRrMPTz9IQislsFbyinFEYUt2J6hQJVoCXUGdnzP70uY4VR3VrjRhcCcGDOOEZOmra1rn
MrrrelD4A9kdDO7gNrrqywt4GF8h5KBC+vRvWOkvmw6nEe1ykFtf6g25GGWYlSB+b3sg5GnYZtUH
WCEIpGoIM8Y+u5ZR4waZ9gxeWratRZSSMTxPWyN2LxcyIURwrgKql0u5Edd4p266XZGmSqSCW5JP
fTu0gLwfdK2TYxLbu1PJvc5+AueDzqrez45mKxssFSgqANZz+HJFl3h2XPT0mPXxFZkQIkMGcdrC
2swdfVHPheoKLqmG66JMREQizsca55U2XKsx9iVinetmYwChHMswQmqTb7zoTwAEehOoqM1ZVaim
9/GLIE2V76xjGIUsy+i/jWRb3F7c58J4emK7U23hzZotxqJHYx94g4JoolFfS28CGRPjuPUvnoF2
qDxKPxgU/TEdIhZGLiHzwifY9kODCci4BMy6xcJ5fWAqw+TvnU/rSAZqgFBE+jn/l+tfVnLtpl4A
9N50KY35ZvXBtVqhQwchjhXFR5OtQNdAnTfVTsmY5IHDjyPJFx5CW0i6btR369dHX6DWvP5R4fg6
FNPUA9G6Bvap4+IKZKfSxgU1Et/dob0nGKcv2uRtSVnMpOymwd4MTFmSPKnj5mYHM+qdB+dtSzyM
a0BRGh/8h7/HBch8h8izvazDNIuXGfgUepmELFdWbOR1+rp2NCLt/K2jkfFB8jS/t/BNjAo+Ou1V
QkQ8C2T8rHai8CkDICG1heDf56WG/D1OilsvuH57JkV+t5MQsMbWodvZCP37mm2XdhYCyRCaTVv4
TkKR122bua7/E13dB4QBGANHy0HpB6BBhwubPwhYWrSn4Skc4k41f0fPN7vHNq7Zyx3Qlc+YZq/N
KLptUbrhug/M6MayNBDLph582MfDkUQ2yrFDciITnEYAZraIxR5IV4tE1BU6KewRiZmwI77hmPK4
QZZRJmaMX7FHn9WF6uH+GhZB0tp8EUzRxp4y4C4l0tAV1sH6p/RIya90QZn4mu7X0igpEnO4oJ5E
tqRFguIXD5PeyWjKfX+OzMysY04H5Oc25M605FFeFrMoiwlHIhzNnAOUZsS8x7+DeVyIucP+0Zb5
waMh8TyojD34L0yHAcmErFW57jlD16D/CA9FdZTPfVe39TR6bSlL4GRl/gmKPOpJZujahfICVBYR
ThovRROqMrruUsb74UPen9Tkr9EgCtUxggFKuOsEvpXaBaOrKNZWBlPC89fCoJSUEK2WGgUStdn9
gbrPgw9hdnRh/IuJBRzzm38iXtkMkAdrnSEv4SZf79xxPXTpgxtLeAgUu6EK7XubnUfV3WhIIxml
PKVFPL2XPptNn1iWTx8ryXv628qwsOAFUwvxUTQVFaweK4laQBum+Wm7d4jgWwvfgKgLPsPtzvz6
t5+22igu8ViYDGRYXh/PjR6PotVoMz5R5V/6Czrjg7253XODL0GhEo/mcI9ubXATrse2xBWHI4AZ
280cgR/9oUV3g5AqwjPC8w0nDUolT1WIxvbnpzilH2UVgqcqNxR5QTHk/VEy8Z7/JsCaYQtvPlYQ
hyiPNs6IKuZQHGFcUN2bPQRExYM4KD1RxxqA8RBJMhTeMpUk0IsZC09zg0Vq/jFwriuoY/PLFnIV
4CGhjWox7ZB13/iKbgzErwZu7s6gr1FIlndy3VY+A05nq/eAShcjn3NoenJLV2Zp3jSf2a9ohQTL
Xn9+rPVXx7n3P46wP2A15oGzjerh+R5h0j/hYuaKfO9JdNbLhhuScBo2Gqf0L4JCiIucd/XXT5Aa
zQK2qN/YRLbZdWD82UEo5MpTD/fjvW2ki91wJYV7Nn2LgNbtKEiXrgVPOIbjIgAYX9jXDqKA+Bfw
UKpcG5guXlXzMr4/CZ47TehZJSLOavyf8ffCOs/GXZGm6ROR5nPfFYAV76BJI+OSO5on5U1weFYh
Zb4jSNppeE8+rF1dYr9IdhiLBo5XxyrYDlVNH779ked+lNc+rIOBj470GQLtY5zV9tXVaKTbeEUI
GxsFyhnEVnt2oY/jyL4PRTYBzvzwUqQAapHRqDCTKMqdNzGVe/aS8zwLh5b0kQKv3IOD/hK52AKT
7f8qql/5kRQTS1hajZhDxns24rZev77IENB3aDGhXHNsnKhcX6MyB5x/5yDjGiWSpO0j6MCpdTSQ
TuIpAjDO3aRGZxgb7x02DkhykkltBAU8JuNc4g5JNocJX8sHnOzY7CKvipgJjVfbFlPM2l31Md0M
2R2BHVq6WDCHpxkoyjZBDr7MFd+9L7c9gQ9b95lvLmow2M3I+QxTbAlMLkPOxtLlwjZBBihR50KQ
WTKKXrbw4Qrw62+htE2bW5PINrjagO9CINygwu/Rvgv1jsT/3LEqi83B/L8Z0+g4oQL2s44MbZu3
igOVKiC7jM2Z2NeeK+7fM4aFxQ44+Q1EbYrF7B67dkoK4at1ts/ddiFwRJnisOMvyn/1nIjyuYh9
rnraB6rMAhPNm0C48ko7/lFEfAjwj8864YZ7mZAkhLcj8z2y8XPzNNxdAYo+SCmSPsRcx76GGJ6M
XP+2KgTH0/RuYd4NH4ngUWR9R6NVY/yu0ViL+5q2OPWn4iizd1GQC1M6ukbTQAfxhjJ5BAPXMWxW
MknhylcGT4tUaPmnf/hy/hovFlMZEFb3g5PzEcewJ+yA/xVjnBxhNXx5DZ9sDZ4Gx5Xn4HFQmBpK
9BxX1bYCyxNoj8J0beg3YFDVeKitu3q6oFzHpgKjm7upxygELW1wCOop/rBKMnEfsUvtLUso7W0Z
LnUe9irQ63amP2bzcoKlZis/hksIY7yHsMUsdOHattKWU3HLvNK0jo0azCKuAPcG7wt7gGPc4qEi
j23rob2hEDishznU1EiA1UFE0yXMZTVbXte/id8wqgigf3krDmIOjCxRYp90QUqrmc3pwra6De/U
AylFI7GJkaqGzJeyi6ppWPtKT2/T8FcdxrY1oqRuU+tqcJ6kcP5KG3/opn9aCn/SzEGPhSWQY8Mp
yTx7zHAcEnTulI0vp0nTJoJA5D7rK0jCoaDVKV1TqnV1Fy6fTSHs8ESYDU9P1RondjvXg4c318ng
602bvi7N++gWEHH528YHhcGe6rXNpLirwHogLLZih3AHPGZ0uUsiuzzzRupRv48g93vQUqzFV+h2
ZKT3zoaQyOIg10BxU2UZaYsYiwpMbcUC0YMsTvJ2pQ+OPYjGnuThbYKSzJHXUacpjYBXpzBhn+8+
T7jwkNS64Hw/yMm4CmsWLP2DKFKi5mKRz2xMFExLHLqLX+nxG3WoWlk+l7fXTDiQFdx+FURWDZv8
ezefu9NTOGfqYNvK9zUlRYjCmdS5VTkvMBfPdQrJVttwptwDKGx0uQWqL07CaA6GwQ5jFhfLjKHL
8T4JOgFPJxAiIfI97rO3B0Q2d9RnUlU/VTv96zQXIel9BnGLBoIIKjBWL/KguJLrL4te8ibXZcmT
fkFd+H7Yy4QikMq0PyDWayCsJ+SpATU2fDIcOsAqrqzqe4arx/uIGnRD6PfhL/J8UbBNfWFeYfP/
WMTQiFN/LNYY4uPtHdIfe5k/WBwc7VOujz3Jtb+nvdGrGjS2e3dWDL++tbLel9eXHX5DEyLJ5EYM
wYFhhlMaw1cHmQ8iIMoKM1gzbIQD5voS2TLLjp+40Tw2OL+Yr9Ivi+9xZBW9Lt1ZJgrUqS0h77bH
Bye6Ut040krmzTiPajrLu/OHbU1dv5dtusuWwZY6B+M+n4FNkEzbcy+ViC40745TSr4mhGBD4jXs
qQjxtHTo0IEDb+ERihhibXwPdxULK2mUGmOk8oACcka1VddbXL/aXG5Mccsf6+GgBQPCqUfGjdKn
LSOsndYf+r06TtqT7uRMUmJWk7Ky/b7zhbxiXjv88qtno+mxtHlo7zImWkH52llxxKG2I9o0OwBG
gdEC9hqqYlUsNlpMNRU4FVKVRucg2Hu7b/4ckx64FQm1/EJRJwhcujTYf/FYbESnTOoh0IXZUmMc
qyGT/7j8cu0xX1CyM2r0XQFiFX29n0ZUhIeKIgg6C7CsJFva278gPfj+Uwkt3tU6Fi6ZcUp4vEZY
AFQ+sSpLWC+xLOvBvlGetC8/2vmriMEOZXjWwqDthPj5HilypFfbqq7UjZHdEtWapPi1vAdZUfSS
M9T6ZSisekguouBpDH/y1UZ8GEZ1izG+PCrszQnXHT/i2S98y4IIMXOzl3z2djXcj1e3zhsbmOAU
wLzSacbQZ1S/GJw1P6/z1EynHngiupN7m2QWySSeIWdy10Azm3UVOMgQfqUhVcjRQAxC6HG9hikM
zEW5p0mFVHL5w2Btu5YVwEiHkGyVA7/WtuY24oF3nfS7Ye6ZM+aYE1U9bg3p147vCBoZ6cIDgYIz
e2ZI4LwFcZ5noOkeJ3ZSYadV8y90FgZ4D2JAr9y6sFChLXjpoxOovOtEXP2xilRLlfGCkcCLNgX2
AAVGXdHewocGQE0iUq0E6TN+ta8gN5qYG+fg8isWmWLBq+1PEUbxkhk8aXtL6bAQY88XzIODKd/B
85ub58dg1d9fwOXth43N7xxCqw+fxawbuUfHRDJFXRa1VRS4FJ+3FfpD3Md3LMxw2mf3N2tbQbpV
Ss3GOp2apPljCoRzTZXAMIRtGTWLNQq59K2ost2P9XfR6SMjQS+WuLcJLm3f+MBXy2XNpdmg/EJ3
Od8Mg8d7mQ5WzC/EN7pNG6pxqoflOIuG7x27BdeOBkaxNX7bz+nTvPg2V96w20ggvsc40oZO6oYz
KVTVLIFyRUKz+xZJKAKRKhnYGI2dT1w6bhQeeHs7o5Kc2f6awXICaP3kiqCSy1xJj1DrMILlGZrU
sd1iOTRudmlqgEPQgB+Pvm3BvAsBCVp/me2x3TpWcXQ3y3DhFPJAwa15YoPvLNbLtqxMBqXoP188
F7qbDxuAKsx4NJCspWAS0fFnDFmeVAWdIaQbAJzy59aG8yWfkxP/9amP62/arZcenol1VIyhz0Pb
uZspi/vZNDBQnwOk/6uQzE7QynwSSFJ57NM0bzjnJeuWZzZGUfF1sR6XtwW2kKiccYRZ1CKkozbN
sGM81tFOvQMtTPMTQSz8pzAedMEB0nwtAf0O1uWV+oJx3XfXVgFPXxfb/B5tC2iyznhoD1dsVd5L
eo3KJK/mY+NiSCivrkauNJzi2RQDf4Z5M7c/7elELv8c8xX8tHLODg8UCN/bgpoYDL4EzU0d25Fx
tkHi57NNhcbTT1Qa6k0x4kDE+HVAYno2DzEzfVw6IX7xmvKNMP/2Ly/mQdfSJg4frUZ9EWbddqAY
0FVfrjWAZa/A73Hz6tVDStpOvoJ/sA/jrlnUtb3XCQN8NGepc66pPblHQWXOR0YL7ANYc4bjmxXI
/gcxqvp2YL9IXMVgG03+umdMSUiVmK/N83QRDKDmM0v+9FMzjAt43yD/zBvqjHiA1cfi3ePvPi96
CRSX26ksx1OO95ACcRZsr3K567E36Wct84tATsHxklrOfb8kEE7Rw4RvmeqYQwfUro4ItVgyjCwz
pxxhUAByeXbCJDXzS7ew/XXKj4jbTJoiqRr0d9hUVgRq7VmiCkHrZM4+9u6dhBeLoYJbfKOSAsV7
9KmDE9gvRWNjzNsQuvQUe/nZSAvV2mXddgV2v2QYyJql+p9y4YQztUle8PbYtX9oHyrcTxOTN5aA
Gz8wFlDsLmf9rxO3UoBwh+4m8o2T4/II7z+axTGYz1CdFNq5XiBIDd9OZMNaF7FjPO+ciFrf23hy
ZLwhVvobJjWFKpETEacZd0qFa8XZVfIFkHotTsUp9pYtCyIdJNyhl97i2nEaIkqBYEPJ2cIIoVWF
BcmCWqu8qJWc4Yv89Z8j2y5AlaDJcR03/bQj9XIXOljKI1TLchRe5pCPUbwWD21xMukrbC2ZlYxc
5xHGBb11q205usbrO+KP0E7rbz/njmXYg6IxIL1mNzbzcDgOMr/S5zjiDfWsfSX0Rlk7kNynydOt
t2lyMb9wmsW3P3Eqsm/zVMZHcagNXs5WLkFaAdPRrRkgexSvuvMylGS7/PCCVHWItfkQxmdTJFO8
wPREu63N0c63l/BMzCSz1q2Z71zzHbBcCPzLdTFikLTOL76qyFGXBnTapNDAgzftzORC4dESiNz9
NBxOo2jhHJS7OGV1jMFj6EJnth1tK4UYPT0oMFXzu/+/km3FXuTQWDXAREwcizH7YkDmslz3Qk1i
2dYBNV08Y6DPemFhok70l849q+1Wpao/Malu9p+CSipF9BbpbyQLTsnOVolMr47KfxDxS7hAQqeF
i+Tdg+DJqjUEeUo2kPHN9vphFohHUhH+8OV7robAOz3BNaV8vC9hrQ6Wf15FCrUt2NAgEQa44Ks2
FLq7r3UEUSOd7+x9gOWML5INMLXEhsG5JCJopJZfFM3GT04Es3vj8l3VDH1FKSlfWwKQQoULVir+
wv5mI8Thn+1rSkifHH8iluLdBV0wwtqOMv/o25F9oLv5qCe5YbaABxaTf0TSbEjgxI//7EkZuQX/
fpbHnuN9YXWAfeVQQD1IO5NBkR1HmmIwGTA7q7YYhzXCWxYkl7V/jEJUchuZHMoMkcIe+kilpBOu
/mpByhHYFJsWFNFrFQ18CsEeNa7dTE59ov4sBnMxm30/OTgnfFWsaxrrPjMRWsX0tiShGu8lR66w
GToWC3CwpikHOuZBNaZIFBSYkjjvskg2/T5tjS5FTe36x5HrGiAQmAXxuXURC9qX5KAIVoibQs9v
g3Il580mD3x1Juyf1MDVEUmUwnxhEN9II050wHXxe/tz6NTjxGZgqk+n/UrdjrbGiWKL3/HclnRK
38Z1PyoXxg8lN4RZGIaIbGsd/MjXOtmxI47HbPnGlEAbfFyS3gnsb76lgstmMl8HlWdZbCjYjmvp
VUYh02d+JK7hp4vxiY0MGPXnAxBsgfvo+az5K/Gcy3vexhwCP/mZd8xK9nVO6EeiZudxDock6L4+
7PKWDzSxwKcS6P3MNEvUaQGfTQS+uvfw84DbvqJXaCaeP/q7e/eaiDwe7CxQvlfIatGhEZoVjoo6
wtaJAKEOiPGEUs+CMKrsqQ3WIo7PDd2fvK1AtwSZL7nssbYv4y77rcqhijLIw22QYK7pIEnEn+HP
eN3pYih28ULsc6Z/BbxiFeRXI+mtIP38BXOK0bcfHuDLqy2HF4P5LIRoGvx5tbhR+UEXBeQ0hCzS
dJbxOnOMSi+KE2mWU8q7vxWfg7VX5VlP43lf1EMeWB29A5N5cHPlWwA00i1HkPQDCtLI8YIalAMO
WvA3RAJYvQEsz2uDYAtoLqGzqPrfxReJk3oo2OAsXdzvpoYtwwxxBPlbddoWK06M6lk3WcGlz+Oj
P8Zl6QEYcxmqrKHkQbJPNLJ/rq1/3ev0QS0qNKz4iIn7fDrK+JWEKCBVrENr0xEher0YFR2vCMiY
NE64OhwNet6XzYESZDwDiwPFPaZOBTSX8IZKT4LWNt/BtkEk05Z1eLMdJzWtcFpaIP+B3aJiUp4U
0Iu1ZhlaSIi/BUe5mCby5Mk8FnvAq4ZroYhgoZgi2cqRtCEZxy7ymftHSfLsEez/oewHltktFYLf
iLiEQ2NXZcdvNdn36e80vnz+snLHsj82kBg5GVPx/cjpFSDO4NES0cWVvBb609VKfDHZhApy6Lwa
GXvfgljM54u+ooXbNjZd9CruFLvgKteh1prW0RkYQ3n8jCeXjnO+A66Ov72H3l4hexb48Zj60b0L
OPzQGRB2joGQBV2T4mo235s/vXg7xcnBeA2dPW4vhYWhtvkLawqqNpZz8Nd/YPcxaDORTQu6jetQ
SPE8aXeaNL1fdg3vU404nmzdz07jjeeAS8GyZhjKRrZq3wnp8SHiV4lyg/nPKsFRFRRVyaXpPL/L
fy5Dhyi+UxvoyDUq0dN0Py4P1IJXZd5uPS+TkejbpIJ2xbqxjmE7Nl4BW2OvalCsf4UGKaTyap4R
l4s3PFENdw7jZBwGPsFPBM5ZV9XAOQukNWpVzbmoHqauVG15Ce70PwM5yFuSZOrMwI/uSWDvHgo1
kS+dXc3YWwrp/pJxXMSxyfFllGr+01LxtpIAsL5pms1gfj9+6NQnHxPUutOkGvwtzc2oNt+aCLv1
kram9Q76BFbJdQHs9LeAAiNhexcLlw4N0zXBjG4AeH0zffOXw+lzsNx9zYEFkG63ZFs2W5LACOI1
Fg0GoJdGnDQD6wov7E9BGxjBkKO81gXxJrqss9MB0lSlE40a+87c25CaoP+j01S2OMyepivL2782
6dE89D1DwcrooyIn+MMbsZ9K8Z0WUJ6pa8GhLgJd+wYTdQTVSyw0uE/btFQnK3rZm6wNY8M+S4a7
DZoV/lL8JEFHQpNhSYzt24kDyC09zKuue1yyJYEaIbx8YB+MBjT8lzVkCkQy/MtBbmeMC/83T4Zd
2pETuPgvIRCjSoZuPPaWbPPwVKgrBWWiJ7DhkQc51GWW850h0YrrODbEYZPDi90xVr9UboNCRY1d
cXNuJF/BwOBDrle4cMY6IXV1DeTJ3FNoVdEKbnaDsWUYc9lwmWt6XnKkMDEMxp9PpFED+73oK+NC
Uw/I1SclkyylNKh9iwfKkluVAGVxvG0ZMGClmVWfaMV3qKWosm9+auhGO71iAV0EjG5hJ/Ovw9XY
szTd7pT2iAXecwg4OUvqPrG7ecJjbnoYe5tI9BN0IZ/R0mbrX8Y3+gkTm6hxA3fMMSbO3sE7A8FE
yf7ix/8B35iuJUV5+iYu5fOHAQSeHJBrQkXCp387kQ1cmHka6qSnVSdhuClpugdvnbmrwgIqMmbE
0x1xr2EX+mA6ZBC9vsfFa4cNt0irztkgowCEhSu2vtDjK3OZdtHVzA0pjg1sYni/WrbhemxVZzPS
Koe3v2tmyi8W8sBRjcUAKKMVkLM6veY1b4hsyVPTQkd3F6jPW4+mDWZ41wdgd3Lsmgzx+zus91RX
5f+1K1fQlKUVGT7y5oEJXED0RFaDqWlWND6XMF1Vyx8ssODa/s72elCDAlT8JleSzoeOWhwD6pFb
e+kO3LYTGjt125s8QTEXAsG+2jcl58O76a9q8fjmAuyZqnwMihSwcIv6gHBbyjtNTElk8WrY7SfO
AZuh2931NCs1KbwoXT6z1JZBR7xhoiGey83bACbSsbljTCAnLZxis3nizi9SJcwCRbJZeG2c8c5t
GB81bmeINRLyOf8K06wY9uPbjTp6jKukdkOjTNPwMBP1ZShfVGp3Ji8GGHh6ZftS4GUyKZUNi21E
yj8cW1uTCKF1T8QoxmrnUgifqaPvCab6k9IRRbF3asrtGvAbEiXoM8j16X2G7ca5GTSP5O4lyeE1
QLY6sARGr7B0686OSfLGH4AlGk5XEmPrPvC1OVQDNU8SUos8VWDY4+verheh26jzZ5yk78dCadZD
Tp9gkUMCqujE3UCZ8peipyBmuAuqn8JE5d5ONwfs6jJyeRyaIVxK2ayJ5paJZKNe0bNTP75EFfj1
cNUSokzaB8//D2n2OkURRtC97CQfOiyZcgBi5ffMJ29f0lYEmjrMYdjNJnfKMv+stxoykjRCDHNn
rFeHydeXuHnmeZ1maBOqOqJy3WSu5ebrqGU+rC/nV0F5kn/1Vl/0tkiQu7wc6+dno18Thmhe0cB3
YYwkQrG82FbMFUpsZvkoOlCuURgPzP45QPz9atwX6Kts5e4zqb32vBJd464B7aB5QV8Bt2raNx0i
WOorgrE3rth73+KAzT73g6d3DwPFGAe0fFz7vO/YRQuoqW+R/dCv9Ydk0VeiYKKhL6SfG8p+t83p
368ZXrTyaL+leaWtoMe4yYqwQgNc1KYwicIAoVfqCqVk7RBjtrTq5O1wdVyy4oUbflPFEt+RJARF
IVxW2/G2wfuFitaDVomAYqu41tHOdAXM5yuqv0rfxWHkHUigoibzGgWBDsL956twlaPISCZAYjL4
EkHQtypBdJOiFeAuGbw1j0v0XB7jNrkXAqDN/kGUUClXE3IkNpd8Vpc+h3U1raHTizNwl8IR0GZb
Ojr4Cn0MSKQVeVfR2V6QirZBIKRxWr3f48lvIfikzwPKDxErEnkuFZRjtEE378nSIaSWWGbi7Z45
cupIsOCS1HipqDPMJ9RGqvJltQhXF415Ek5+0JMHYNwRmtKmQU2u4YDhx0dX3R6E8dNVLFxVFJ54
/Df/AKw7CUZ8yMYKTmChc80Gp8bDn1QgBrl1yxB1Lpa37QIkjT1xZwu6NgzJPS9JRZu898SezsLf
qGnZUYnUg3At5zHO//SrwWW9YO6MYe6OLVzugkImDTLDif5CfBCG0m7eQwkqfMcWhC8etEENo9Ug
ssrLwp1D2KMZuzF0ZNYCi8F/Q0bYtDSTj56ag+4nZb9xQveeBH6dm9rFIoivfxgL+dbktlkY4ATm
rooMwcxvuTImN/trm9q4fyt2zBNyBXP3EtQ4IPeOgjpl2SXBHWynn4PxJFVUOl4Ka138oP6f/Xm6
5ymmeul/SKZu1wt3Md/PE14XRrU/AXIyMAIkXP6npTAlg9/Dj/R4aZQTYQ5MfZ3RkIN8S+cITZ7X
BgVxhdHR83tjFCukUptk5Tj3wCCm7ohmaeqAEv8+ll7+n61bcIqJWKvVKPqYp8y3rUk0T4Hyia+h
dCi7yTTsOooWxZZCzOHBYSyqd2i9GRU5bw9RD00InMNmj5Crg48KwMLaofNernbmix8RRlV57Ep/
CcKdIZUaBU7AyAZDVPW8JnAht820t87hdytqpw8gonvJRA1rHcTk2nMU1dagUHLnhHsW7EwGzZsP
nSgOAP9hW8x++hDWZd1THp1JIPTRp8pswgLXqr4Lo3xeii1tMecfzwOvkWCYdU6RNcse+xUNuTEP
M660ZK0JpAxBkkqdq/U5dbvW5zlbqP7H6YKsxVl2yQU5sbRrO/+nU9yPQPK5DAr5Bb527y7g1stz
yUTjIOTdwe9+YJQGUJ1eFmx7TRH830N8gh00wonWhHfjAMhiV5aDZjnbfE49hcQdDMx7Re7QvFSm
sJoFsNlc0tGzivpxBekkoXQ8+G9GH0zX5tx2KsdZ4hmY/flWHAIvTXNOlGrywYCF7+n4cVYlkUEl
4FCS3NTMVjTSxh2QXDd5m6v96xQeXMXPwIDRq9/pkMDot2BahLO/a4oU1OHYBv+Jm/JfWCgRt73a
yyrIIl4jOZgV1hr41QFx6sEH47Y+uWCp7d1XkbdTJDL7/FAhfvfSIfEOLKuLtARu0bwhnahu5Ek2
reESAolqkIrErGDXSI5apRCyRbLFBa7yjCWSyimfc3ek4v/ScphagrcdOZzHjYM/+AGPZ9biSy6e
F9mKNEsYYmonyusLuDjwm8ZLX9DlyCN1tBDB6SaAX42OGB6zLaD/QEUINNZek/TJZS6lDxCTkWZ5
KVjLIRfvltqzTlRDNP28Jy6AQMTbsn7WhVs1EJIcRJKd+lsxESoYgt5DdWrH5UVmHU8E73u/dETf
sCQWlymbT5DshYz4Yzazp6vAp5hd28gfzGGN2ApKuX4Uvt1vDRe/fzh+xksGxpG3etg8nsbhLycf
FzCLxkCI7S8YZNByLIjyubxy7B9q16eGikZ+TNMfd+OS3gB5c4RxJehdGZsckCTNryQnIMJVRKru
L/trAGl1F2f05w+teLeQXEI1D2e6HtouIItHwiC1FZg2dqaPrZad5lT4tOHkPiunKDdt4yhmxlhn
4ZOk9AR16ssLZqRfr+vmQEDuwj0qI2iBt1dZiBkOxvqUGDNSAxbryJJfct2jx10Ac0M/jRaWQmZR
blqsPvnCVHJoJthJtwL3+8JWimi7ouox+Qy4u7GTrv+Fz13iRjwnW+0k85y7GQ+CRYzMsH+r2q+n
Xogp3Z0vCkBQTWuDT2N9WUYK+sCRrijuYZOz43cqUtCj86kz3myOTzJ3Fy//blGeR3HleQ6KCUE2
J14J6C9Iq6j/n3ORreNM7zXpB5ULiq2SKiOhNojj5JDgTYt6a7UdE+IkCeTDEj86wY6LprAF5Inj
tJS3QoYNx5BWfZwOkpbjRxkNewPImghzsNTrUJq/st3abaXz8fcsfK845gkszJXouHCJj/S/t9D9
/cKw+i226Akru1/umjheCGY9ihyCuEdE7ZxYmE1e+r16Stw8aj8lu4V9XZHHudAzRryy66xRdptE
QdU7ePQpg1ChwvF1A4CWlPuCSIayW/xumZAfkSs/8AKw2fISuLbp1DabfauwtYrY34bnyHFzwxDF
x8cmkwcPA04Lgq9rv5ZN24woEgBoEk+sBPy4uGfid/VN5Oz7C08i3Du3f4Fdmx5qgVXtuFYaraW9
d+lzWLUZLJVBinzjNsP//9XtsZET3Xu1yTjdR3NETgra7JOzxp9EWbWhSQ3fKUsxIuZHewhWB2p4
vgtOWfgJlPk/e5olox8cnMCX8X9UHx4eEYuxGo+z0edVbB3WZG5NbGDRTu4obAfO8z/iN/rof1V/
NtczGX2DuvLOxc4M3kNjJDpT4gWrESzPYpY+l1Q85KN6Rii/4477vsSMuSeBnpBLbGtBvgDaTvTY
HG20DGiCsRVnGbXkhS7xix8OVEcbHp7G5hwN3SVQgN014X5abQTqtQyWLBi6twhfldvlYQQxygW9
6/jgP31BTZL6+f00g47ZC3xkLJSxnqb70ZUuGeRfpazFuyyogDcIRkIEzK/8V7EhEOpXloByEvJ+
yBYUEAy4Dd0zHQJdow5kf7U4BPW/PATPuHtCsgDA0/Uc2lxPRy/BdK0Ve7NBLhcHjJclPYopA74F
gwMukIZH9ZCV7cIJvdAG+adAElxqUcrhlgFdtQglB2gNTkrQN5NaUbfKytH7lIeGn+FZ38T9N8Bv
oSslcWMDxndD1t92FtWZs0wPPWwwzTTMGw71xW1ev5k8k9GOpta8VDCAK9ox7H0w+OdcxNmlTUaS
Uj5wMENpbsaqP7L5/J6FTA++eGPzDSevHVDmm1QyVy8d0IA3zBM5nQBPW7BrF4dZbnAAf0XlWieN
xZu36giKHx587OW/74DN0ykNDQoYOKWAJMM9he2vghOhz3+wQbraX7TiS4UQf8IOqqk4eqiVsf1s
CP0ZorRbyYDeMOt4gTmTdUGd+hggZxMkjHrPC4ZwkJ8f4SMI23qDFhQ0tHrPoYGbksjl0HMm0tHV
/tOii9tlxoBXrhjPI9GjkGA1biysO78c9BNVlpSvj1A006W8Msv1Q+Df1zNi6tmvG6igEXbK95Cf
F5lyc1k0+/F6YJ6ur9k9e0a1FTOF2TRbAdAMd267FrloeyGUAGiMXorB7SpUzYKbcigV2B7FE6j2
WvI20+BGIG3SJxbUdMjXCzdeoini69qdToq8rlgVDHMjaA/VsR4cWfn+m9IF7UuZO9eS76gtfHkY
3CZXDK9oExjGKGVs11TsGvnllhBRfWWqXYviMiX3A46JrkWnoHnHpGMm4uD2lx/grFtujhB3dPHS
EiyaxsUJmxvGaaeEVvortyVMKGcPpHOLNBTaZcO7i2T5Sx4upTn8N4581QdIInl70lAPr+B5UVWB
dhP1G97bmK8sIZ1jEwgdBeraCQhOnn5nzOKZ9ihYeosX+MDFA0+RettCUSNbB7gz/GzaapC26770
I78/yAoP3bYUaUTrChZFZP1fO+r3gRSZdoTGcZpW0QPVSXgZrRYAflZ59onfqbLYxGRJnScVdppR
cCixqbc5rhDfQtcfjo3RuIHNTUmUCvIGVWBqCV9uWQBM5V1/ETQ2S+y5g4F1rBEbadv4hAbVFr0J
NVcH/SrS0k+wfaFkWYzRluEsRHuZjArxEuElGuP4LwzjBtBCb7EpsI/oOgggdwNj1C1HCtuPF8tm
tpHl/IN3x6vl4a3YjjvRRdfNoHTCRqIl/3ix1saLPlBbQ/Nf6zdXLhOai6YW1t0VXNwDclGj8k94
zFtYqVjaTrsTjaOT9S+F/4e2HAckcRZH3uTmB02iFxphd27Z2FYq4cFmpZ0Ikclefiq6my4p+ccG
1wjW+c2RIqv7hNBJwJ1YIpYZwqg0UFIbWnrAqXBxbH6gpSbobJgJdVuAaaYa5jOpPj4FRGR17lGp
R6EgldkS9hb8MznH5m67e8SNfwhT2sRHMv+QszhN+LxFW71uxOnpMzWEdo2GQnH+rwpdGLP0vpKc
srBxyypmkSdpeFocCDQYK4U8yqR64SrISKDtYEKsVsoav2/scgceLWoPG/iYO3QH6KSlnnfD2FAQ
vV4xdw8J+FjIaajD4GIF8l++nTNVMc1P/XQIfWGirQkKg8OPR/vWvcVbY1qDuq0+dHo4+FqJKr3L
tts9wO9azpfPT7Q/e/xp8Xzzj6u9OrzXKGIDwWVCzhlMt7H7PSH4jO2gLIJdcKuBNcANzxHt87fE
O09EMNQWPC2ggJeXSx+KGLd/q8qIKharfEmBI+OLqdhicKRMYdmTHMCH5DLHgRjCThs1o95Nr8fn
sMrempL8f8XaGmtDZ+2HDXJ7V8SBxervsElnZ40SGqe18a/pQtVnV0d4AeAPwcov9WdXl5oKhL8G
NsbCL6hQBNx6/Kt5gZLJHrfwUs9kg6RC/+9E27sCSHU9CZjRkYbcXKo6kgzOqgtolvsYSu8W1Nlb
fDibB9r/yin9TbXzSD6EjkeBSn0+AMtDVAe70bKnj3oWD67Hzg0JF6ctY7xvC+1eEkqiSJ/0160d
jWaMyeSWEnd4/IiTdBltD2ivdfkE6Qdox6bAqlsB/rfn6SUlnXSHKSNFb1dKLF56AwJ1mkGMgATz
wRxKjajjmsP3x1w7O42yvf9QipOcRIBOaxfXf67XciLVzb9TInmXEJNqg4p8062bjSOjlXhiqRVR
Zj5+cSEfY/jVABdMovxHEzVEzQa0zxF+hRKptdffNBQpHNqalxW2wWJ7cj46qVD8/ySt8szBETnX
KyE5uyk1qaRfHvco5KhV3KDx//TOH0R2lqd8zK2Ri68XngDK7BWMaqBMrfvZsDLci73EFi0fR0y+
6ygx9urPCCf1PS882BaxbQaC8AC7KEhelUaceNpuouhKG0urNo2BRO0wUnrlM1jIxrLyuBXvzisi
iMU3s1GxB7WkedZX/5DodmHkCzVgMbHf32kA/LrtnVp0XFNc0IM3tkrp821X6IgUSge8BEe7gbs+
j4OgVPk/JucL7ig4ea74ikyaZYJESFAjlRQLvjeycquCW11b8lCGpc48dzvRC/THOaiAjhjojVUp
cj7QdnN1O3WXa0N0DDuDXGbjfJzFnCpq4FD1qTv9cSnLgQju8Lk9TYvQHP3MqZ1QNhKjkCEIxRzR
4FHmdr10pyWUGnH2Ad37XDkJFBGQBMPvSnHA8NeoVkcGCY4W10F9DiFsl36ZIF7JUdas/PCpmEqe
ynmbFpjIa2E+Z0vC/svaTxmEtWhhCrT6COwmvoY2GkN9P0TairiCtFDB45A/PwBVkj1d4GUaUANU
qysZIMIty7JHthbIBg/PKLV3M4pMQ/+px9SUfLsr8m1bkWPWHnnTG6Be/ZyQJtAdFrhCgXAc2VCW
gPNAGdwOvDjjbNS6tG+zLndIyfeesI5QbDl3b4hr+x0BjUplqSah++X6qhEBfPhFjNLjor+HfOX4
FnZlu9KPg7R3wleaR6yJPrV8Jnw+ztZpMwBK/u9R4QGavaFFPt0WimmzNdAFGvocOTDAVRBkJsc2
ilkWutsev0GPrribTLQLBJoRh96ZEg0FHg++FCqMnb5ksd6r7Sy7rILh3iwQkYyE4aJQ7QjhT2ed
rJTehpIySHWCIo8BW4FS1XWYhA4/WIAOTV1HWjAvJ5J2lCzP932rT7FtGphBcDLXKiGkRUCisKc4
R00hB/4Rn5pg5A4tEYM3Q7vnOoFxagg9ntb9ULwDuwua5TBHf1hTev3tfzWDYn2npBgyQPKVcUuM
O9sg1Ma8vWLL3YyWdgNf97mCbPJc9Srl1MeEyCQ80eqf19EOsDBWvOou9Ky3qK7WVOhuL6hs/62V
gWraYnbTqhumL2GIGmigjkVYzdrdhJAIL8xSd0bh06Bv10zHowvdM0nhnObZU3mmlx4vZd3oOwPX
xiTceVbj4TCkU0uNqc90qigZh921Q3gm66MuovwYY/7nzs6FenahDZlKvVlvJjap8KABgROhWNAr
HMMMvSwKprdWOnSLgZs5OZzcLg7STILfDk855gDYUe8sn+ZQ/+5buOpl0gO1ohFzE2Y7c85n8Lxd
ITwRGZ2QYyss7Bm+09azWoddaL3uWkeE35siOvLVhYkp2ktVdz9KKVnHE6cNZFELPaWXXUfZ4DB2
h+gtDaLKJKRyHQKeoBS8ym5H2U1ZnJySzFtja0gfdZYxAZM14r6w0FTKJinFjMr4k5FuqzjJyNn0
zGhsKFTbtymDq73M+znwO26eg+sVbnd6rwIJOKn5MXyUe7zoeJtIbZhiTQOiznp+1kxVeLfZCQpl
vp1UpkDqE9pqSq7mZErt+PBOk6QRoTR5lDGtOqkNwHFQ04Jp3d66e8rWhx49mkc6tRgYy0eR7nqU
sZXqNDVY4jIBDag2Eggz77xtJi1sbr5f+LDp3O4Eo7dxVutRB3gzXgV0uNKeEXEWF7o3K08eaSsC
P8t1w6ce+1/CbVhVxGkU1RPq4oCnMDksK8rEV++cFvC4Gb0uZEWrwlJz2QrrdED7YwAEwpO37Log
C97bVmaMCLYZQ+NzxUEY1TfLtSIf961WPremG0ldmFb7tkAeoFWwJrJd2TqAkBgxdxFbeeKHaHwk
XgF35bhmZFuGIDmQ7yh8exK8MIxXB8xdEbr0Tu2lX/Bv0oCecVWp+1f0SXbPDcMYLvr8ZxXgYBP1
bt88L3160GZplOTsS0scesxTaQ3pTRQacmPEOfiq24bOcrtIOy8kqUptmBRYhz4tAaGgfSxOYc4V
vNTtnCvOE4jPXrPxAq0QxN07XjYwNx9QMsI0t95YRekE/CjgD/Knl+0hb2xJv7aQDeskcSLoEYQU
LzJhXsO3yAPgtP0hbL4E4TqEXpZC6oF+AV5QGkC7O4uO68m7Xe7V2Wd51l/uz+DP1iavFxE3Py8l
UhFk2+1YG0m2wnFeNTFiFK4vSyD22+xvgp1F7y5wMwyXDJvKvMWkJHsQ8e8WPvZ723hfoo29guPd
trnBLf+ai8eDUtJcKQgecSUOwjhCzNBsyBC7P6agh/J8Lm7bkdFziD803DL/jQfb5eFsCeS9Nk+0
6cpm6WUf+Yeoa9mfJPHO8Cvyn56+hSznut70/ggESPJ9gAh7TcHkQFdsArhlUdhh0FfqSe1iQdh8
Zg8tItvJMB7IktKQZ86y5JVvwUKhMeiV+hC7DnDrEgIuKxHILHIxX3YxfdmrLJP0MIsvjirYSD8C
MqAUCKXdi45tWT0GBv90W2wvyg3tBlwS+kTc/UvxNidvIKBdPZzmevIwpWHUUaKh7uGodNytAWGh
VS27smJ+BjjVhabO6rEzOCqYGwit5h5trlX/07lWiXNkxrdLou29cb2F8A2zrelel5KOhOQUbPGE
vDaiunURrqoAlATXYQqe4sRQon/iocs02gXWE7M7AxkyT6OPhVN/sRM7ZiHpb05U0rsqnDxrF40B
kOmQG0sZOQMwHAA+5q0XYA31GdMAhE4nZMMNRyINw4ccUNkQkkWDMgQzSxRwdTpVU/KOqOgCyf8Z
1EMaj9H29deaYDy1jnLoKecBM+bEzGxmJmBHXJ/35RVbue3HiZU2JLnScVIX6wVZ17mvhgcov2kr
TwCt15knFYI5wt7shCooWgx/feFLth7U5hDEZZ3emhP6TfdcLzcDNZMA9uWKz+ZsmOQJEzWiNjB0
Z9fs8J51K0zjO91avfZmLMAbIzBi4uOLRNuQhFebklCXCEzgqC/r9d0kjDm25vL4bJsCvVxLU8EJ
wMxCAf73jBU61I+HKJLFQ05CVt8uvDqhG/A+yDX2WCoHhEHGFaOhkiSrV1MjYrhniNdLZRBBZOkt
vY/q4Ca7lglevNMCwuJUuGhOUE+T13IVZb1TedzumqWCXqdAFlpLDViXojjkuqguHXqVoerB/bB2
7fHNvlWAhjAvb8oHkzsqY0qPFejZc82Jqi5omg2+rB+i/VKcv+W106TrSjoUw5+A4FqrbP2StEBJ
ZSxnHfJUKnLrx/RAPHTudUWCu4fSF1q8tJ/h1+LjyuuMOfELgol1TexB2LXRCcnBoGblMmQ8J/cp
SOanwZFifbiqkKXcjMCX/DSIul6lNM2PDN7j/WLYwsFvTvr8XBb9C8RYsLkte6MI6005LHd3N20q
nEEPy/qXlS7qZc2s6V2L04VxVl+zbqWG8GnpAhirzHLA8wnhje+miyFZWkiHeNkrMTivCgy7ZSmm
+b3H9ZfsW1FqDfAxX6mA/Mr9dEJYjAlZ3BgdakG7YBjowGUE5K37pm3pU3qxsETDsNTBOZBmLU3L
Rmux2vWhAi+kixelPF48aW9kqsEFO/S3iF8SSuHL0j0aY3cY2adMNVfPUGEniRIfIYAM6H2MQDNJ
OGWw5JfYpxS3Qns4ERAUf7HK1Fp+unahxnF0i2Wlzb5hUSyjdSRUIGjzcCpOTodC508b67ZRTf5Y
F6+dsy8sCiDNoGNIQrGirBXDyDqVegu0c/+blvhwpH8snhz/Jq6dleW9f0zJZ9e0lVqC0Ny8xB2h
83B8Dlj9IKzvbafjSdN4WcH8gq6BaM1N7a7P1jeKLBLbzQyU5HdQeQMQNLuzg1ipzydl777DBN0E
IQV8cyI5GygeCUpAQE7vT7LEfS2Hr/+oSuO+qtnPYTBIa1vQ+5dHk3gay1wQO2Wa+bpVXXNIQmdW
G3lglmWjdFatMLCxYaYxetj07GTIfGKXsZZI9NKmT/MH86zmbeO88fSBvsJgVJcDQp6m4vAblHAd
SlmlthaMp8tw+ECYoBK9cip+MGLZgO+41sRV3LPKIz39qi0uI7zXkQRtPizLBk7J/3zyN8F00EdK
oVTtLTZ9OE+yDNKUwVV3CZ3Tsa+lasRv6p+m39C/AHds31a5MDh7gsg2idRFbjexgGtae7hUgmqF
6Qdw6Gb6gi0dUfHVtJpCK88+w92HSBauABC6nGnNcky9aNdMSfrreaFy1xrty+QCnuB/u+9yoB0Z
9BeKnmYgZ/YFTnLu4oFysGW3TWAG9oORpypt8PpW766ZIibMAO9iZ7OkJwASwjOMPkNxympjhKg5
o0ViEOqiWqqgjS4tWZSofKKJLGlm9i0yVKE1H+ZFRmAN9ZcqCVT5R7TamT8k2ez7obbL6HGQDCeX
IpYiLa/kzR3+2xwn9ZtZP2Hd6KmIOhX4UNh3G2hhZ0abILyEwZr24tVsjMzlO8VmS2TlZO/Pglkq
ciAZWL5XDk4xoQIeu79c5WUUWE+S/i1HgYf+6C0l5kORhUU4TAs8uFUlz4B/+AwiETQP1UYGUXXs
0yPVpYHyPdgiSfZw2g0gDefwAPRpplSpV28LdeN+mKJsjZ2I3uzAqnM5hFbJLE+R3fN4AfTmllck
JFqcL4WfA2PMJ9mMYFIJK445f7hzlmHosdd0wHAGzocDfYHd7zXhW2Hwb6Rah9SSzAdvvMbre++L
JueKQUadcZ9/GFG4uQPvsDlR8owO3srEvl7qX9sH5DXztMt77Q2CLyHCTb0t1eRCQIu1vZjwuuh4
2vYMA4Uuys71VSFOA6zScgVj61Ig9r0mRYDtv3gJXV6RtrqMLQFoVrwq0JSvhu/JJy1Ov+ot2l23
KQKYO5ivTDAQuYzuOhBWTuUz2Uu84yb9FDx75Hmo89dnFKuhzQJDkD7/1IZSn12y9cG6wcmMgg+B
qTJqsso3qMOB+uX9eTm+Nw9kRBVLpA+VnbLQP4ehgzvLxTvmgWE4CASEptqI9pfTsCM7NtN9T/zz
GVr8GkUfKgeTcHUwYefa2P+8Jjy03I7LOLPMocSgZXgFi2gGhpvZVHOFcUlvxxZ+ESYIANQGU8nh
vIiSNgySEWnQeeta93uEN+HCpMl2hSuenpvDhZyBms8xjTw8AozRcUSUAFN8r7OGrEIYTFd8fcN1
T7YlW2+SRheKYjw0G020JZ7Fp2SMoy9tVhTFGyOyBwZX3mwuURyWe4bwAuOXWUGjo0RIPYKdepHg
kV6exL9hypnrRzggj97lTZc2U5Ql1o+78zeeHGTHPBSAGHLH8Ps7XfVtROVZk/XK8Cp+sUlPKFTD
TvEaiq0VDbH0bHhkBDk9KldAa9uR8qGJ+NwhpG8k+GW++lU1NpuGGOEHTiTO8/dUCY2V/8bhcmn1
f1tznZR8qN2APl/MmzFXfhI/hw5jD8x+IYErVNodQpEBiThW+oNMiHbvVLTLMVh+dBnTqUKNhOMi
RMLhoycMNbqFMgaomEQmLb8WUVnN5o0N0MMcsuXZHozzVGUHGb+qvTzxwGS7TFXyP+NJCiKQ2gk7
UXEDbzfqqnhmm+7ZeFGfBFiikptZO/5X68+2apN4rTjR9k5TYKhWoqTJqFSdPFru/TmroDfS4TDX
ET0zfsn1kw/45VQgxuw5xkiDJm4Soblm1DpUkpsJf1PjO+Iwz4d1DoXtYcZZvVbcEMuJXDnrjLxh
OsmiIv80iWYmCijWuuY/Djy56+fgoSIkNVk1ZDk2QsKDqk45v4aQ8/cmU9pT5YAFhMFfB8XCYgLm
6PoHJvCslWbW4HeW1Qbd/6IPOfLuZTOZ93I62g/X2ONcdO0VRCMKeu+/kBqkrLqfZN6M8xAQcXLp
y9G/jfCZdSBSMioguRtamtJeNh3ZTEUJqbNfXuTMvnuJg8QD/iT29A7XqoJwdk+KJFan31P14jH5
VzrHMHHQooZjGe8ao0yl8z2EwUy2ktt7+iosmQokZdEWwrSRiIHFThF2R5UV2tW73N6KSIj+ioYd
Xc2bTMIEiED0QwiAW8GHkNwyJXzh1LDd30B95IZAZb6WCbTrXwLyJVUM3HbRPSfcMP0TQd83YdUi
dOmAXGIo7OznaSgnlWxpN7tA9k+LNw9bsB4XOBxjuhZeiSDMrgAI40BvEpdHVon83Q/gMTR4e7rU
ckjeYWufMLnwjycy8mADg9ooFsybuCBxTiHIQEeYkJCIJ9RGKj93vCpHtezrRuqzYoGUBjZFbw/g
zBpK/jsNOfuWxdEAxa7Mn1hQeOuySUmGVySP2dxziljtmtyKIOEK+e50Hs0xC0MLuNRwf/2yz8Y7
QUjzWOWAIzVM9R22lpaV9kPwxj9pt6PWZmgdzybWeVdOgjknmrM9j9e5tU24s4KnlXArIy4l9qbG
v7yDbk/xZ9bGhy+YeWG5gwfSSoxfMMF7WbtTzWHLagxN4a4LJzKSMAgGUiNY03MWLgL3nfu1J3y5
D48r6u8e4JZs8y2bsX7QEXUxtYB7mWfW9pufS1q/pzuy+4PrVCProxIWcPk3VokGzeVp9KS3Ntxl
ilS0K6GARekj0i4SBNH47ZghS/Ar/y6Y4PbvNhbMS/rpesObUp4jINFR+YCidpjqVbl82l5AHWzh
6LZcdRBEhXEZEjwuuZ/AmNpmUzD/Wu+BrkDnCCitZhZuju0PZzj4wIo1OZmRfLy6X7gwt5WAVV7o
4AiOLbHgP//ndlUdIA5Yrtq6NJRxzK+0fJ8m7mrKjjcNx0lv2A+Of/RRPPYKKpgwLaUPQFvrZBmL
kJRIZ989BFyHMtC3cXBNPTpASTgiCkM0/63mJKUc1Fnz0dvgR4Jf3mKxvHTqIA1fFDjoF5vfDm8S
aenoVwzQ5F8OvGFt13rWv/Mr+jFG2gh95j8DR0tR9ULbdITQWRlsHw+dWxx03owZaNsp7DeMGSpG
CmBpKV33h1QDTN7PISrEXezi94JM4lmonNqjoUJK5oGqsNVfpillRPOxE/T3LtoD3f4fZqth9zw0
nVlHgDAbNWJQP3GqdIAO6mZMFTqnBePl1F+laNGYsnlfJK2aVHMcWtkmQfOpX/+25POB76wrfcKd
Sz+Qg/zzRV73YjdN+HRrAsDaWT76GqBdMqh1fhLh2umOl99oczuT6MxFoa5Pbb1ViASIVy3sA3hL
qix9yQbE2uyGOdwaemrAjN2fzdJvLoHyF9pHJu+i/eScthspa9QWXpa50Y2v2I20jYCgzqd6aKPd
q1Jkj3avi3Ks5gTramVfnkvX3IXX2AqEPSWFExUgBThvppieu/aTfSm/abdLdOwAKEPPH7tmER6C
r1lKfuxqABgfE/kzrTencVWlYvG4gU0OtNexS4FmGm1TP+GtAR0lzaxKArysuTFpTzXQYsXqFQkm
xieziyMXJc1LMGHZafME7NseL3+5rZmazq7OncIlZBeC1ENHX2CDbKpyCzyZs90JPuKHnLguJxsa
pHUYscgrjn5GEn78umFU3S3k52Lo33KIC25Z2e8fCQ8qgAfoxaROhPny1r7dilDmtY0YWGLvrYb0
JcSwk9xTmt9rFAfO1836bwCuCHD5L0vjRW1NgULhXFZL/uGMprBasXIz8UNf9zzcg5iBzJYpo98p
3kxkVtxnX60NAJ5x2+RbqnZrthyWikTz8Po/rX1gDLU+aeFP8r4vxT14KTjBZWKdQzblRSP3g8jb
liB4xv6KdMVu8rjB2srdCXeQrhHoZ3UvrJY4ScRtsRC5k5sfDGOCHH/p5QCBHP4YuHYDsRRMHd8k
Zn2sPz8tn+vYHJ7q0T6rFMp/lw7Iml2WIwD46JqT5d9/T8kehTo4LSbeXg6SjuNeDpGbbPb6Y6H4
FfFa6I2g5f9f/xtp9X9Og1KXPMZUPx7W63rRcAMgzP9l8KMmgsweSYhoUugZ8kYxzHRzYxIsAD7/
t8Oda8gn0g9oeXAspGsOx57YjM/ouS9QynKO5FpdnCRDsxOhz0m+yrW0JqMcZo0qEKUSuTjnOR/6
cRwdIXzT9jjb+vuRl8ob4Wk2vrJFcd4wNYCyOrf5F0jpYLRo4Cb/W7cidHCi9+HIt6XeiLys0FH6
bCTztUxl0MdcRqOiAZei/BCaj74Tv96FH14g8PmvbWDkIV+q7PZToV0DeRAWIhKFwoLtKJyrpXwN
bbR6yEwOblJDQ/JBStCa8TwUEz8hsSUbogPOTmVepu8U2H6whGnkCpskF0WQ2TCbRhqF1uGHZgGt
GtXweTzSwO6lpKvT/dlvwf/oIW1eBCsMFaCrtoQO0QVKL4/ghFQcUXrURnU+9dcCelsM+knN8rRM
M4jQRaYY1ZPoCrzg2j0dd1sjMCGJPdtD1x6jVlUnLcQaM5CYgjKBnRM4fPN2CIloGW5zqGYhurTc
jFXmZYxbei6BwyxzMx1a55rRFHD3Zc4uz08Xs3dGQ+iwkyYzzxIu6oiWm/n+UU14Vwq+SBDIn/v+
jxAv0EFlzva4oQjOweGhu8nt49lTTfXzhS9/4lMw1lUdx/E1fxmGGozGN9PiQxO7kmrSirMDfQWD
cGW0cX3HRLSLBp/GLmO2XG4+SzrktQb+orJdNSMKYeMDeJGegIClLxWT0yyjf7SRc8afBUi/wsyl
1Xi4iqfWKAKl2h462sgDRH/3w9mT+d5Fho9wie8dq0gks/aFL6BK0r+PG8yMUeVe7iQobOGpG6er
P+Gza7x4hZKqs3UzuTi5bn28m0fK9RoyNuduciqZ5kPKUoFARO9VrSRuRg18NYvOQwZfMeNx+9jL
8R3XxyZ+XN+s8IxNBnq2/sXx2lmteCPuTTQ1a2w4GfW+6WX16CALIll3lROZGOSFayq+1s0/XdaE
fHzABZMv19nttNw0TvqzLd3qhqEvMWQTyRNKSZ1NIafENzR19FDuQZa6xJJcr+d2mZH0MtujzaZe
U/kbTC26xwYISpHMf3sY17ZaK+WKpn9v/cNOJkdwN6hY4v5j1NVZNGaM8YczyFS3La54HyP4XLe5
61XxB6OounJGUUMf40Jj/Nb0//HxBXdD0XZhyQP+iN2Z6Q5J1GfoiAeY8ezLjMdkiKG8HYEM+NRK
Z84NzgXiT1iDMkyEutIxI1gh3m7dfJBixlpbaALY3PFO9qjbdnqBq3Cbt+FXo7BjI7KvKi78/aoH
Q37RMbe2KG/FxObMaMmxJ9duLwG3Q6mJvPiNmq2qWTM35f2chqCtVwO1Ft+UU1tB5/iw4339K654
MCZeTSet0lARvgwSE6u3ZlZLY8Yr9cNy6eNxBrhK2OTST2yPRQleSH/XQd5d5EAjEwBPmNAVxD81
9/UgMg2Roiy+OXoCLK4j205Zi+S+k0yUrehipMFsyqpUG1Q6km+mBFwcK3zWrEdpP8o30UJ8JalD
47nCwgghapaQO9pzp6t93VytQY0Z64YmE9diwYW7SY2EkKjBTffMQw7viNAS9Oc5cqiD8jOJwTfQ
6Mt9aYK7Z1to3Ch8bsfb+PEyFt9OkXXKh9OVkni/59CS1/SP9oM40szpM/tJ7NhOMNhjSpH3VD7j
AT9weRFOO7fx2uw2a5FSXc7EZn91eg3iLbZAF0nfINcWOUno+ImVVU9zUzDubiiNpk/+pfEq/wnI
IpB3dA5Jrd/HplWQ4UWQJq2zi9wo0qanmYUUwPivssZqzkfpuG/SydUPQv7x2ziqeuK6oujGXq/u
ZFCwrx+ACuQ4y6LglyplNYDCCWGEekl4KgSQEasvpI5HO90BtTcwV1p/SkZRE3rgQKrQf0JpNwNd
Vq4yCzcH3U4XfqteIG/CQw2EQ5wvD6pIeFEaFoe6y21mV0BWpPhERohRIjhthxFe0jPgoBA4bW+N
OFMHcKVhEg5qZYGAV/5ReaCmpIq1BYE0xuCgcfUK1uQt/PpNhF5MVqI02+m/csVVmqZZb7UGAmMH
Cr3msPd84x3+1XtfftqjYSpAAL+XxS/fp/O3PDslrKDy2ZiD7WK9mhdtjAcCYgRWnGSAJiaBhO17
2sWQPHRc+fZrk+x1kzPtRVHqv9e8thaskepNMmA1LKohnH0+3I3njxIiRw5OIDaq6CuId6wElJIt
+HT8kI+Em1IC469SIbqXPS1inVinwX4pzo/Xvp+lv36lzokrXPcUzg8auWvXHeHrEI3I+oAAOGjo
zl8uXg+5l5hZHDO4IAv3KHBNjSwz2+h6TpcNPCOMSBAShBSIybW5ZA7as6daA12ZIxm8looShzX/
C6vs4hv6206fxg/myWgFYGbtDPw6Pt4zAbSvfGKk/M7md4jqB9kJxdLB5nbwvm4UXnviNgGC7FTf
U95OEXteiBjerkcJkF3iJL/fU+/M6mRh0ph1SWfFzRJ/BQII+zH6wOm4J+NBtSN5aFLMo0YzaJhm
p8mWpJo1HzDMTxHUzrGF9uudzLb5OMhi+1rilnB7Kz2WJezgg6sTmO/UJG7/eU/XSqVwN+Q2fCY5
V2BfoBeDwh25XKak1hHAV2C9zJhtQI342HYk3ms48ecXJ8uHyeHGJAcfiWByOwUKjBkgemb7YyAc
Tkw1Qsx3nd7n7tyhacifDNyu69/pq9inyoSGmh01LPNUW2oQog9CLLqpFU8J7x7CTGql+XO9EbfC
ftEw29Nve9m4y0NVCve4fqYtR29bK/SVjT6QR2t/yEVkznNpZGi0GYfYZyCQEUSnonCYMt1Cpsws
0sIS4ptXQ+6qzfhax35P01wNcItlcAIKNRG0r/v7oz6Pumh4EoANSB66Ktw6GVvbc3jTq3WH1usi
nTK0vI/9ZHD9Rzj9tKUFOQUCZu4S+R0AnLAXfMGTeYZdLvJXZzGbLiUVyxw5pe9wIkGn60+Px9rH
oEIlVWbWMoxZEFwRgez04C/TxrQncjtSjNaCMDAxGFK24mZkc/Ym+jPD72zJgFpozQil1iLx4Ivd
eE3Q+LESw8uHHiX/hhS6pp854TGYTmIauMV/6VGQePRSTi2j37+XEuAftdBoxjV7XFDXFGxfZT+y
LTmK4yShBIexGfmpKkC8ER9Ob81edcPaMPmsY0+R/tgJea0uxSvPSDoWW3zeq9y1I32JLTSFKsVk
jjwIUcyQiqVr8+0b4BETY9io8EhAxOLsnQjGN0SVOl1nMBJXJQgf++2180FsL5VvuYaQfg3Q5ZKO
F7H+H/HRb1wCsv188zhbL1xczc8oMuDKbkZfuiQyTHOnvlIrRqGcXRPU0RIeNEhbkzVLX/ZWdCbf
MMO1sfqWvv3QPFuUDaHEmAQd0Rad1GAixVtqC6fj2BFQpYeIAAXR800YMnXkmiBWVehaVpIkTysq
yu32Ej1j7TUrKyhnWaiMLsQpm1qk///Zq1+Y2iM1KEbesXgZaXWc4qJ3umQxvUFF/vQlt8B1kG5T
Z2HyRiVAq1DvvmWLyT5HQOQGSF1dmgI8lbSvVw7me0PC7pvxBFRSjSFoq5UMW9dqEXqApHmn/wq2
EyAX5byPpfqNvtyQzMh/BVPmYnsTWbukjgT/g/ul+gjRHQeuJTgNRStNatVUTHkYTFA2m5Upjt/8
oY+eT+Go86Qkc5dAj9IkHiAEU9udMNZhKOxerNl6ZTrYUAiFzCL242u4lknjl5ab038qP8woBgbj
2qul6vuhYVKBDlWqj33AuRwvjc2YdL8a2T0MVH+XMgklK+cR6UX6ZJH75hAQjnE4R2zVZLHdKgqs
uBhmvD78mcHfsW8aHxgmipnzDmo657tq+UVOtrWJ3peEfOw7M0n4ojWGqkEuMLGShtidvHc/oJNa
HK8xwTA0GyL9zK/7HzlOTNlJdTS5PwI3pCpVJDh8LHoOciRtyH6qL2go6HhlVyLQLvvLe4WwOrtW
T2AItg2oe/xJm7qVwFTkhRZJuUNOV1dHZuJUxFU2PWuQmYScr7Yhzk+fSeOAutd4ZtBR48lLyrNf
MVnEBR1CMgWbs6yc8dQFS0ScuQ3DMg8LCmOrwsPTD4DNK83YW2RdjSv8aPVPYUM04Xah4To6jMbj
jzfuO+m4WPmq9umPO5FkjIJFOKtPkNczTbbMcD0a8Y8az5xrgTD383Qq3qQnSHUMOlUsDR3meCGt
p1ws6oYioX1RrEVYVpQPN0OiEtBiq2yp0qh+ZGZIn3cvu822i8hT2pR/VKlHH/y2YKCzakkdgivj
71HRL4fUnEJn5IrO9iVhPkfcyrTrPwGTb/ofDGzeb+hdv2rkkjZ1X83UqsiBMbeE9rYp47YgdIAU
BLTOTKZZExx0P3MhnGqraD9OiyJ7NepVCteXi1dJ4sMbFZz1HPtBhFXGWOPS4wg9Bk7LtoSoEWfW
NAdpaHmG04+A2912rrNZ65mAmiy7lXJ1M9nFGkPf0tjeUZdy9guam8HPat15P5zK7/ONdKvuC6UB
R0l+6EEZPsLTW1Bi15nL4AIJhmftg8jaXfd2UbKhO6Kt6f5PhsLEkyDqFjmXShK4qbuLL6zLxWWK
hL67ro7VY6H1gvLzh5VQ32FPq9BCB7kfL7a6vqbYpQMCkog6FSfH8Ie2m1W74Yuz2SeizG9Mp5To
4rhe8lHTEbHQkz+G4FTPdgDqF9D81TV5GiJ4qYvMc4sIE2YP62FHWzoywvabHplKKFE8DkgrAagW
sb6GtB0zAhCnHFUREPMZQTT9fBmnJCoVnm/7FNCp47tB8B2bi9GAeg//iOdSbO+A8gySY+omL+zD
rsr4rnI8+4bsVf+/HZfI2KB30yxlX7Dt6qI03vafsQWs3iJQtof1KyVURCKncl4Fn1CDsJi807Kl
kMSbKmV09xP8E6zw6yg+wmnI/5hpFU972YhF6HBYE0Bv+wfM2LvC+TtMBtP1KzjW0lXdvJkeaLfY
Ceq579KRsOjUjgiF/dRWHMHXgunvxBueR/B4CBYY0dUGt4zzXDTlTWHLF+UW8O/BuL6X7TgiEmfW
iZyo0m6WITyeuytbTdQcIPRGR2KGbABPhIFna22cdcAZlLhkV39z7mvydAMc9cWjB23NXbPDfds0
nLmQW3nwD4zp4TJ/3Z8qGIfsak82RyKIe7mD6AYgMlIi50XETqQaMRktZnmc5BoNgupN+uOTptUG
7VRO0HeV0mwkj/s2rdsjU65zO0rj+aLcy+1/iqmjmI4FldIACsB4cqVHPTFCNMJsiSI1lVcrAo+K
+Fx5BOfSpF9h/7pgtfMOz+Omj2kReOn9TNCIX9lKhqvA00s8Pq/9WbC5xOmF9Y7qeYT32//476BM
EYhkcCLKi6u6VEzM9gZ8jTjMTHf67ep8eGpWfMUeT/S4l4dP/KbSxlj6FTZXi4OrP1mR3zSzYjKU
Sy0CQowshOpIb7GzT0NqPvTUeLUP53/CF9258mEn6WYBQ5h1dZUcK0WuBoNC6VJzy7hEKhRYjmcs
DBtSeGYrwXgDQXbRAaTqnFs/48acAGxKSMgXXPZLJYgel7ONOcFtxCNjaaHPSGsYtCI+vAWDCdzu
ppwTIVXIHqdqEuayoQ7X4IVQWWehL6+Bcl2z7Cbvnnt3uaxGPQw5/7u2BlFdpQviV2v6VZ1Q8QeT
YI4fgLHFoqLj7D8qxII2ePY8CSN2/Bf4ub47dD6Ikvld8uNJE+rVj5dcJdm6qO21UQJ8JtdxV5Dj
ULhkI5YNppaWRTerAUr+lOoG4BIXCQ8M67DFeRlaWJ/VadtiyoMSq1iQYDqeIGtm3IZnk+lMWBeZ
Aiz07E9Bv1iLUkW4rO5XT0RZZNPV987hkj/pNR3anNtD76uy+gGv4rDr3Dpuz/RrNoAB2LDZVnwO
zSi2+FSklj+FRFNVLiJSIHHqowJSJJQ3r7AOxFU646Hf5DI/nARjhBgmJb2/sXOIMI+1F3rVQAhK
m5YGz7AWWkIzGzDBuP90XRV7sLcI+FEb8h8W8t1wGl/o1yQmjCwkuBI7gWkYMBLkiPyGA7OzMHMO
Re3Pu07T26yBuiWSL1vJb9Byfx4jD0fLhl5eXggXL0nu8exBYO9RLF8MtDCIMNPPb2OpvMy7BUIw
yVN3lX8Co2tWkuGyPqoIEpuHvTh5zzw1fBMoSJ4I1cp662q/rmLeK4ppNmstLBuGuEBDPUBoA9Nx
dxE8umNFghoEX4C00F0bwczbHALWiHHnwzFQQa/M/6S9wBamm0aVFe3JzrV+KkPxyrhoQ50uJ6g9
w4hFLI/gGKv0HvhOZDI2dCyFO8FnBIxL3S6UhdkZpFiMyTNousQ/IXfx3IIhoxIYe/QaVmUu/s1q
A6Lr2n/D9lkfxDGYdLpELe1FIe4rYVlE5Eyeow756/nK/0/a+naIIxz4rLuiXL3yuc83u5dmgl6t
dZmiA2zEftCrFhlAOqwX5KNiJOrjq2gIhwJsL/teU4xM3OqySlycd7b46SjnoR3Ui0p44SYglCiW
fqJOfbfEGUzjFF/SHzvyNng3RVmsfOCiu1rr2w9mLrRWDCMglw2fmHbimRBVvsX5Xi9DaDLG0Wh4
qsBBZe0q2Qbzybd6pm3ZFjMKDOA/1WnQ3OHQQWOwFZ+Kf3651H4k5Gr2FBgs6rj3HstotsXgCGAp
Z3w3pUJXX6uGcctZo3WoUZfpPeF04U3PRIsrLeFz8sl+rAP24KRptMeQ5hBm/ZcdKxtqE213Dty7
wonYBtG/lqako5OUyc0sNbzmIrVajZldI3EQh55Pik1JAZleJBeWG4XEoqRqBrmSVkvr190WZvCl
E2BQr13A71hnAvNfUYv3g3vWdoTYShZ5ZMxqelnF4tAFqcIbgCFry4EzioPOQhLE6M3iKdB2IMTk
MjOXHAJDgbEbAUaac9pXaK2tSzotoIwND5c2yQyfn8F955Y2S0ouOWtJaw7Bgmn0QTITJFq7IZHo
RRDygSB2Gqxxe+9aQ4xU1CxW451/of+0eUwf8YcW7vZPAcZyasgoiJgmU2pelCugouVwl1k+YFfK
l0DsFI0lj3fZ/qnoHu/E6OkhXV6Fhd9/HdwFxSZ/qPH3B/WRMzLS7jJzKfP6gMs9a2gG79swER5x
LJY2CzltUQa6mbRuYYGbLixR+i71NQe95cwD6idfY1Re9AncU7x8heCYJGO7b8lvQgGmdQN8nESU
Ns4zkndBCuPpKao0jLjmIYWBTxTEO25vJAPA/V1Ei5mGMQbbbCNgpUaNvby8mviBEodbXeSROyp3
4gFg6nAb/uWGZVNmYqdoBInSuZlr0obYKngwIad9i+on014AKVifyMvJy8w4XDYdUrpYmXOpsoPO
DpsCk+Dv26fAw1ZCv2F4dIANQe6+ytMEJgrEmk4fG/i+p47gebt1kIwMdUkIGh8MMTjIh0j0hUMD
XEzxVKeVSK31O24GifBRCPza9vy883bcAhCgewJSvVKxjko2OOpsZSges1/65zzd4G/aBq+JWQrT
3ft1/bLIR6TQAWnVerGssJdBzqeI/irw30V+TQ7qFM7+/DHJbXLdf3by6PYD0X/Egp4MdKnI6IZ9
9WdtbBPw4wsqxuGZMxIflcQWGSjSUFijUYPzHS5CTDYjCvtxCXBmcbpNzvmezbQqw3VKvAYyKs8I
sjWkIIrkth6QZSNV06Coc7G2DHWKkH1S6WIILV8NWifRzg23XKdcC3K0O5ppXlHBl08PvodCwudn
zI2HDDZ6Gapc5DemC6m6vuXzTztz2quAQKt9SsgHWKukxNjvYZ32YkhTCGjsOybaggIB3hVEqrdv
mC3jShgsGTp4PGucd0ljTR4TIB5FChDyqDeZt/UItTihM/ET+IoryEvq8mRh+g8hm3QZErKOwHiq
rtCkhXtpC9tN4xbyPa/Vws87BLpNszjCNVabxefTjukgQ39lZsAc8WC9gOktfiijqPs5OWf1g2t4
wgrirt5tNxtKFagJCQKH5oZzZES1r1R47VhjYUEvgY3SIhLddlBJqk2zzYVTtODDaaEJ0uivisWr
Jn6K+tVhCRwftYm6hMzxPcPFmbd9yzy4ldhDiQEjoNT79EWPKZ2p1VZzrXW+qOnCuCKiz6HghS7O
FG/NvAjVEvCe4tzIOnuDuKT1XMU2kJ5QUFk+219tEVzm0IXq1PVxuFsRdEfZf6OA8Baw2OMFF11D
DrM8e/39K+0oTL5x2d+pQ3lsroabJO+eDbEtnVk73mv3w4AyJb7+OxAJVt7wHsZ/c3PTloFWZlBl
5rEfnKSKT7CNexdVl12dsTTKv0RObmyU0FZLBP6d6hAgSsFVxiTJt0h8Uiw5/w+EqZ7YwJVWRZY+
3CxyFdl/FZRnW6hxIuCO8gX+6GgQ+/y16LmRG+QcH6M8JeAoMsR0Z57DT3rD1UcNfENZjusT/hHp
Ra/I+yL57X0tyYl/HhxuJ0KiNc5x8VM97VhS7OTStLimvVCh/DbUjZ6hHrMvBfoF6aCEbDX0biBD
rDihhsUe0v2ZrLMn2sF5sI/R+RUUmroTzDRedw1vYegsUQwmG6UlYqF0++CmLlmVYfwFcXczNxR3
HtrTHCEr6gQnQpvp4rJyy1XmjzZXOsvbccOvIAUm1gmt6GTkq5r2O0Q+Fq6Y/VagonH+TAEhkbMM
ttk7Q1wkFQUGX4dnpMhJcKab+vydIPWoMPobUwEljRg9sI88dr85BjYxBvuR/p8seP22OgfEbfj4
J2Z7ZUo7CXug/3FHtRsQtjI8G7mHYdUy5AQbLv+uY+VBlJRbzgNY0Ew6JCo/eB+Je41f2jS/QfuZ
Qve6yd6XDlvxi94dCyMj3mpVcbg/XB8061EvWBpweR16mFif1UtUBA8Un8rJ6FXBmt9DQshCiAMS
vZGwGTgaKsK0Vs7kAPJuSP1x4LSxq/RJ2lAHCl7Eo7ge3IjLOZMzO6xRw4kNHFtyunuJorhzCLTF
APeGquTIRnut/mkVJDfd3HMTNRMdjAJj82Z002jESmmvpHw4GGagmkTqsA89Wmxs0cNS7sHtP4wN
Iy/XSBICucBm50NzrkZtVsNWWLNdY6cFFOBKJyzMHNyGrAsgUI/UhCbzPGtPsKoBKZZAQ5Dm01Gh
sCiVJexYKrJWFQEd7GzGYv7hoDjuD0gy3YTNaKXjKbMynRSZynS/MXaMdz6P/1L8wHKNBbzR0iuT
jawUPn39QFjuDvPFh1cxrEvgC27NO5xNl7nApkSkPK4/Wmc0sKeIFSfWvZz3EOf/++/b/H2X3oiv
JlKXrLYVcTDrxcQRdsmQWwlNq12Vgawr7wg5sk/HAprbtIg6p5QpRRQsuJAZita2Vt548suj7TIL
YfEQ9/19va/iKuQdGs5oF+/KZ+RlzxjM8pI/Z+2ioIVRpPWEQ4WRa54cnQ+DuVy8dDggQEMQ9b1t
IkuQ35kiqask5ZYR1CMVJLhBeTHSLxnI2tUZPyUredRLBB/fswrTfU9rwr0S0GzxdtjJqBrgYEWF
RZGYicFcNvqXSwcVNz4gXcaxzjr3o7jNVsmt586Xtq2RYtxaqZ5KOGZ5pnk1br5gYFIlFUSEjQrO
KIUKdrtFErgeuX0gKm9v3oC12FvadYMZRFsZUAltb+mJURYPOscQQhbaumsAZ7OgLGM94f6LmMKc
X4YWVbn+EekfwCIT9eXOwnyiI55uS3cZeO23lDocYhNNNEIR4HiUTJvvTWq7eFBRFugG87HBISpU
fwlYJX3mH+a8/hSR6xIknLrf3jE8zm17hMOPUUzpKr2DgFoSMQ//CiOR7S8SrtPQQJ0d6iIbaxeF
qW9cjMoJzrIIlnjghDtHUel+fw1xqXeqCTOG3u7sYWb52jeo49NLg+Uqg6jshPd9xeeXryLb5bw5
48qVx2l6vn+ItFajtpEFeEugXrQ3rVSbqdIGDkdNnZSCWQt7ch8UjtFBDrKYSRF/W4huMHHth2Nv
HR1gT55UF/+qQN7wAZJH5jy06omB4bU8BVPao5Jx8Az7ZAsJb8PpQs0Dep3FoqaiCUDBuot8l52q
3BQTsbm2owU7pY2mPQpPDqZctTXjvpwiCuh29mqRspXvWgyVzKq8Ww33W839NSV61qqKROImnRLv
FC5uFhGxd5XblEqOSZFybu468k52CTJE+8si2tGveBPa6ZSguaBQfmFwt+7bAM1DjdsgGkTi20vi
3Uvjx5FIqHJaN/VFK4EmwSYCol2KLE52ujXWAPAhbAdIc5yp6HEswwGCi1rY37lx+NUDmUSMzvgc
MPTDbo9z/trBwEM6fQB14q2xCcvVdA2zQfc28YgDOihxmflr33z9QfxsOCxIIr2DsoNW1eblEtFY
eSoC9xUgitqkNrvbw+5Jg3oMMj9kfyqzlDpLVaiKUKLW0hsUcoB7AyWoqoS23zcbeTM40ESc5F+1
CpRsWnyxhNFUqdbhl1GXTpYU+CztuVoChMO7KdnKAhQC0uDcKSnkewym++kqAWQSer2ZJB7L2mb2
tg6AYgGtzfMmaUXq4NLJ0CRQR4lD5kwov0k3lYm9rjw9T6wgyl2rS7v3sKG0jA+AzObZVoMFvCZ8
pN0yaDtgxoi/rgzOjkWuo6JIHfLdHXStJg91qGj8tTIkN7AFbhpUn1KZGwClvqYCTuZ2/GgYbq41
PXripqoGh8gIw2gl6KtJ7zA/yeh/Dk7c8EBLk1vEnMJIg2epXGihIV2fRBr3C5O6MzallrV1rpqA
ZT4sosU7r96wnsz3WQnElM6MzyEAkYWBKhg+lkW1hZWXyFjAEODM8aK/RI5GEB+wVnpk8QfpI4n6
6v6hbEw4s6RuBghJzSv35L5zVUkW3rGmVJsBrEaa+6ZJx7F3GhHlGZ+CmOJduJzmUr4QcArCZhtR
ghqHQhxvctf2QzUjpD5R80+t51LkEWn2pAYaSuc0lQLZSzrfKwHUg3eeT7WaRad/B5xFeHW8Fhkt
VlSX3kiHKD90RcE3gy7KwQqXqZTdUBqn5BnA30/7VEucrqxuWQ7wUUokiR4PWqG2n3+VWTSWaLhh
mP2RlAsrPsdy3NtnqI1G2Spt9oiLoJhy/WlZllTu7zSNH1cxUsQVUMIsM3ENEqyn4h/9xCc6M9JL
WV1E7yEtnGIncTeT3feA5YSl71AE3a44ooiKSyP0nvgS0cYN6Kz+Nm4DyOXFV8d3Ki79FOSO7NC6
FiYNh4uxvvjQqPLn/r1JL9MKWF7rvgTE2WYof74ur3vJ2mXm3Ykj14ZhsiJ6N7eGlEHL5xkly78E
kQloLWNUGArNe018OKhoWXido2wDR3STG/DBVHSOcVGe6c1KcHvVyctDAy7jSPjBPdd0YQG/oMch
kMvAX+UFRorAu22rzWz7iwFLVNgz6M02rdOVlGXny0mTzP7SCeQAQHW1UsLa5nn6bB2ZChvWM9WM
g89nbTDGFpCxqpfiGgHNrSYsk6x4ZTYL2mYmFo9ZSApbf2jJ6IlErl1Uz/3J5KprATz6ZrNB97hN
KU2D15+GS+pZMKVBlzci4h+NVtLSFhSX4phA7C/y9if1qDcodwJHCVqDJLR29vb7wshPGZls1EB3
nXs0Jg1z10dcD+4KMjL8Q8OP2gVbwszMYqiO99IDjJl3dRSPe5v/BazQKprrfQxwBnQnQgL5A4hG
pCxH00vciV1MIrSMhdeBLJ3/PlowDCBtErmutsrjSY/3NAo82HdLrMZpmAkROpl2KMktanexZ1Jj
+m1kcGlN1yxvAI+1EibdM5omX0dGazHuNxth1jQNWOILRxMkuUvqtE/9C0v547Dhfiq8SyEQ5F9t
2moFGG6s2KTXTuedlv5gC0SoX+U4b2JN8LfhV7PihzNTlu58hfK+ZpGGFgQCl2n5F96bWrJDraWF
4vKsexBzDiYm2qMeOc/Cvr8uAS7r2XegDfltNYRDFWB4jzLmXjF6U4mcbKZQelx4oAljzg4HcuPq
SDwrGinhIWPfUcTi/cyU+Y8uevzBhu36Px52KutmTAyIDJ29Fzb5wMmEKm8STEbHPoalTcxlhpjg
qrnNfiSj9YYP2q0SsGHHD7RZAMk4YRqrUqZEOUfhVGqK+G56OpdHnzgj6jC2BNBkh9Vf0DjaHH/6
1yIvKeil0jiCB6eYLtGx6QGFaXgJHPoZMNtNHBdBVNo6fJJfd8mdlGCITQW6nDtW+2QOdy+yWpHl
I/1LwTTee8Jq3yLaYi2/uM5Y0iwUOzxRd3QxY/jA3udhH/brUTw0zMvt7IeFMFwYXJHhSU6qwqkJ
zl9lYqbaDPTskJm1MZMYYwirELehm2wTehZ3/3TP6NvXXyF9Px/ALQIrxeZWVC6rwS6S2nIa+C4q
GHKAauAAn8YBBU23784WAcayZJbu/0sqyqCEPrgXcxLJ7LsbD+0BHOsVBiLfA0LmNqa4OG8AKqv5
AwLo5KFqdenFbT7IBz4XrtL+xU/P10rikwzA0XJUNAvjT4yfOGDQG67Hk/cJIxDM5iPQm1ANnqki
5Zr+uqWr/QoN6R0MQyEubhIH3SGL3CPVtV1BSTq3AW4X7e4A3UuhpE78+0HC/QeQSjMyOZ10Vqft
cFXFOF64xV7I1C/EIGEqtep3t2HcDrWuuPj0hVgBZxDE/QEzzTX18IKQjQ5T3cdW9SgrFHQFE+Gz
4nKYQl4DtSZQ9ksOUzyBWTnQ6dWqxB4pUnjO0ojhPrRRT27F4DhJ06Dd1LJy7seS6ZDTnaGeksMc
GQwgPcH4bqHRqiBWP6KN9b5x50tZ7f+fo4ZdzUWtyAGKbpAssOY/Jck/6C/8bADVLFVw8ZnQAjTd
d5/A/ujR1EFkdUoNtJ6OXz3UBxMlANVJZmj0Du07X7dz0v46/OhLn58FHk2CTqjHJapdLJ7bHiG5
rjA1RPrD55Tq2ztdQWHyfYx6p0OVO3A6EOaYbwAdSLLrWzVu1VCocWVHuHcPFIIJC4tciZZenyli
fwRYL+LZWRbkzUcManVbpmPkJXpnYTidpSBv7v6UIqn8txlJDRWVXa5EfAnUPzkvJftgfon3W/e0
pAJr1jmwiHekoyu7G8tdEAn8d1sCyvVsl+jI7dwEQOXtPpGF7L6aJVCz/WNYbQXNLXbOyOaZZGue
vtvfXcCo8D5wQYuKfa6M2T/7pgjtf5pJ44LqD19XB8HTOL1beGuJWowF4FRy09S63syXauwYYJGS
tXNFdmdAQLb/7fc69EvKULmRQAhxW/HLSR3JvhiAWdNjzG7QWspqWuXCO/ydDzwiifV5KpeHdBsM
FZwJSMBkqk3Z0IBb/SCMm7GmpY/5RN9rXkqOf14QlMtLL+OWPfgDi8eEFH8Myq//Ngh2U9L30pgX
LCUnojHtUIRxSD1MUQyk3AGEF8XwYwxdnznmxPjplhj0IthtnlB3GCVENMnzaPr683wyDOKIqm5N
ETR2ZzH5KnE7U7a2cp/C1BUtg3LbX6ksZtWnfMNjqHAKlmBHDyb6slSHadRCwuDi6LAncgTbkcyA
0vr4B7ptbvSFi9j7YOKij4G48NnbP6qYYOma/SLqfwENeSx72TsrDJP+8W0FIj7eJc9eQAor6EGM
YCHQElIxbpd5ks3LBrGQ7Oj3MnkzKYJwwQcBIEU3AReIvKPUjAM5S9cbLzYz9A+rbWr2BXC+qD0D
XclS/YfKgxLB73a+rYXRHzdMevJ4+xdPo2b4Pp15Lyj7h3NKvd7TWx8CTGBg9hlvZsISKudi86Ax
KkEgy0BcwG5kPib6LtlAJNfCgsx2HMRxgaNTgF2xNvpfWfSVfSVbZKm/TBOUlYMaVUEUJkcxCEea
xdchLAGc68uFV56Qykgt6xDZeT2MUoxNPXyOPcESCu69nElrtpJ0bneFVkkqZ1ddP9ZJSOq5jfc3
ArtzeXNwCSITfLoSTEeXV8h1xcOWoiuv+DY2nnfhyp5b+35IRRLRLSNfGyLZTejDmvsqYqcIxrKk
P4PrsCHquziYhkSH7PQaY6hdTqVYfde/gbtpQByElV6SOuxNypjQ9FCVJxvjRryq3WsfVq93niND
1CBDtW5NR6xHHLg4T66c2BVnvnr+Dun5ag5HYof8SeYOwD2fw6qCvJmM5OShwrys3pTBCFloFxff
gZ64E2KuL7bpb/4FCOH2sFeugh2uFCHJMBk80D4Ff0io60gGb+D2feRgJbO3OPyYc/TWzQxIb//s
9nnXGPcE8soV7ISz1wpBWCpBigVWf71luZ8thj1M1gRICbotlaMgqszVyW1GzzHqwJCEuGGv1CS7
Llk9/tpkBej9MG5VG0sTvj9WW10jpwubwKITGTzS600xRsdy1V6ELSxMm03rjdaFGg/D2c/kCaZa
N6jpExg/ZXcm5eeEQOpocm1P3vWqVSP9x8zTNt2fQKEDco/bhL5SFmf5DWYnJ9szGTktBeI7OmeI
Dwu0KIJpj6IJb0cBEoOSQeuA+YvVvPX1OA8orP/u7cT38BPf31gdQ9KXRBypdDSN6eGQIw/P9W6K
zed8kfJ+mPPU/7TmEC4RuY+0Q90XxnjaJRC31pyoFLIA7eqXxLYPoz21XY8xgih9poLBICN3KskS
IyxK/OKibfzl6g1KiLygg9E0BD+FTo3rZ4Yj6sQiGTYA9fL0J4BWce4B072nPxTlUHefEGxg+F29
fkYP18whWujOfQGMnoAQ+IPXjNMCxu4mOEGjW0iAt3G5r9J5w9RUQBU/cAr7TaJR0AqyNgRG9P/p
2bcEH33kC3IDPUUOeb0dnQKKdApTbJEV51jIEwJwhGm5JRIjjD/UOm1MFBcnUtnC66c1juYgJTuu
9cTLDKyKpwss+37oAZUP+KWOAPGV9RiAH39QtUXiY7Q+Kzt5kgLh0byblX33T+1aGJoZ+C267P87
bPWZPB6+5zVFroS2qjy1jLBndpm90sU6Tac5PAliZkO/lUYrjZ3qbiDFdoas8zlxzdwgNNB0TNb7
x5QrSUJrcu7eWv6mg//kcDXpf5/7kxfVhje/WN7ZXwtUttkB4yGJ7/h/IRWAQxuPo3X45HGD+cfg
wPw615Ow4shBYkslHKdw9wLzg39HsmiPtnatX13BjbFt1cgG740r+fGVAMqJ58qTSTfIp+S+q8Ce
bBORiRXYsn7gvReN/bGTR3NOmByfpM54Q6oSGxmO1tkPi4z3XDa4460LTsqxfJLR7HKJTbAbr7mZ
KVn4ojsK9265izMK4ykXqR4PZ2fMTcNUoQnvxxXCZPeEEB13mvTuwDqXl4FwElcQcvEr7CQMD82A
Yt39hIZVkVzO/lJCdjJqpfBoJqn6mzu2Ps/xloMSkbH0Q5K7SxVE0K+uBtmAUKfd9xW4S6pxUiA2
6XDSNrkYvHmJ0l8duOEtQzIIXADXlbO/Aq/kyjzFS5I8x8oRd2jr7uWY9v08gAfoYgYHL5L7DNqY
NQYkn/6xBZxI7GvyGaHu/5VwUXBsRL01iPs38S+lzZV99vcwSM8cqbyrURVE2wMKkin+8/lYDY3q
TiF51ogYkzU6eSsudKmyO/1UBhje5G7alFFELqNqkDDVtzPfBsYnk5H34Oylunn2EopX/I1euOfP
RY1hpiX3O5/wA+bGZsrh84h19I4QD+YWVWMx2xprjyNS61H+3Bbubev+CksbEN+uEC8OZbYtCEpL
hFxHXNVVDzV8GLnoEE8KWuEY5xzaM8YXV8Jg46yRVwJlTBOUxmOXu4HQ4LTBz3rJwmtuqrA2HcS3
J9V08kVIDeaUYClKmlSi5yvoS0rxBBQj67CZTAhWhnLvLxK5m5wLzav/Lyteum2CWXvU1pzzDiA5
0W48v7lc2IVG0CWyxNXNc3z6TRkfMi0S6DcNYwsNOISDB+smI4Ibtuu7Ifsg/yvqXvpX38o7X1P4
MxC0oPPOxwml9ngYctAxgNtCgNFaDY1WwzQRMlwemCKsoU+K7obH3EGt1Q1Jsxb5wMLTy9ozNjqs
YhnIirayCxaMHG9RjSzY/Thzpljh0y/TWETZsbZrBO/k7HBH7NCriEXNolajEIdTCWP5dLsqLO4b
Kc5r4qrkB1kdcrYVVs3aEG/RcjykkEI63foHECtd9pYUmK8h5oHkGq53QIVVgDSEjjCv7Vrjm4gq
dvhxIrpuQOf8yJzNKxtAwGANWArjz8IcKNoAMGmHuiR/qcoBT5Lu/8rEaIqgGYIPwtW336Jb2g3p
VZf2KYKb1IIcbtUsV9qZ/LHpOuhaSjlb/m0+vEklKPZx1fU7qgq6nnNOm6j9rV5Uy/1vhmzYH/IF
Vnla4ikcvmZBUtRklsNOaWIyO3wbcZQo5TjYoF+Uk6YSKRw3jX0MOT4JDf2+6VmUsne1q3lW+Lrj
Q+3Iy3Ie+nOu3NMzxGB0noViu1j2AuT7t6Rnir74c7X6L7Epu16AwR+bY1n1VfWdeupES2M0b78P
njj43nh0aezMlIr6CSXMwgDL+sl1CdxAOibExU6L9SCQgJedxzB0uz3ZyFfx5izp487k4vYOSS3w
mzy2w48By0RxrvTg+MQMrrCxA66ie8JeY8iZenvLr1KgAL/nlrT+og/DVQ2UqQM9QP8Ck+ksL9Rc
1WtYEH6Q1UaKPxlx+J10DvAkIVkC2WMUWBhixbGwETufqSs1s6OAfYwBOgZqLuoPnxKcB1dEz2x9
7S1b8uxjQirB+4GoAU5QRlcHQ2B4rrAOemnE4TAE26ZbTmcvkYpnQobG/NDEPpjXsxqXspTQnV9J
Lpy6XDZkWdcMZeZ9tbyHvZafDgYPmBwCJyHOUNrNWXmKQvQFslzE85ZXrwveim9Byq8aa0Trz9O3
cTutZHqQtV3zD85g9MAt7VTkyzKg4PpZxx4loFRjErdSvdH+KL6cdmZBzj9hm4geEK+OLiPwSTBp
2nexEZeLwFrTSXKre6BGvZ8HpkW/3lRd7Z/NfWc34Zo4iFFem934ZxVpUocfhi03KBuqd0EY4nX9
1GnDGj3NwvZBDjuaPo5e5oPiZKFb82rkp5zMgQdkrQxOEKBTmoyU9Jqs26Cd5hWRQCa4Pnmodzph
cXqCXC6ybzRy2mTCjywSlCjgTsfy0soziExXcOXgRdNpuD9Rk3KfN7I5NxPpnk6OLpDSTMD9we4E
ecVFjkXI/8BKVbJ9OK52WHc6GT0s4Cggirthd28HIlUsNrXmt21GpyfzlE5/QBIf9D66aiMXaIjW
TMYVkzs2dIxLY+YrqSbF1KhJ1kmfy0bf2MD+1Y2SWsyp4QUC3wKExEw+Vf78N1Zp+RIHiJknvaiW
giGaQzwO/WOgWYkeK1nWE4qVhtTDRwm2ABbzycjUq0Urt4frwR9ki06sQtSjqEfd6nwnmjmmtWfH
RIXqj3gh29mj46d5wBTs8PBu+mvqfDmBL5ekwJHRCdIZWnc0B5lGn7H4WgM5ev6AGcNx6xwW919u
TK2MjbBIMOCOAJ6kPAlB97aDT9iVMD8r42bzpNqcchHf88/VFUEW+rbrsZBDnxyqQyYM3dIb8WpW
5Yfcz30ar4HgNRwbp/HcbFIPS4lYDexbd6aFJrGYE2xDtnwmwCeRaenYhd3MK9iY+1DkYoRXyl0j
uWpMgNqhZICQ1lmZyMTiqERWi6XEguANHGjilvHO6YQ9EckweZuWP7orpZLYIPvBfnkJSYOr3XLj
z2FXe7vaOO/S8+9RvGuitaSugM3eNBKpjWLVI8L/afiqIcuydhzfFPYe6LOmON4g4NVZfZb2SGZT
IgsAnF595QdQo2Y4cgqQtv1NyQBip+oVoDUmikOzH8nRRDjVEOGkx4YzDnM6YTcCx6wlyNkUsXNx
CbV86wBfeZ9y5/r9iYC9RUy6BtR4/xk7ms1NKCRC6ykS2u5Yvrq8yv18URQwEmQCMVntwQrGlpqI
xFpDnPx5pGebvjadDyqj6zI4TsVBX1wjIS6tl1ix2qIcBwZ4hXTJpsVM+fHHzxdaqwGjJT3xyL9D
WEQeCHCVTdHYqGtYwyyZzOE+cufOQddqzFUVOMwnFGjSF6eEm23G/5LVx2dKc5RuASr5ZrhtK5rT
oT5eKAU2yQ8YM4xg3wDRgehELGZnhKnFbO96Oe577pso9otOawGbSQpDlV3uPvRipq2+BEt00O6W
yxYwaBvu1p9r4xeBsJDtTEv9cUy9bbLhG9VceuYjSX+THRcIVyCmOqxyJLbOIgRO5jaTR0GAih/G
zeZoofeJIvkzSFhG+c+eaffQI2tz3exFvC4mjsRuYjnaGF8os6ozN20SwI/oCJYwBZ/XSqD2+8D7
PjLt9Res9FMbcSjUQRRC8RF8/q+qdL6m8zd51QetPz5Juf2UHxjm1wFUh+JeyBSWd5u/mm7Wfe6/
9FeRjeL75Q5SPsBPcpNjk8PRG8HZojPMDeAglL72O4e/90gH9V9uOawICWKbNM92YJbwhlNHr1ex
+h7FbsaydpxfcVlIEJ1q+BBmM6D5S0Bbq1msu+1og9Ll0DrDmu/5Wx/jee6GrVbvbOVpH2oXffmc
w61epywFJm9AhFbR0XDF1DJ++YYObF6tw/pkaViifm7gbY/fXhZLJe+9ECpvR2m+dZxY8qEIMwJq
p8a7t/PCu+TapHYFQYRkuqYa5Ft88aBfWca429uTHCxY7nj55AbAV3rlwFUhePm1Uco59v3i7ruY
5vc1ZDf/W9ubH8DkVuQ6Jd9mmPiy7pbGNtMrLeFQRMKg16YtmJtpCS9nq0m1qz+2dbOgZMzyU/5b
tNi2sCsbwzaOYUPV/+u7Dyg7Udy3LX6U7QVqoZ+eXGP6ngu3LRDNjD72WWpRMjaoAKvFzqJig8d2
47MMcd7m1AeOFvV3a3YLmekL1TA0YkAlsAMvlAED+Ze8B6+Xwhd5UJUrKeOPLvK+Nm4g2E4nEiGq
mn41PALF49dnFcgS9xkhbHK0aRvaWI/P9+YpsW3K+nlhKc4oigVogKg/kL6+BmXQRumgpNuW9BHd
OADqWQHTM4SaE4BbQEtzBufTGdsKdLPToAejZDSmEFndxq+8+DZiZZlnIrrejKbQiWuLUu40rDM6
t1ZHjZWsw1/omsMapCjRBokbP+ioK6t2TIpBHfrWZbRoaMxMPyIQfCWGfLiW4raVqjgOCL9L4jNb
oJwvW3lAuDjSu4E38eCMbF23o/8MeF0nelRAbvBZNt2iqK4Tv+QGmunrpx3Bd1yKNmIP4rnQuAqp
YGbj+snnFVA6WsZvDYA7vrVhhLvNDA0WtiSWXBUFiVUXRfqQb0tVkxfVnUC7GdWX64Ryp2CCcqIV
u02TL+iSF0yyVXl2mMz6jlxjLd7tO+2vC+ZTaf5jDx9/wPkdyVZRimml8JI6Fi7sVxJPcSL3OZF0
HKlSKSShE1bF9C1tWSPsOOgawG3CoELDOaJYagRdb3ZVL+ihUMU+yk4Z0G1xB9xOKT1wzOw5dNgL
7KOAAR9rhYWmkf4fgQq5TICzM0huHL/VMEg9ElsNBumBAyg4h5AhoxUORLTbreybHsZpz2USWAb+
nAY1Lw2bIHKDwDwQMeTEvxM9kQfxUHljNtyqXbGobuUct/94JzTF4rkVSUYKYZ4bUm7Xf65J/cGK
WDAqlOnF9nN11pECkVVzIWNxK9cyJSVD+YBExGO1PhhB+Bx0+BfD9gaXYDgkUrYczDqFQBR5otZC
dl8Ohww7tOqyEYGdkKfc+dPjaCAXZlWM/efGIL7oUWtJPTQgAAK+5vgGTL1UaHCqylL6DBdOdhuC
U/WLnYhmiQHPKXpcR4C6ezj/MtF/8NTCuuztx+nY0GgD5mapmfZsvWNjHfP3L5VQlKdQ+QmGtgx2
IkUpiuk6LGfdmAcfGAS3nvENgSZB9gHL5F5809QkKF/H4YhCiLLdYfL8fZRA+LHbbOfK5OTDx/Sr
RrxM0Bvtyb3ybqIa0qq7b6/mLYfb6cU1zBwntiBtLIgFRJhcmG8NCkqiTK2qQtGuJRgXnDwer7nt
9ZrVxAvGfEcIOlhwIQTWzPyDqyJp5Ny0PdKga7/rHDvJJWWOUEqZoj47HdCsxX8KAKCtuOITbVbn
Ed+BFZDX4WNfL4mYmITvPry9aUdyAUbJdFydrwqLelVBzKyi3+HSj5xT3q5u61rFc/cLmHNIvzx6
r4MZm9YLuToVQ9nh9nK+VIEbaH2o5XHxXu/LUB1IKHOm0mDJyus76qUlECkvep2OzYlmbWYhtIFC
K1+tGhTeT2/VfHroWtSJ7ulcE0k/ODNasHk8HIjzcA2n1tjNA6jtadcjP8HiHCy9x7YzzrSvzuIl
HrbwbOBox+ojxjgAUi/83+xkonpYeRV+Nl+CE2quJIlJzOZp12ButouwjmTN8D2FRRn/cGVgLGu+
8JzDRcGO9EQBxmuITDrW52NUJWHot1SQQl3Qxtj0e6M8OockMztexCasWLQ8NSs7pwcUXHUC1Hi4
6B3c5yc5zwR33coNo9HCd0UVzulNLB6pbDexOos7HwZp9DXlBLOJRTqG3oh5QMd+XuE/hn0b6lEq
9UnuP2XHL5wl/DqBLh5SAW+4lmimtfPJ2FGXfgc7iO76NwqRLt1OK20gFXXXjFo4iEJQo6O0rVOz
lRPybZZtFcLzVl0x7fzD2FMVX69W3Fg4t4Z17cU6YhIZZylbX7w7kq8F0lo/Yv2OkBTXs1OCDSIg
BmSZXXz2xAS0BA05SMaq9EzcSMqUcnchIwBlhvsts6yLfkR6qp59U8Im+hHV+fpMuPCORbdeqAkS
fk3xYXjo8ezjgO3iB4M8DM9ykm4JOWewxrEeomyKahEYe+G1AMKcpmbTKLTEr4bN48QWChss+Giq
OiMb4kmBSIseuKYMzxZ3G0Dv0N6qZ7t3uCvdU2Ios0qimp7S85hF7XDH7jmf9mBtkjAltQxPRTt/
hY0/WMmpB1SIcJ6CdpIH+E4tIpGyJfZl8N79U9x6eoppcWaMKlquDteeOFSqlGpIL54PqNNZyb80
sKx7uUP7vQLn2Arm22j4RVTfuSIGKC6KBHojpK+jBCLrp5D+JuGfKv4fpIDAgprc653IjqXgQuax
HfxIX7FIh+bh0zOF4ItS5szmjqxxK6aAq/w4tHp6OjCwP29dfGSRnYSPyb52T76PKGZhGjpTD3de
N3vmUlYmZ+Jzu335UmNvsyl6AYwjYMd+llavUoi+qLBl+hIQsKPHV3Yuq1FuP+g4uCt0+M3U3W9d
+BElibzCtcFLAQErAnHF8EwmjcVosnTnvRvEzrPQgUAw2Q5GI9ZvICaDeNqLd5sK+JcMPZjs3LZ2
oQTeMQbQ6MTNo9sFHhI8ZQDJBa6QhHEjoyJiQw8/bcR3tzouACizveIWoQp1sxUp1YcQYNqbajsn
+FqK0S6hFJqc29HgmfwANphZXRQ6taH0iM24ixcSHAo6nERXVqPRkgSOWQWK9Ic78TuDTqBz396s
CyFIPO6oZEs8dIawyLAJeQjK47/heT6MhOTn2Mo/a/gUr8eXFFnEVR5PdMadjSVEr177wdbzlTSV
FBEOo22lWkewzcF2iUe10UsN3ejXIlkpC/3gz+CSaKeua4TW7M92ryN8DEC/qLOrsTjBI+5BLd4h
lPnxKu38LvrxJKWp6cCwsZbTSB7WIbaSm9v397gUbDoChWMlQMQhOSQs11Nqxr4JiBMGBCoEA7Rf
LmUKI8th1AnPKpgwrp4DhokAnMqXKBnmRtFZz0UmeiMrxnmXxarv7OCIePl09bajMH2Ol1GO2i++
Nn62ojlcglIlpyXs3bMtll9F7i4pbIzchwtL0OMAVBd3bKEiHuYhPWWbN3PT9sReUczs8pOuk8TO
V6KwZg0E3zZftWnr7zV9iOZx6g5Ck72QRgG9lloKD0NjnsNvATMaA93TjgOGlkXi16zeD6yWuAmo
xDQdjkl41lh8gsTSuqBY5Et7u3yxmJGApP5+GRe8C2ESdpECNZBWn5HHUUoxiZ7sqK05O3NxVfgj
cnIvzVrC97te14FuxxZQfswrAsVLmX0fyK3zj7SfYOHGxyI+AcclOuVfuMVv59wNeI10tMdXslrM
t76fxjZPnQWhtvYKKNHxD1VBFRPLcxLIo9dYkQV4wgc9H3kArQxwOzUWT8cOxRkE5hvPCFZ03v7y
C+F1sxiaEdqHIQPuDsKiRiK8o0nhfK0OH/dMDjITqbTl4aAbabNxhDWYG9ONOy9z+T3pEpdHPs1A
iMPyoJ1n3L7vCMIahZwkuAvAyqysEiq8lz52xbiEyQUXSp3wwzDIo27xEnlnJxvIlE3L/kYPYSid
NstYFWqK5HySXtXNTwTXz3oG0mfn64rp84y3nZN7OE+gHKruzwhSz2H+SguxBfLeb2k/Z87YG/Uy
x3QfNALwGInXxiQYuylusWyQlRByZ37VSCIkTLGoQGeIRqU9m0UPjATtvhwqWyLJ6WCZv0+k+15Q
gknzmp6x3hCAE8PWEiXdvHXwJSvU7oiIMOe19jvpMnMZKXrke8PXVsjO6FgdN3T5NLWeW0rnwsRm
ESLXHjwrsD4Nt/x7peyantIbR6F2Se80zWZbMJp75LRMTXzEMmp5U3sPXrI3QV+++nJC+ecXYEwP
A54mZ+Vx089j4g0If0FZ5YWWDaFL5ULEBOA4l8lOmL3bDv9nocsprTwLUwS4++G4r99AgjgytfQT
O1xvg1AVyqh5i3HvE75KCpS//nZOoebFISBRhL7fDEm+TRa6/5CB38E6Hx80QO7WvjIs2BUXpHB3
EzVDRtGN9bKkbFTmHFrv8JJGnWU6SSKd8Lx1lYg+zysgiiEvRBbTzvYAPCZr+iILtLT7b9AEMq/E
/RUZaIbyote2T5YZF/6n0l9FfSkgQazG/4gkyfLPYs6bXsyJSjlk+r/XwLOpuuz50x3BJwzuoZ1N
fpykErcVOpKcMn2ygZPSgKg5AddXRp3CzGaT7ySrcrivdHskmOKVX8okZxy+AWfC0Aa6/4wzfnV7
NKBdRMkNf/hldb5m64yGNYkN2+BB6sMdQD+NqFFqywujWXHx9gq3eJuq9Xa9F+BTaNfBygOCkiHo
ZwWBpeqgaaE6yDjHvYi/SnWScE8oeEmvx1cHKUypQfstlxRWBbvN+MsCSJ8woOZU6H/OHYVzGvuh
GrvaE9juMizEavm+nAvkNtZB/XdX9YHJH6566KJGWg+7/2VzA05PMynE9zlZKm0+BCzeNzmfvW4m
+P148VzPM0iCY/YpeTENQmZhmJVS0jgU5F4OeXHe/kQaDvkFazcbl88AF4O6btJT1Ja9BSxOwyAh
j6N+Ma8hJKXonTb8NmGdrpWHBfs/ftbZbJRLqh+vuJOE1ox8pnWoIEl4rBwQ5QF4RB03F7TqgNGd
vFxJNP2F60NxpVBrsVwJvJZ8VnYhV9el1Z8kf1U20K9gYpR2aZ7V8JnAYs5oa98jv/uarKrGO9kb
9kEryuO6ecyXmpCK/mQRA72Z1NYTIMjcNEbLjdmS0Si3ZN46g30BNVfkEk9dLqo6X1dyncl7oHeq
7KKQSvnTK3EmvDWvSzewGk9Y1LVIe8KMSeV1Xl2y6y8HvXwDz8v+jp9uOdeO8kztOxEjMkgpxRJm
0AiWghB8kWW0fKB4ZCEB6daVwKUY2gTnlaM/tCd5J+hlkPofznf0m1BSF1mwin/t/G5o97rej01f
GbIkboVRVYthamzvuh9fFyQpSDpbntaQFurnEiRPoGDmDS/4v3mu+klYR+kHU91y+5oQwg7ZRPm3
6QpBhZaCA2bi/7sTy38/01A4PQUEu1GHNGd/VLCi6ujYhX3IEm00Atcv9cR5yMLI2qVgWlII0Yh4
CHrTULtzSNtIAgmVYUR/NXz1gN73XandGkupXMO9RaNetmO+9AJwFaw35Y4Qn4CPiKe0D88Z37yd
dVMvx++ElQ8zbdv+bzhRb/4tJp4Tkq5P2XFNvwSNxkuj2IX2PQ5DJBaSPqcqm9yqoNoNOgXE0fKd
0eop3qURtVy71O3vwSGGWWnTyfoa+UeRsXO8UQkybntiMTdFxrzS8tgDuU7Ui/62ZfODXeRJWYhS
HZcpdsl1Q6L6RWiVBTfOcLakb7N9KtecbD7K/U59XYr1YNhu1f0toclf3wdPcIDXD4o7mkfNFxhc
H1ICfqc0SCl1NV8Zrvuq+cpLnaSuFLuj48K1tBS6r1qjcfGOkkkfBPTndpFNGb4rU6mXe3fM7aG0
18js9mhylNZcXz8rjxZKz1onuWomZs7yr4bukLtcSfUdt16e8oegB+knK9yk0RdSNGXpc41OHaGm
JDu+2vTf8YJht9lkm1f0/3NtgtkafZTKrn4ZyLNOkbnMK8tKeHUaGi99IuYEUnO0xPDMAE0d6Oyq
roflqVf2/7wIWhD45ik6B4YqjDwX+c3zGj9dUah1H0enNIDrw7jDMg5OTU2LGef6IZljOdaX5ns9
rD7PKxw93gg18BFPt7H+p/gjZdf7CqH7Wq9N6626CYB8NNYgo4Od/1A2EDXt+UzJ82hayIgtpmu3
CXBXs9XEFnunvG25sWeOgKYw8TuOitpBz92iRixmoKfyhw76pdNVDEgJS8NfCP/z51NkPVZrdU4f
tIVGPPW52New2wKj/sQ3+HBqvy9Z6bkTxcK1Eqh0gg812rJd08cGm8oyX9STk34F2fFNEBn9VIDa
JEK+B5wm5lDhERDh4toeXCF4ZmRdK9VJx6oe9/1gYAM9dcikYni//bcvQLxT34UImHang87IRl83
BJ/Eqy1pDxu0U1psAWJ2ehg8qPTVvnElqtgKIdgG3Ot+SsYAFQi3i31NcVFUpV0NBiMaCqyGZ3FB
ImFzZC1lsCHnOcOjUtltGgWm73CrSPEQ2BtwK4E0MqkBfnA+xyTTJs/dp17L7UDjTOHju8e0wyHb
ahnJFq2CcKnzkot6crcN+26NMZUvhaCw5hfwTxHwwLVwJhsgvssquyzOTYDIC/AlHBN4hpt+rF3M
d7pU2LlHQ1M5yl6AW50JFRiZKmhzQVTL+xX1PZJFEyhyzT9Mon0PbpqCFCXr8oNAZwFQguX9ruoF
BbVx2wMC1O2wuyQQNsMXrqLWndB4tweeoADzs+NRXSyFqyBF56SoY3VfR4a4aAdValLH2f7Y3GL5
3LNf8z9HqK8Fv+ufxAp/8m5uHtJfx2FmFcAqhzUW7aU2DdZ8DUUw7ueqL1BGoWi2RWadJcvzKmi7
x2r6+W4r/cZ7u8XFYQeyCU9re5jwM240Q1svG2Lcgckr69b/Aqfgn6mSeFwECVSDL0dOlnOvi6j6
QxXmcvxXd9XyWbr1BVYdJZtxsX3bkkUlx7Hhcc71VRaXD2TU0TCf9P5fFGhRqs5qCwcr2UFRtexq
0ew/v3j4x40gwKZ6tPDtqiR8Ednz4I2uCOGzASv/18ttnZHUvtvVVB7dFQl21a8WpeITqAliQDBt
+qWi7UHzF0QRa/nQN3ta+hSGWTiRaJ4O+dVa64mgrJnqpe/8JGgQQWgA6tsUtBrS0YJssOl6IfW9
wqn/Q6SqbNOKv1nho182I8SYoWZg7Q2LS/O0XHSQY4DFcYCaOFHABPWxcVlppMPyYki4QYWKdLZa
mzaOliixjIrulr1toyaju9TygQTAy5GA90HOAek8tSYRWd6baMGFWg9GsIEtvGQlEO4G6p1g6MX8
y6hrKrVRfHAkiD3j8Ob7tRD+qsh2/mYrE5O013wJ+QWO3GmdEGm6KCUq0LU/9GQ4xt8i3BsYGPcE
7IB7IZ7oqvGWIQlM7EUDQ7C1/FJWenNo0nDJhm8tqowbvxPHlcCeOnt1l1O0AoRaioZ7Zyeh6S3c
bI7ZDroOROY/2Jce1KWA0NPhv+dXqYWu+gDbNQuD2Cjz2eIp6ux9xS97zAm5P9l9CZVNM4p/RAOa
fJg4uYyhSelYxao2wqodywidz3E0rAq8Q0FEOA7wtHo6kfwY9CqpprFWeOgdXkoWsUhOqE1Gqof9
NKA4eAUmvUcVPxVqgSwuAKokaO2ucNTQV1sT/pe9/39Wv2vPkPuUtv7h27GRM7b6dMgVmFhv/C1o
2Z7+M+Bw0AENNXDm+e4cwcUnM0mz4ddjQoWUxgCDStngf6nbWxRupE4AdX4ID6m8K9RqJLZAQrgn
NjDw39emMpMWxHZXfyKLPQVL0VQJAC4GCr3+cb2NL9Nby7KE2iDaDwbgzdFBMBXaWRt/8Ihd+aOp
0xOwVfrjeewufgLLVqnolcvSNYaG9iL2nqOdT9aa4ZUcNRD6m5ZRSKsaCaep7Jic8toA9am/EbkR
AXghP9FV7+xkwyDzsiUF3uVKn/CEIpqRqovsOtYA2ss4I0oDVfh/UtIvuMcDt1Y4MVBFbK2xr+i3
XJuvJnMglmEgp4UVzZOc+izj5X/f0MZZvTvrf5q+wVcBrA3/Itg9H7tKMERSIA3uU9+865kvPYaX
x3dDJ2J/ns/P6qV8aL7ZWixg0NM2D5ORtnSAEKI5BibbPNEkc2sq672Jr8YnPpgQajnrCyLbCkxZ
Lfv0CAplBRLi6CB1JhIXJ8dmY8EAi2LTzQqSi6wEhBZwkl7nngwNMwe6p9ETsg2k6k3iBykcOH0S
17r3V/WhpDx+0GEajuq3GtZ0JFLy434XgdFIhxdcom6dyE8REgB8Ce33MM8p+0UkEssz9D7+PRVR
p36EUoC6pRvuvc8wJC9w+A9Svp+hSKugWKNIZzw52pnCloFMFOJxOfTB6zo3cT2UiEZLYRGSKoIR
wi3CiSN7TwtOLueS0pf9EPVpFwytB6p4NqOyxoHk4Yn6r6vyxbukNlBCQUOk7CDd8RApGfkmNhUh
e14FrUQgTsEKOGbDqQTIp/TCzUXKnSdNrf6BgTV7iOYSBPyGOZ8+ayqyvf+DwfdHu5lyj76bCSKo
hhgJE27tlN32xHpibye4gpPpbm0oYuAPCujzxYqI0GfyDaF9G090jwQUjoRBYoO49YwG31uBFxCU
fZi9SfNVR4/MvSaZdkjFKX/YGnS2WMHrVweazU4OLeN6iWS/aFbw/gzoolNd/UA+uLj2iQU+ASdx
7GYaoCyl+VOkTzDu1mfXpxqJfFi0ZexQVlztr6Ky+Of2Z1gYyQixSB88KK28Z3hy71XXcg+zjG7r
gbHN8dZMNx1V2m9mckb+q5ORm7ygEUKI5vNv/oIpyIG1FsHDjuO7qYuafBaaLBtfSaX/R0UitbTN
C1YK7optvw3m++Dwi/ASrYf6csyQ7h8R57fkBj+EFZUNxf6fEaGJofN/R/ptUW3q7q4hNtyulWba
omdoBcdmcqr9p+wVytqa4hpg3x4FyKur21yZmP9LiYjpeCL26FZ0r6ky6JCO77sGASeiqQj002O2
/zSJJbUBLKxangBbFypXD0X+oDWqWI4vgMsipR1HLb/mYxHKcM8ht1RIR+4iSHRHWBLV3zpFB4FM
E98JjAmbTDJJoGhAXE8KM1nrKwxNxDEBqBeXHKaIZYRbOAybXvw9NJVt7UM/42waKMQT8laxr2z/
NzUi1gGJaOT7BGZWyx+f/FC7pDO2V2tHbJsHlfiKkEWv1Yes758YMpyHH0iRpRHE6q3i2monv34W
iPN4ZEmA9pk3S55tm+A7yGCEPq2FTMqs31U9jGymwXgW5tyAxdU1+Z9z+yA2xPAg/kroSyPjBZU7
/LQ/aFjwfT02+V64QoBoaubVx1nhrcMmkqx8T3jJJHS/Fk0bdOWTQ9RDvJ/2B1wuIxGLIDu6+Axl
0VIPruQNb4XdEAYV2qjvFRjfNuYIt2FQK3MBq8TssYdS/h7CzDU1loOirFxhmgig8y0bXl1sVI6S
B9bhKBLPry5whPmAcjiicBQ4pvr1eK1vylSk7zN3wGVg9t8PDprQ6KvA0MmfQdToeAldyY+54VTk
hu8iK7qizEH7IkPluP75iJ0mQ0wxdpqlzJR8wFyRTzUFHHIo380kE04kT/PpEeiuUNZBMB8bW3oA
RDYqvySOh36JPLk5/TiJ2Ts0KUuf9DW8Gb/4RqmAyMal2c00adiz+WoCnDoOa1l0wr1ej/5ValX6
DfGAK7ZF6p8nqNhNI/8M2McW3HHXyTZ5mZSQZDabeaSm2dqXP2o4vQU+Q4KtDK8wLQB2Eq3eV5Qb
/JyQgCXsgCHiZoavouD0YCg9ZiNRWgG1Qa61V0+R75qNCfruT1OcNuAdKfXyZkM9ZUu8zL2hdGlL
cxI92WMdGub2lN1gIxikljXZMU7ZUEfung8JZN2gml2zcAPd7myUWPZRmH+lMcsnKSU+UBjRh6r6
TyiUCe7GXtKASueAQFNhcfhkL2Oi/Jocmea9UStL8tPonbRvFzamtXu750c6UcGiiam+Y+iDY/wf
sHl5tQL/OJkiFekH1PQnAZp+96EZFwkhCucpYBiGeLM2KaQMcvs93z2DhbCcEz7igrg5fZsR1/En
bVA5xJiDeH1hXfO0O6Uck4jG5mAZrtur0O41TZu58aDPOBjdUVZJ2Ruq5QUQF0FxGtR4NMo01B+q
NBuvlOjN9PqV3nJHylTlVVskgOtvL4tC9uN6YIBjlUFfiTSJ6lDA+Jm2oJIVClMaIulXSit4utvK
b9t5yjHgh+O6fSM/Y+M6SBBaN3o+Iku3GPd2dLLAVBftsVT/m27Iy8/nej4N3IglU+gXN6n2sPoP
sMLy2ZkYU/AR+1kPVo9kfI1Mb9kzWN1+ZB2+fiBJtBISzeMIgZJUPkxtS0ejHr1io9no8UqN8QNq
cfQ4M27jiVxWLPufxbGWsN3UKts24v2eJZg9PPEWvawDubMnm//69NCgcx/iUqJs30sbNsHB2sjN
v/d9U0OBKDXW7hDMfZSHjgnUGZHMMSg8dS+FeKDvrLib6Cv+mLwsOLXW2vksapPb+TKX1GzSM6vU
PMfSwwoQpFS6XpQEI8w5sFy3rr1LTPW9NMaHfvG2te7YmhLvwFYmt6dbH3aTXX9M4Zs2Ulq44BGC
TLwGjhwJxTPXOvySGGNXJ0NEebUHTzhp9h3HpzpIlde/f7RlFpqq1GZz/2kN/L/wj3MJ7la8z+nD
8ri1nFNxqvn9cYIWKcimfLziB0V1e36t1yfN9oeoftyeaI7z42AHPpMOITRZ19AfrRxkoARpHuwU
j2kYQaMWzYIyZIWvU1UMcLqc8aTNjE/+JcxlS454W7Np+Aacy8W/gDqOJYknEm5e5sdigxj+adZU
v77jN9nEuV3XIQLmNW2UH09d0ZijKTHXYWyXy+rNMDgLom6mPIvQCK1YfPnFFCWdQqdwRNGIPKbx
FubKRge7n6bgEqHz5a9m5c3BpdyGjKaq8GngEDsm5tuojYyBmOt0vy7KSibA+SvjC0NsIDBLl3vX
kia7M6PtVwWqxVADe4ikUQbVIhkU1YSu4n37b0ey+lzCvvxNyVPNM7bATBb/iB7ZAQIthBQjiGBL
CidtLBVsNN8oEk8E7XsNu/EQPR914wsz2bdj6PI3H0MWflY+HC7XfHztBHzN8ZeQDAat0+Oto462
ceNYQSLQqOGwSPi6pqK4n+hbuY7B1rxZgQu6psWvYqwFcN4bp9UBanoLYJvp7wwXhaVir6lEKKEN
uxJmBkgoYBtwp3QRuk9pfcaNGge89V5dCSeLH5EKJZ+sEYIUDHYpmOxtt8N86pnkhYG/4wc9PwXC
TT2mkuJoB5Cjj0LJ4FeIqUrl027qRAVkmbt2QySXqKJXCwniWR0qLlO6w789riq/OuaG44qT8UtN
EknW0axHgLB43bgMSSkOCqiU7t+X9fIQ3uoSBkHVAHGNd4nNoBaM4DBCiX9nIhhFnxxagMuepyDi
/ANjNQaBPmfMYnCBCaFq2dbUAkxX1pOa4kcUA8qGJ39DsEcsLxBq+jUHNUAs+aFC8VChXIV1A0Uy
C7JTcLSV5bHzvCltAhTu5b2VjGqADy9IkRdEQ9eNJzLvNRNxC4HgJtQsAboV23XAw8DdtYxa8E/7
M8zkoEtF9oVi5ugj9bu0ZzGK0Mg6J2LAd4E8zs43jON7skcwcido6hLfdiFSqJnQIHVSGNaufAga
WMKm1R1YzVZUZP5hC7VTTQoVVbEW0knmVcdvic0Tcl8FM8nMDBNyIK7+NuFTJO4TalSzj7RXBYap
oWOMNWfBCMGK1PGNoqaoFcCJsdLpKhhD/i65IdXKrylaJD76Bv4KFBYQDrmQeE3aCSvrXvMWBtKD
1TLy3oaPVVV25GYXb2/GTMrIOHc1fvQJrIx62Tcqrh2nFAMPoNiq1j22dqvJuPjACnNm8HFfqGB5
IC+zuKdgdEVfSeafpMGRsHZsk1g5AjfzcmQGFhheUKVUFxuOAdd9yfPGSsoAbYghYJasD6cIQxnv
x76SszSiPNOjJio7S5BA8VvC2dnB+n1Mavs34z4uP2rZwwHuBj5MloqvMNQFxBp0taQN2uEAxua2
+0mBSqphEjrvieVuAmBXjyYbAuETZU568KzGdmbphDfqz8Xa1jul187ZSBCQWv1XLsv10W9+oTWU
8s752I//MYoGOwwkIu/kMyWuYjubdvl8bORbF6as4Hg9AYcGtvKgLypNjIhU0ktQ5UgDDqHnwxSE
r1V0JjbSSW4bQwdRWQ5HYM631geFw7tO6XRYvrMlQwTeLGYklCJ+M2GQt1haTR7lbu9u4mIgnxek
BDPjRsGgWKPE+mrWmaNgyCZHBtDbClQrldBvou/32N3MkjtnqmAuNEo29lA/9icRHQdNlB6sPbff
stE34cEYnyLZYpBWs1Uyz606pPYpjp9+Q1hMjzyQhW1yOp0w7M9d/fmbZrsut4QNloJRIOdBkWah
uj2XsdSrGjlunZhQdCPcaGfNTpwgQ0YUBI5Z3+9J0LyHLAP3mEo2tgTk5h9J5d6PpDDfgacI3D4N
X8FiY6AoIO/jw6RhyCAjbp8gV6NDz2YoQJSHvRCL5VERSRP1E0DvBuVCNnJ9H34wIG4SMltdFGcu
gAPsRN2dWEoCmyjXsupKS9J6ztj6BKqpNUumR7K6reuzWqhvK/zkDMN7h+NU2Wr89eQahzpCNkw0
T9WBnIzUENY/vRHMTA8lBcaGO8S8W3C28gapfNygUbmfNVfcvusQqXIzQ+heHzjmAXTpEGThcILP
N5vIdF39JzR9gix1gcqyo38eAyJLAajyumBAqmJaJhvKu3peHS7F7vmiEVd3TXkGAdMAj61hwxN6
eDwf5jtw8AAqAFIonZ3KiW14GL4NdLKSSxtXJR5rzL/kkdUWrzIm+T5IMD8kAmanwLFmp3FlqJBN
VTRu0c/+jpr/zcLrizTKDutHmmEv4Hux+wRUO3h0mb1AxY6TviDwWfArxplUw22Kc90YBRVHZ9oV
vOoPvHofrEs9uy9rSXY7UwacS8uB7SoHURW8b3CMBqC0BSmKEjOUHdFVRcEqnBETXAzA2FVbIBXy
9tatryrlBT90nd2C8b+Ar+Gqp7jO++a+zKxNsqMnmnyVlA/G0kvsyp30W84oCM5TVr0DAymTWF5F
MYbEIMPuOVs+OAzWB/V29I9oUMV+s/ARelOFVQQhkbN2j3rn1oebjDiM/1u3rriUg/s9UVxpCCWS
tWbLenCJF74/qmJD/4/cbtxAgTn43scLOq1bn81blSSxsO2UdzqA1+o5JR3BlVEad2ZiQ/R22NOS
fZw5SznvYPIKIvJikX9zrbJ4dcSTDxjUNrqzKLPxn0jK2h8FxegRp2dbhtM0xmdqojJFj5Uv++YN
dKZQPxPqLfAyQIB0CYBkFJVjNZ30iXjzkxgfQfETf/ugN8ATCer2ssFBrwkYVe7TSng/Pit7y+wr
ymeaGSL2cA1NOn1tnMdXv6eYRewDsRxW4q1BiA1HsYLcnkSgiZU7tXGQufnh+QSXwmRbydP+BuXU
lazeNQ3JDV1mmD9G+3DEeBLDYAmp7nSwxVlPGfVs/tIayqR4BKm/uO8sMd/L52YwQbU+OS0Fo0WW
2NhOz6McsgfRSkYnti6dL8H2heEctUc2yJLON45FbxMG5n7yqci4TZb+v736zjz5d+FS2xgwpPCS
Hup94Uay1yavbu1OSmxntpOMZ9HOo4JY4iOZdZ1tsRqZR21UxqvhI9Meb8AZ1SeF1u4tTUfZSTa3
lqRxHWy7jWMzqWnw2gIp1lJ930foCUKLsGnZtawu4BvWncfm8D1FYV4kQWdAQuCAZloMi3NSkIqk
4RqPUyFmYio5447T325PgjW/4HqGobIJ5akWcu8AuUIzzuilqZXsrbC6B0SCsbCkVS3tIpG3AyUv
J6VIe8oQHaMugR8tMxs9ddGm0e0Sbj31nWII7q8+HD8gwOIv19owUQlCHX3XOz/YOiNBNzhxAd4K
1bL40e48PR6tsmqDZe9TWkOWYJ6hq59eqQ1RZ4HeMDHsv5immtMYlavOoRxDj6iavpXcc2pIyGGN
2kMwseDhHiysLtUX6gK4GM1vbzgsIZ3HmqicvbmJUfgzDmfyPlHzHpFz+sBX/BVcD84JkFc94XO9
9GoR8E1ps8yfre74JhAlW8IuWS9BPd5U3pZmEdjqnrRnGkEEYN35qppaRrcxJCjCwp7BtPVQfX9q
qx9AeLU2/psYngdfo+ZCTWu1E/KUIA0bVY9pChhvTY9Cn/QEVJQyrinwhQmC3lKJx3yH3dq0Tex9
EGN4pte0FevpnRdvznmaP11z8QOd2Avd6u05NY5TYVVaSE5PH9gA/Po+pM+iAtVx1IP03UhA4isZ
6ZePg20rFMrmIhH1Yx5mClyIezQqiuAXjiwtlKL8UEiKRguFlHlT+BBVWH5SfdOPHfDpls7i2rUb
wQj0hJxksCFCie17vBb8GPfnxeDNikrA+rmK1DSf0GP3sVZagDAIttr4L3MD5bv+r4uYe6lnS4Ou
dhA3SiMfoO7+DAksCH/NL1YOUf1nRGc22xFhcK9xjVXBaWpgu6tV1sLB1FbUl+YXJesHoU+cnwTa
n5xzy87riKcN/hf0AKfg6bh+wzhN5prztaexDv8xmzYL8RsbPZO+h9NJ2telRps3rZCFQPGhaXsz
l+KqJUCgdGVUhjPZeLbqXlVJfVSPGBRxtbBs/Dvnb1y4SX4b9QGRrZUSAnczLNBKgs4MEXStRzTX
AGcq26yMhPhTSTx0yQm/cajVtVI50ubkCNMpeNn4qJ5SXtn/rEPmWMiMpiy5w/egOfPjLn75f9NM
FYiFonkxFKfj39fiZ8tOEeCrxvE7z47UOdD9JlFumzCkHDByikRTJuKCGrIiaUDzd/BswhM4eCER
rdNExRmAGDy7GSnxYx6zFGvjmP3k+Z9As1LHm25YdSf15rcpWom++uIANnZWOCBFTamUd1sAwMkW
rP0x+d9HkrnZNI4w+uPn569WVHo4FYRU4cHfVjpnkxV8QjLAhK6zjk7zD5giPIqFlRtUSaYY3PuI
8FlzLkijcVeIbdYfTatQE9+lL3dKOcDUyhGA8D4sNrIBbewTdsVDb+OXuSxYxMbVo/qPuVqyAx3U
wsGZbwq7ysqmbV2bQ3165xZE/TaZMcGZr+8QKOeY4pS3twx/xf3u8xU81NB/gNcyA6fcl/tjaBRO
9UDT6+OiXEyzedBJMcefM/RbFz4KmCoVvTKrWIR5+D3120PQlrN0Nj5vcIhQzNtXGYG1Mw+eFyuc
nff3oFkeuIMemzesAwWdhY9vT8nLZRV53GDqQICmOEnYhdX+H0puJEoc+JWX6c/3FQXAGK3nB022
vxYtwrzJ2s+cXBte0vwelvEWDjRehLB4Vx8XGgIENd7+e+W65scst+pk/KkEKVV5YIZmL4TEo3d5
yESIFW/3zOcNizW2/fhghqiMMUgrhhIFmdHg4JgdZCAho/OK2Cg7p3rqkOQxmnlE1tWGq78HtqeD
Z0IkOppk5bMj2BpbS3/DGoKIMy5TEzvkfHxVBuILclsIYw+ZOo1CUXKqpxE/vMelkomSaGr7/Ehe
O/iQX+wdC5Qzsia5nYJAf1NvUY2YzGNHZpHxHPUfRRC7BjrgE8w0JPaE/hHUC/G3orOihqv1HIUS
2cQSGrTzMAD1auAF0aeRDW8nO9Qfu/1xHyAM5KnCbHEPRSmy8Bt00Fj0pj0SBmZ+/N6fO/3j7v/b
XrPnYio+miGSZW7E9knILSis7YxMZII5uyJ7iAGwXFbwWecA3ai2emHctSZ2xMhMVAUTExGegakk
M0UFhiFsoeNa80cEThPrNn2mDclgZbHRFK0bVciyWcdQnli+IJDRTrHvx7kEYYBqTwVyGjeFLyA/
oqQ3q5hg71dnbiNkrInlMxGzFgUHUbJhhxWqpKeP/Zwt3+YVetT5UuFpBX3lpbxs5qRKLq4Hvp9j
BhVL8RIwLYDuynEapIgE1Hl45WygIeb/sp+oi6lRKFozpjRx4o8W7RZ4PH4LFMe0GpdQWMh+eMZI
zD1OIhzegeIyf9U7c7FWwhWCbiEqgN8AJcvCeChLjdn1DBex7WFBgg22AfaERYp5jZYiZ+VkLi7f
Nz9M7tIcL94cSBu3GtZRb+Xhk62PlpI/e3tKRLTOZlk4J/x0ikJkVk4YTfXcRQT2JrW0I016Kv0w
sf6EVGKhLYi8I8hSvWkSQgo2grPIm1RnB2sML7AQ0z/r1Q8t/kAyVyG43yDfWrT9B8Bh7TcHL/11
Kew+gF2TyZQ7RxB6VVDjhf3LZ/ANf4eXTjzNV5QV6wP2ccZU/fEYUjsMLjxInJrA5VE2/h4AtYWA
CTxw5LZUJRt7GbWvcaCVkMCmUoRRm4ckA8BvYzy13dGlxfVLe2LmNtYtKtCbPPJuRmvtypLTvGd6
qBDL1fmCVNW11AaF0iRReGdLv+Rbt2yLLsgFmzxuP1POPtuh3HqEpZChFHfG9BXsBgf893+y1lmZ
6TwsP5JwuivYvJkGHznRi6F54XfZ/cUDy2h+lWzdZBEgSqb0m088NA38K+6J2wLx/hIyXJ0mDj44
RuOUG0zI+iwKDb1L6OnCAADDN7bsqEnH6NJZTYFvHdzHdZYFsLSdpi0XbtdsxgFPHkYAFfjUpBe+
lPJPr4KVkdQixj4xtOFrc0ad6P8xHOpQ+zcp/e/N1FC3erwUSPB+v2hx3mc9PK6Vs8iQKZ00s57N
/U021ODiSNsZVb45iCyPfMqtSl5UeSgvaFoLWMu0vYgrVpT6xEpItgOqKF4vwJGJNEwZaKuMF0c3
NYZTAAbpSuZvLvATGNexgsEzbqFTiLg2v+AW+Y34kU6HmzvxoxJGLLriS0umLFGTz/Alr0b/mUub
7/iRpCBHIKCVVgbfeO/XITAVgIXrw1nZO+plTNCGHCC7hoeZMpUKjhXsXetmfGjJWc1Q9JzOMbbD
iM8LZzvXTdq+BPeoFPQ3iyP6Yu3QE+/68kIjdDjTwbKotqkzJoBdTdRTnFaj7oXOhUfL/vq+nHrO
JzqB2DF8jQUylv6mhgPiLKK0O/h51s0akJA81zPX9VrmBjeX+mtZDWYp7L6TjjgWpXsZDP4DHBuH
QY9o+ITKAvoWnQRa1Zbbe8fbYqI7yebpdOsXmAuvxUYE+WTjbufTH6+tYc3q+xgXjaRFzVWVVVqB
neLooYxhKo60PWLLTg7FlLyMv2ag53d3a+HRCtcp1VXvdLujVd9M7r8+kK/6k9DUj3+6HfTFEY8h
xc/ouyBC3jgJ/5rMkHWUdX7UxjAQD63qAKFtvRirQWUqyQZfbXpqBzcAF8nzTPZbrQ/MdFMWGCDK
9dZXJG9KDlmcQM/lJPGrs5qUuGL5MqNwJFzqJy6ZZb6/UJg9WhPmDEJKLsjeQy9hgFiEnJrGsF8U
lXL+t7MOirKINVYh9RmV+y12/jUxEgjyGVpSITDBBkcF9roet5y01lqTUNlqn5E0RGUZthVInlsB
tQ5oA2N0mGIw2rH40/vS1Ic3xx/XYbXCead0v3zjd5xorHckZlYe9nVt0Yir1LbzxpPVOogrPuMz
GEqefSZAYlhyjB4L82IWo7SsYwQNgQtEZII/dFnJqajhs99VXObTiiuT0XGaApvOT3TCJksx+r42
ulW/UbZiw/bcdw+duMtQKzG6JzdOTwpdqzx79/FVPslUtZ7iRez8OGTVSLbFfjJY8s9ZFwO3NUv9
g+Bv8Fz+qaAWvxl9DeypS4bPZlWpQzSaibmbHrrjncG2/fNyRwUhTIVaL4xmXLiwqoQfbTJVGUmn
diwqEeLwlTtc+TBZ1zwZX3MqR9ou6QOHn5tO2rHqrZOjeNn9J0qdSNEtcqRJ8uQt53CpR1/kEOsg
12JptVvo/trC1IdPFr538KGC2RwHisx6KptPVZFO0SWibGEhvrrHSZiq2mE2G9q6Apz2tdt6rFdE
Ip6xJMPX4mHK1Np0bWbRedGdxP7hRHpIs27wl921EyKTjw9SStWhcni5d5M2ZtTsVnx9pyQSvWJD
WNWTICSvzLYaClvZTiSJAEnhbHchKQK2AqVjBiMel4HEn0/kUpqGxdRbNP8l9hSIeCUThWlJ5ZOZ
6oD2LEWdfZ63Lzb/mgEVFPoBrofkOplk0YMRz//xD6kXv26NRV3uS4SaoOyG31nhAUpLlv3X+91P
5I14yKrZRENmgMeBIuyure4/IGgaiLJwQotBCFoeEnoGkwq+e89UNLa4jKfBVIUBh8hHRIS0xsTs
ilmcFz2dw7y5taTocFCrXhaCrIhZ2n9pXub1xk6JjEp1ySc1i6qWTiex8Jac4um1c9oVzUdcWqun
e/t4B1RLZF1I3UuAn93IOw/hDx+vqCqSU8bPwsNL9Qrh3VnZldDfQlBhD/b1LPNHMNpZqSqwgkcc
9vVKKfLzU6Elv8P+s7i5sXw/d9W7VyFQ2spiBlccrjMIkTuXLqlFf7g8Q9BJcDw84wAYn7g0bBGT
EVK4lq9vJi4V66YZ/krNBig9Bn6XSpmRBBmewEKt/eQNNwn4zNnYZJkxHUkLaojauv7ege11Vp6V
K/ymLOWN9dksRC4tcd86bkXhp3pW5lkNFYhPL6Q86VEMMb5Mn3DErBNjKwe6HKGHXys3/56hycoW
F1mpoOskN3aiQwcGRY6dnHwzmvTrGukJmAXUkLHe+77Wc8j5jbm2Cjswuiv6P61w7oVbkRxlEt0H
R9h6q810DxD8kBL+4NbeHZkslC4zaBaRz9UmlWmNHzOvj627cySHVwWPmHix0S7887Va19s1yzbh
J85SOeAks9Aqe7Vek8Fvhig5IwKCKX7Ec6uyIjwibBW6sW4nc/p4WcEeFhDlaZFpA/SK1WSokpbb
o3uRrbpG1QUAZqSehHMOm6mG0NnUNaYoyGXrqeHK3lDIKu2hOvhfoU5SgwnWwDudgJhBv8eqtCCZ
9esN5MOrlrQSbO5XqXwbLWK/kq05af0+S+4vAqng+oWpphVWhP6lTRY/LGJnH0eFLv608IPumVR3
YG+KZDdR2vc3A+vpotJST6DXk1Xke7MiphGayAy6sy/UuZ084IqveBqDN15qSxaYeQ7c/EKxlUIt
p0eezRoYkjsrrdB/DaLIYMQqORo6LZ0xwrvfbiEcBQBlwVlmM215ANxCMx3IMWj6g+sc6XLZdmKL
wlV9oTn6zkSd0JssI3RDae+XPPv70T5SYNpqftmhBLdbSeZ/vC0hKMCvCI7azRMnC7jx0RrbLcm6
Rc8UmSXK1cosVjISLKcinHjEssNvDlwVQUBS+LIQk9Hxm2viZjgGE9kDY6JVPq+b4uMjwSfbpKuu
GEQX0xG6x/Bj67+o8ien9bO7ZluJ4FzyvRfyECS2xQ7LGgacRBs4TJa19+5W2+9AdUty+cc58IvE
l9wHDELHdd8tDwR8ek0ShwD50XxajeTB/INno6ZSP6rtsJob9ZJtrwqD+y5EP6gSV1AifC0XLKjC
CREe0M16ptQ16r/8F0su0GzMbD06gzYX1KAyQUYiyx0e7vcfXPR1AezdcnEo1C1YaRIxwYo8x0hT
JOrQJBcsJUMwe1TK/kiCvojlRxxzo8Zk1+BygpuPI0xyceySvnff7TBvBe2TEsM+nf/Gk/GBdu6t
2D952rdV64aS0X7k4Chq9oN3MI1Vh1VhQSVs2nfochm9Kzq1KQjGqwp1X+VB3rI0tVWE2fLIgsiX
65fylVq9e3Q0jluZgwfGv0PJxfhQ963VuRDcsFDtFP6ea3H2LFERbzoYh1fMnXqhWhNy07ohaXfs
WmMuoLdeIK27XgMnHIeqAelZFAYnTB4OlUyn4tQyzgLV/scDhKIioT0PRQrcRgTvj5qkiDzg1mwY
TnjVbd1y/WT8jWO9TAgrSsR2gpyHNxZolgQC2pzhffMWXdgUdzlxu8ulOlpg6Jc8WiA4L0MkscA9
z/cntgOZhlqz8ROIKIJHR04OP5AjZsnrzA/XQensDSDDd8SxmWNt0vgywtGEE6plPv63ajH18LRz
pZGS8ff6meeCUSsU9h8w9AAcLIWK3jJBAVk74ztoFsD+vkR3iQow/Rl4vFqLuJAZQufQC70+x7vY
go+nl/ud52sX13vtanIufny8my1JupONgQEDYGK6EZFDUMoM53EpDpby1AV9WaYhBI/ZvCZ9ju7s
D4jZqN1esi3jdLT+DjGqiRHo1z2BNCg9sRsWZwJb5I6Wh9/rX6pB0rxiarRhGJf9ZZ9/ptq3K1ic
bkL5y5D9BC7fHbzvA3RF9p4nq74OCjIuIKm3ttRkcrq88oPrTpxKD6S3F57W15vhxJFPEbJV1Pck
pjkSKSMlJU/sbqdIwnF/NClGRW/1PZv9O7ncftgkurhxXgeRwu5JXPqfuM2o5RmJMqdZBJnsPUF0
7Z/qCcIj/jlAUm+S6JIavE7gfNO8cwsRzr81xWmt5hOvDFh2TbYqhPQ3j7Hcy27G1hYMrq224U/y
knKNFGXsbMed1T6UwbpBkQOrhZWtgrTAe76FaBJNgadOo3eNrfGDLgVc+T1ptxtD+39GZfbLm5xX
ISkM4TT1/Qi5rLBPjsYFMF47MCiqqAzVWWzSo1k+ewmx/p6u5ppwAmhnVuuTtWrRLz8BL/xoLoev
kUsoFUd23y2CqBH4x+AakKudKog4MCROa9T0ncP93p626NWnjhPNZplgFO1CfTwEaOrY4Mcrs5tk
5sdwXV+CAQkAXYNgKCTLS3zlI0JhDSVO6DekTnZYVsb6Mhxh577IehpCVy+X9srMg8RkFWxjsw+q
/jSvFqewSYgo6oFGcRNtmNLJAyPM+/8CRNNKt5GXrte3wnckMH92PWkOIN6FmjgMWrQ2EZmbh0ow
sLT9cvHL60FO6t/jGEUHH9LWxgZ4PyDVftTNhiPlPbjb7rLP6npiu5WOD3kcsXKKF8HXISxC3u+z
0917Drx/1AjDiItQFB3o/VCCdL6TOT4xqquyVATwBb2N4AEAHjYSyLPDQxaJfBE7lm6xtbWq9CbA
qh8JHKr+eRKgSlRPJS0JGxpVo10EQlPX3WQZLWH11Fd9/byvFjufN5sVyf4wk5pCODnvWebk5DSa
8D2ax3Fz6/Tq1RYrxUBnpuo1WQ0XNrPULAa/vyGF0eJoYLKxI1Vf9iBeZ9wQv0MjHr2bKxdJuTeL
JDQCA/3Ig+UvbuNFBzXJ/ar+8JXmwG+vGIVQM+uAnu62rkBxHw4EwQjCDQiWJI6j/zLYaGUzXHQU
DpVispbsKqoXCcrMpv3qp+RFgBkWDXKpV/1sKYBpzRqduhec6wwN704N0Efu4HtAjgP6PJwSz/Es
fqyJhEShsMLC5CUhkNYo+h6W4QJS7Ns8MCNX3gRp6/vYZFEPmcYRzGcB5F3xN7wnzqot/bGToFPy
ZZxXNeRDC2pKNdWyRFBkBwoEGkJxvopkEuV+e8f3geo3Jop8kZWtMd/e1K6MwpvzNmwOqHTu3pT9
0bsTsbkhxHB6bhEwt0Q5KszdDBoj9HstEEGlgz7kx6fJYBLonn8apj1G4psjQ/E7um5HOvA7j6SH
zfWCJgvln+LhdxIpUlZfXRIVWPHwS3PLBb6kWjfx+K/YSvsvYvTbs2DzDOABNlV3+oHY0UluFBwr
qiuOyhw9vBVyuyToaTdLSCyqZvcHcdcfj1Dabz1ni5utj0id/v40lh5xabw/8hlekuvC4XNuIGRx
4dKUh+63bAudHlSZ1HG4+YdZoCNYPxZ3RPnsBfPbE5U+txhOlCMESUEypT4vFr8no0L/sefPs+/1
qjd7r92BTcrLPYS3AdLd72XbQdC/B92YxyG7pUJMh8uMB0rTzqw/TmvOajavIDX39+FXLMkwIael
ycBn9kl76KsP/jbTRE0PqlY28sBoB/llXd8T6/Ip43iCXtGeozOsaM0KAk3rcg42aBr8xmGqsYR1
ZJLZil2rLTQmg0ZHsi/q7zhD0NEfo9q0QfZWcngHh5LNLxaDpzDBWrw8ggrNbFO5CyM0X5qycBdt
yKfoIXJhSrBpxqFGBiDEwLsec3LmMEk/qkQn0mFdpJHJpYU+RlZ62qC/Snsxb5tErTZ7MYNjHDtK
XzrqsHnNVXSxTNH7nbBWDLE40vzowhfBvkF0oiUZ6XJURgEx3W57RUTgUrHYNAn0AxT7KHk6VWVt
VwvHdvWpzTlI/YPBAo8GpiEG3aeEduZ/foJQ+MIXIeJVDv3apjumualmtiNPVr3qkQEOA2eIif1s
7uTHXravnHuqEZhFK32890MNzjRFoDhauOnGcXGG7d1Vq0S1tQ9T2kKlPckzNMrtgGo333b9FZuA
rAO9PAKto1M1Bi0tKIqrZkMAex2whtd5UF21hRwfh0EDbjrXBDccoZn0sQHxnsBLFCZKgZAIj9Os
rvGSy21tD7+iXmCbUv09fvHX/3Jf70Ld6vDHfZeeCA2pDJcNl7vURhn02t5CvUKA/XDMJ0fVvxby
DQgdZ9iS8tFXVh5cMZuEw8XzD5xuI7SkT//gS/mZ3cic7ETZKJXSvWWhOK+gBOsjBF8/GLW9V++0
ytas/2EMHHZIsYeGQn3wVh5H7+UKzbY67LLMOTsr9sCez9fFVbL9uOe0fTXqIpje4Ok04X/G9hD6
jJGomxd6qFdE4SVBeR+GL7C1BtJWxqrsoF2636plGiXv3E8XRvfwy2F7H5abMadQOEq8OHMrhaZ8
Shl3bBWasy9Et5rvs1RWO+oH8LWZlFTSqg+DKzA4thRYP1/dEWA8TDKOOAMItif+6BuFcru1UnCZ
qHEmPTSH/6DkMZVZ4MGtNRlmeupqI7wk0TcuNprVGCGcPtNhIJxO6SOFSweufynV+tLEw+odl2Im
aGefMZKQn401g0r55ZqNTb67yuvK/83hD3bGbioRMqQpmMfsNe0tSg2MYWGWqxpMOGbpqBBHheDh
8f2YEhIssZ5FgEJhR8NUUOS6NZNciXjHZWi1IWBBsLSoeVaVDmDxgJpm3YS7TY3qIQMen6EoVs56
lejCODXw60v1hC9+DqwEiO3GEINQEGbj/veb508vYbQE0/ThcuaqQbKISUHi7iiJFf33XO90XiOd
ZC3awsEOZc2kj6qWVYlNNP2/WkxZwkTVrO+w53rWTxD2gnezyqsPfug5PmLGss3d24Tjs817R8A+
YWOfJTUfEdS/X8uBVau+dSSQT5IAcUET8FbTnlAT+IXUWiJHs8IRDRX017bVNjHMd0G/97FijKKm
72IDMIA8jc7xapcVDahZWR9svKCsS4vxFBCBi6ZYj0DpYR2Nk7sQQaGubFAcO4MQnkB9NzR3jG1f
JOHam97rqPY8AnJLdmtqob6C0WA0bD6ODXqGz/flU0loS9VOHAVfSbhukIHl0JF2OiC+rqxl629E
LCyrLH4QiTi6tGtgkLjk05j2XTZvez+k5CXnBpDIOs2d8LvtRtoepYQ9/CJr6Ha4QN5QSw70oCx0
ROP38bjuEayRrdFCCHMG9xNoJGCEkYCxXqau8CGAZU+v6vcktRdGqTLFdHt0nxSiMkaPVsoedXa1
+1/ymh31zt6E4uR+zq6qSHI+516wwiMucxZjQv12U+VjDPioM8pDUuPrHNSqOnMee8AJGHkQsuLF
IISy1QFac34JqJRTKfwyPqVgET/TtCNPjU84MGkQdgxrraK7a0MkZtGRv929vSCgkN4Wm49fv1Hx
RyTtB1DmtXDC6bXSWts636eKKjrJTNt2+GMoNa0RFeoBUPAV3+Jn+eqBQmTQOYZUR6pEguLD1zeb
G48AlC2x8Ohq0MQer8bUgmhziXAFZ9MOcplMfwbVREdJt06XZ5hB8YLFO7eMo9qwTNwdpIpLXHKQ
2vUAPyusz59C9CeqYCIqFYgq64aY/W35v4E6iJYJhFuqkX2SaskYU2B35PR2PZ090kTdFTcM8rp1
7CJ7VOndvaKUZiOox9gFGtdIkBXkhYbVTrxE5Wcc1rxCM7iiWNNbhKXAZDrDBX/gQ3MgYbaKZQxx
KzH/tT/yzuRqKlQfjSpwvkrQ90VQOYwI4R+5coG5TPHX953sDhcSINHleCxYjOiy7XZJlDFAhvnZ
EcaCitzh9Ohk/uDk+T+f4dMf2eukWRTgiv9Uuy7q8auHQCBBoTDH90Niq4hGb/JjEwKo7Biu4Zei
Qk3nLkItB8Ur3UJM1+IV30oyHT7pQMQuuB7psXU1MC+hwzoNLEXIaAlZild/Y4uAtxixd6KBQaor
abTvCwrP+KKy6tIAuzOzzWf9/38klJEduY4H38xV5kfAl+zegN8ydS0EMwX/d22m7aJGzm8zeObu
3Daku9hrT6eUSlO0lJrNZ4PY8cAtPnA29x432PcDDyYf3bRo5rrIjC0Uktx4WCtnH6iXg2WxcSGY
NPY0EZRixVoUp+Khcyk8aDSwU22eP3ix0EN8m+bhhwjw1S1y8j1iwG1EYcf0UrfHZXuEDbgPonFT
Gr73Ycce4avMUYtuNNlFZENlBXzNegi0Ba/6IwqT+PqGY/fRpRuKl5SRShtrHD1cqjrqmg/HwA2U
l/TfV8K7yX6psNb0PoasEXQbujlUCIkILd7a/xk8udPFEo0sXmD6lwNOQHamvN1DoOxhpvkiV5bI
UC+1x1wi5nKQ96NfLdkG4Y/azuhWAHBCSa4ZPB1+aHTB9i86PStIxoqAiV7v02Ay+UvBEMbVYVjQ
qz+5zpxyQFg02o7LwNKy/v4tlus7ywlcVcOTk+DUgd065fLbW7uqkEWUcHSEpzJOuU9ROn719BEs
g4jnywwvVl20px8uLFvsFeVoVW8nk2OOw1ROmdCK4uvv7keG3ImPNCckRN0X6dOqtGmSKRkVayhe
WESdvfOjdQiMLEh1QHxwYuftKaWlSYg4mAh88Mrantng253OsM+lFfBki9NaJOnXAmO6Kn8gw48n
z1aUw1ZlIr+nunrfixTsw6RIrtDEEt7lNiW3q7x8DgU47IJpOmDmQM1EGzuZWL9GiKUVgUkvny46
7QS0WLu7TgXTllpnW3c4UirTptXyEhYWnP+CuwOXsqUaNjwUmvpodO662Do8K28XfAXYt4MSn98V
EaqD315MLQ6IKyh9Yaa+xcl/DXUl00SCZN4+1dFaynaBaQJML3x5d6SWyh7N8k8SNz7XmYEDF6Pg
Gi97g7hXop/bj21kiU4iwfT5KqZnu/d9g1ViI8gKg8b78krtBB3LtL0EE855hkD3j7ZQD0wsiSLq
i3tcIR3q5b5TTvZQRNkbWxGpBq5FqNlnWJElCPZOoXojWSNZl277LzNNvgJcYCBMIHtbkZIrroJz
VZi/RPYmiWir+xt+5lpsZCKc0l4WDFEM/z2y97jrQx+/nSebtoYVNvOttbBJdDz07egIbp01rsRc
weruixxoemPvsOnLblgWBQq4WV/0XqkUEQOlDCUZeKsNxd3OPphzCTLT2xI7XBUXzip9ZLbGL0v1
OmDdDsoZiT/VL6wlxBI9YhPYB7nitcFNZrrmcfebodDuh0DSMhUVWXs/6H/ETmJDAn7O41zLSNAA
3iiC17z5TUC9iGBFnnhEbCVD+3Z1bIEoo8W3TlgZd3lSBV5ilOh4R5cbl1mc4sFyyg9UtWjAseoG
v9+v99vpy9kSifYgwxroY2QdS4K9VCybdnziVR7TwT+JUdtzxMU8FrSvuwYqoQLFxxiUVrOkLzvd
vXAO/qJIalzDPnjLo+xZDSQ68vIoOdSZI3jntoaicL1CTuQ4EMYeT6ZrhAXvYN7YWbn5wIDzlmK2
iRJemlZ4nPA+5M5f4rib95qHb8jOeqO2Q0DUlewpOSaU6Qvk7DPmAMaGCDSVKdz4ewNij2XB+bQv
vdy7JtsfrP04tiFNZxbCykx2NuMBXUyMfhlDd7fMILKlea9hXP6O4xURy/s3y7mf39GRF+XiW84P
gsWPQHcA1JrZmsX2z3i+k5bbnY2FiHEv3nx+8TYFu8E3GNm55vqqTi5VyOwkst5HofcDwckrtN/m
suOkMAEn89Xb+gvDiiUnvucVxhLT7Yc6/ZWb5boPe4jy3BfDlUXftxYp/oXY0WYX+KeN7Q1R/HwL
itRKNYmAhHI+MLrU5aYqzXzKaTAudITqPug+uh0J/pxtNfmfUSxYrAwvO2Sqv2UvS1nl30MMTEio
26IkLDR4KrGhX65fc8Xiq7OhoiPYwJv5e6VRpMrgpY8+cH6r76JHfxCs3Ur/3mK2QtrRe1k507Ig
C8gdxsH9FYbuNEfdAW1fNzALq7Yj/dF/KJCKsg+YPtv7JqKKDfcGlRYH7kQSrvqD+hYRzYGI+Q0B
OS+GHFIkyCsJFZSSujxEwkLqjzEpieEMSI2w6Byu+DvJZheIWR2wDzyTUQvES1K5EnuWSR146YFW
16bBqiYEPdICvmhJWQmNSS4MdtmXWwXnpw01EHlSl6fEvzKF1o7DwphKsyn+6oU4hAvwWA1cN7ha
WyKFOesw0nYdf/U4zmK0BdKI66ir9b3GEbNAIcwC3bDtvuUBb8WZZw09ULvzmq0idt+iH1f/tJB4
EluvBxXUu9x91oeZQTzXjbfaji8HGJ8iGH4P0k4fF7bFBVALAcj+soAkLk/TL2EwNXFvbbG0FJ89
2OxOW3ZsEKjSXTGMVPMX59w4rUJupdH5yXDvCTE2/OiLEePXMOglzXi28MpbaF8XHpo+8t4uXMT3
kbcKsIUmNcPlHyzD/0GLRUixyfeBaG4dUeARcHN5ozBofKOCECs4kseVaJ5GiilZCPXLR3k1KBKx
ZqyhW+B4AwTIR7Fy13EE4hTpM8FZZTF50q/ZZZ0KcQHwNl0LhcOKSg6tzCk/rKJH5EaFpLv9Vejx
j5rty+saHitt05V+5RSVLzVWV4xFjvBKXMkHRDX23E6O3DN1kSQvlLe/9l3Ho2j5T60hfh6j6xMS
IiozyKQiznCyO9own9ZzJrlKC59cv9WlojCjvd3q2tY+fk01XWbLiGVsRPtqObvz9WV6zH1BXuws
Ze+i30YnaLPBXTlB36Dq4L/kN/Pco3hXxxk431BQNEu4g0AchIEp4oNOmXSG8QXHnts9jHyPSEHr
YuqLtRCA8vVRCiImt5V9RG4DCXKXf9M9RSX/6KORTw5PAdFYPe9pBu4huW+7brfV4NGrjVjsBWAg
KDtwngRay0NS1gpTfKmaneF/wj8GvpwrJeU3ruQjWbUnzubxB/7CAwhBUA9IYpejvEVT8Ktg/vjU
Y93sze/fB9+vQLIZI2u50NltDk2fc90jN6P+ge4mme1XyCwOD8QWCbO7H4HTFRazptgdGOUoDBTH
GDTP7TNYOAnkxpCfUV/aExT0YIoxwlL0k19vRZgktXISPryfTAaxYY1EOZnliLw7PwB95dN4Locs
xcLb938e23aY3QTZJJlJoDnR8CFse1/8fh1jliDG9WtzumfvKkLfRD1ii4JrtCthNuHthEqqJsSS
5dZ5zAnrfEvihZdqCVAxY7j9oSNtg6B4WXF9qH++Fd5aNoPnE4cP4rBkczpVjgQaQQWNHllqmpeI
kJH7KaYQ85MO7+Rop4UQBY3ZRnFSvbojcc8c9Q/ATzsxAiS793oGiU+1HuZoK2iJEq2jvpCkxC0H
BN+BJgM7hFEQ4zAW2hPftZ5BDxE50agWZnVLhW4eCAmPc4NBVZw/x3X0MuBy13oRVKSDE+HJqgyx
pnk7ZheZSW/YkE65nFJKcYfM9ATzSOnXgVWtXscBw83K14EcK2OTFDfo2scRCq5+niAyparO6kRA
u1ljQYL/CJVYxliOkekVPFekbBB327S3h3AHBTo0UuPmSaL+vvSP4uwtIbrIa7H41SNAOme7waiY
iGm/lxCAeTSwxeAx7Qoaxabjjl2WJGM1woRMkW3Fh279CHI5BwF2kwAm5wtcI+jwXGrhuq8NcUau
V4yOfsh1An2Ljp4HLU82ePzsbBMuWqy73NIoYn8djx7E5223BHPizue6bW3/F2F/rAVnuehBJMvn
E/loakKK/FlVWPxJFw72bLi2UkRAy8bVkHM8Vny7QNz9mprWb5qWto28mYyN9HLaGcojouhBupfT
I1J2Fr3mUZcQotsh+DO9O9WLpeGSufRUoOqFCuj8tZkYYg2mIAWMkJZxNbfDn6O4mymCcdmSLdY0
IgWsaa0oA4LF4hiZJ68AXrLY77xclpCF3rVyo1wTWbrK9PmwuTv1IMrrFmUT701MQX6P4nLvlSXD
0V/pqLvCb0GDXNYf5r2Q8yij1ocyFJeivYrh2pqJw+Hbqbpp4CGNQMw0eBjlmfA6SLOE6s6nX6EU
CPheohWJeNtYDAbzf69a8zHUKM2IcU77vvgc3TV0hJXd+qBJYnxfl3wMY2IMsx/kWwNHWBMi76Fa
waDiI5Sxb+W7h6QkfL9XDyJEjjzM1TG6Cr0t1IW6XPk7gVN72HP5MWoS8yQ4Q/o5MWBCa0bwrDM3
g8BpG9kD3M0ndsdoz2PD/WwGm9kPoqghyliEwR+m2Ao5f0FEZE2kLJmlrEvj2gHxigXcqcMLoFcy
d74uErz6ZU2F39O8MvD4oDraKyl4orrjxEpBP6Tqas4I0jGFTCLluXUKZMTmPv7Ns2QbYP8gh/ip
CXvBAzVrCy7/b60FntHwmUCUp7uHKJ/ub3EkceqWTqrrV+XAL9cogp4fm11UzfhnIkhx1pBycsd8
9IqEBFZ9O3/tuFGGGW46RzgYogvQGBD39PaPHiUuonFzSGoOiU26GXx3tHxug788CSRGjAfRzkZD
VxaZ1iA2PdHP47kBXPoen0zjkCo3c+2PZElUVSL3/8n4Dw7CULUdtQUPHKc9mY6EY2PP8L5QE/ZO
nFBAgiVCWC5JXj+tHp23yq3PDlKGhXgbDDFP6hEhXUJ7KDaZv1orPBTtOlFYtIytZQC9YDjZ3/Er
d7miuyladNS5U36S1XexWS1ftSFXfM6tMC3b0RaIDM5o3dIy6moJUOJrKFVjo73YwtUSTTghI77G
hkpVF5wz8DTm5uHAdJy2qPN9AE1qu4tZzin7CGfDY+CCagThfyw/yEt0E54pw9KcpVoddUFPnlpL
+bs71czIRPtAc5FcCBRYYF259dWVAdLIRW/IXMgQ3NIWUHsAS92zoZcsZc3zi4Kay9vgiPeFv+W4
/kOv6k6OH23sQ1Xr79PGA5v3lBik17AiJo+1BzKVWMTdYwQXAep17ONNEDwdIqSARlAvDcvq8+Rp
fC8Q22NDFTvx15lavy4Hy7TjrLpi0tHSwokfvLEvh5N6dopNCg66lu5VDA6k9+A8Stk2tDFzYpE3
/dOqoc2rBAs9Ua1IXSAB3znfOcJG7CQkWoaF+GqtgbAzeJ8Q5JRGWXLtrN68CjJN6siK9LFZsFoN
2crgjJzOc4Fi5UzCQMJPlDGBeDfbtZ+N7/w/FACg/QHtnVqarLKfE8OqEp5fWz0PGSMUZAfX5h0Q
R5OwcKiX7iKiS7xQ755T8+mKKT0Tmy/PTRzjRz+tKxSz+2dN2VCMr9QAoZUZW0R6z74k7U6gY5Z8
YmRSOoc0qtnFS3VsFjaCvLo9ZmU4X2baOcgezirUV9FvjShACQzkCHGRDo7PxdT2X2DSNeL2ZdN1
QOHmejC0BnQ7hYUX6UWalB+L8CGiVAlDPFlZqJh9rM6uXfDv9FcTDaC9N3LwrL547+8nY8TaEmKt
zxWOk2epq9ShHqJMeRZ3DkHILrwPx3TqiWZkX3qXSBUxennT2IDlaQsBT3j+98LrCEphfDzaWRTR
O9Z+80MWfLMGQT31DU+jkIaq+LGH9uf+/qZgujJnb7u5PoVP8gp3Y3nN8tdRsxvnMc3+fffYhFAy
gFaz98OwLdiLBv9UeCYFimxNCQj3XB3vpI63HomRbScvjweLeotPo9mBffx7Eu8raWNNbhWJbaJz
xDM7I78L14hieLzZ5YHVoseg1QZ9CZbE8CqiWSWoZH9MZYcloiTJh8GB0wJb61jJSNKER8MQMtjd
uhpc1/QE6VJOJNbp/uTgHG3XCllyIVIQUjweni5Hewbnjc3YgPssCWr8IjZ/OB0JajVCfxyXlTDg
bQ4dF6xcMv2bZwo4MgrTP5FNWSCDJCqJgMFqXm8lCKdLq10pBGllD1bO8Q7sLU1NCj7AZ7gZD/Hp
oqAvHdtngRYlnVauwBN1EDn1WprrZA/v2aLL9q0v1n820a0JANygLs5I6QQqug4vAWvmiG155MXw
NA0gKhomwAxpkgcLHsBq9ik5QiD0qakx9zw06iCW18Irz0KEQnPS/+BkqP37dbiSNG5FTHG/CXO+
yLsV8qxCiK4+jMdHlJzt8INUW1eIvCsLtvr0+KeHw4T941Qxq9k4qdkJQ6q3alg1D/QU9GsWEL5T
0u+OTAvKVzbOP37WXHMLcD25HY72p6rqlSenWwxWYckuJyUkWu+jzKA7AY2lRjbmjunv6930cNbl
RCKke7B8gxkNfjRIe6xWHn0Z6w9tJEdb6jtZ7BriMEs5cQxRR2mDxbKeEbyDN5E8am+YJKtMFgBK
jSV4U2bruP79h3zJ0cKEO65D90ExFdRUZ6oW/exwq4IgKqhUCYtD4Q8tEaRtzfArAjHL0gEjboLX
pqtw/ZQoANA8rcPMCIKKGq6w7UNaPUiGcz77EZlmx5H5UW+fpogaRQCbfou2ZRVcWgVAuPjYEhzy
4p6LCgeQQzgORTkJFS0NzJYP7aKaWjLWgHJCB2LzWeCHf3MQbOqJAoEcsXB7PjhaVX3A3M3fYzDL
bYJ+MfVfOZ6aFYzIMPNWKrAZHGZ1K7kv1NScyStaPhU5hd6t3lXIda0pOs+/J+822mAO/r7tvgIj
Q0zM1Q5BxhMuVYoc32LB0MwWtEMa7lJnkJxcswdIG9iNYckBRezONUXxfgxDJV41gPTc8rLg5KBX
JaBTKQjMRdPWhi0tdYrGJu8dZqhbjcRyR4uOkx+9kYLfjj8l0iajGqRTKV+AoK80WC/1GU02fwNX
HF8rosajhYy6PenxlK2HIzYEAxRz5l9UpwWKy3wgVCl96Zq+y+0qnLugchedu2Nf1q/KLVvoMTa3
dD8Y9uzU3VKvBS+IsqpysaaYWsE8k29l6nSTYZaKJS7O0j2or8AiTwesuEDby6Vp4EdDBYCFUPEB
wWCHuu63iWk2chpg/2wZIFP7yYnEzKZDoXZMelJzUJDWcadve1SRrZpfF+uUvPZtndYMA24x5rhX
uttSjcyagxQq6OhhwN8+ac7ign+vEOBGXWmabA1vueQkUAbKvqpMbbDB/ZyKPY/XgPfOV4W24v9g
DKsOE+WVEmbVZr128mqa9cB06Ow9rGdPdLK2VnzFk8Ji3QOMfADv6ntrYoPJLQPv+Nt1tNfvza/I
wdUpWIq3IEZuqXOQFjZAH9tt2v0v5AnZriZmyN4SGymxoXNKFi2CUqQwCkYfOjW01htZ9HHtpTl/
8DVWTq1BbPGCiu8L/Qp68jDGXS7ga1VLmvVJLIxZeCnxJ7HoiahjDwLn6Mxku6ayVys2T0TShCxP
isRMU6BVdYbU+5v7VhnJb48Dsezxln6ttdhhKDoK7Ih24BUGUNTOX6fTmiUc1mkPmRMPdL0xTrCb
mnjklz01EIwg62unTrvNdcoq3mFQXOZceCHg9z1OGoEa++pWEU5dHxWndt5yEFVvwgd78TMqx65R
LlfBS75FaN3Q+usFT+vtGGGZQxsUODu5/qegfYWDtKjWHCG9GN9+6dzHWaJPFVklgvHn2KDRDQnp
sQxL4hDHijXZedamiwL5aXX/qV82Oa5YgtQ0nnm9l7hHsQtml7iu/FDIZhAtvp+kBKmUTIXMWZMc
yRqF9YYZD/WDy3hbNmtaXDTQiCyala4ni1XnlEIwBfzfh53U3mbHmbTOWzkclJGBY8Hm34RWPI1g
ZlpMLraMKrBx5scgyzboA0sWRs6EGV7yxULNYuXc9TB32dOs9/y3eeaNa1aq0/Il0lEnxAgSvwp3
prbnv/xVuc8tfhpwwa4elxxgyyoaoF/W4yPyYqrZwR8Ygd2clWJ3j45CDW2R+qj1d3o9hPrLtjhS
YmdauzfrOGh6KKGeE/cnok9fLbG4Fjh1YPg7Fe8hOUqBBN/p9m54fpj5hur40G8clU6YYhgB8+Tk
Grg/YG7Eqf/80NsAUg6LU0Ifmu0lYEGy673fiAgEBHAFbKJcn1LQTrtAgf8642ozHL9ji5gMQevf
PELyELvJE6EZVrCCIIFEwDZjkvNPEWejz/OSyUhg9YkyepLnPo41FTcbpTR2z517SHaNTR/8NI+b
IF4BN/slfGkgggMZeE+61dWJF9Y4OY1qyN8K2f9mppsN5D2YUJ7GZnq33UtDwTvKhbqkJJdOYSqP
3gnWpVjWzVd7/IAUIKIA0iazjHgtE629AyrLcEIebdRzFqCnpaU+8Peem87+WuOpVt+2Mywfpy1I
lHTsWRtfUgXJDhtSvQDqG1uzcBz1Zg5WW7aia7Wvmk/QT1Ru/RjOWt+lzNiq3omWWHrx4rjm8mlg
JmiL5rYcrK2HTPxqOMEBk/jOv0scIarYvxL3jdvmzVa8kHp0FqSmmGvIFrMPnP0dsYFlm0z6L8uZ
kT4Pg2G5Td2zfzeW8kJNQQ4taOn4CL8mCMDDtTX5h/+Jn0X3ABmWIqmLa9O2Bg/fxdoE4LlAZ++I
70fKmZ1piJ+v5MQ9Fa/iaOGipObZGBh/L2e8Tt0aIxP1EuxJeerXtzEfRy5fAt4W6HlYwe29BMDx
KKv8qWYWZskE4hQzea/wRknmPCtnhhpppnatZA6R8NiDy1Jmt4u9pHs4pFYCuiL+cS7MMW7wRGcs
c9tElogOTNzNnSnL4TRlweXoSaUhnB475vSqElalyUzT7yVC/YNjmh9KNZtXqyBzy6tQiSSusyOc
RAZ8Z3AcUeuOR61SHKhpKX+7D25p1nPppxd5fzDl3lqw/vb66/RPAbmVIOT7klflEBwbe7fADhR9
0F6RvlTQ6cs1Z1+l+SK5kk9VdsrVvgXxVCrpvdcG4n5YvtVoxCRXGG3/2CXLwANMTXWZFS1WERtv
TRMQ3XvPUb8E50TceEWkMM61nKSTIDErHOdjKgL9I28v7MhAEx5dICzn/2ZHI2tluSjeSmyb/SwB
ZAFrvA48a23Ju5+sOwvzUAFGy2rMC6KgNRRx76TwbS6/AScTN03Ior+S7rGckryYKfUM7oxMLWvp
roS8avw7HD5eA9ZTF81uMdbO0yHIlL/7NtRm6kC9YY1ETIdbEf0kj8g+anz81rObnhMCpY/THBo2
+ZwJHMGGvVIwD+ucjoPIXDuUG0cAc3aFxu8gBK394T9A6Kk3vMJ/5p5RDl7S/GCXCfsVI3VxktN9
OuMn0wKKGgUwcxZChKNGAMHxqUq1Bix3nsjSf/uF1kFBijtV/ffpLIt/HikquYNIWDcF9R6YuwSq
oRq9cR3o6vAZh77quijE61UHgB3NPI4MFi7Xh95lRj4lCkWIqrzV/LLg3OUrPGngAhhuts/piVXz
2o/tD2hlsukzFPSZegwo/SszIlqRBN5dIPffBIpwAKM9ViKGfKYHhYVfWQTO1Z1kdXRU/328x8x1
yB9gg7aB8kkOUbouDmToBB6LgXHeA9N5i85MEHzo1XvBtiGTWZ30xV8tlW4RgsGRkfyzmFMcjjhW
Pxin08LO0Br4+w367ihWyGP73SxyTsYXBV75NPcVMwMWUUU6zrmap5Phvpx/SjUD9xEGG4mKyibi
7sKTf3Wd/QDLTtjaIYqogXKzeI8UrSuu7Pa5PWr6xjK5dikWWf8q/I7sG+V2qL9EykF1TEheRmpk
hJ+XI82QB+Xty/wrYzTnKygpOJhfzGyOjugTTUe8gp1+Bm1R5sKriBmgrt4t6nbDep6nTIo1HcmH
t1qzC+5TpMXOfLrZBZPcuKhd6fKJ01uD3pWu8vLN6AL4uXSKv8m1ryGJoZOLBLSsokdV+OE0ntxz
Ew9hVHANfpKtoV0KT1imz9vKUtm2/Hql4AhutHoAE8NYyq1FBpzV8RR6igFsv4jVAWoKEMDdZBCx
wEhTksHK0Y7vX9vdTGhaCXLfsQoLQ2Zw6rhDfzXI3yWrCYHO79shJpQfOxI8Am3XNsn3pdMcdVCD
52VEqbOYBbYuSoF4FvJXNbcx4xnwveqZrr31LRvcWlpz39TL4e7qCO0AuAtoMV/h/e+6KtLqSEGA
rxqRb+vNJ/nPA8J7UoGtp80BdJu5op6727W48lPE38Rr2ZEXZJrwQCN2GHejBsjWDXARRQKgQlSN
fajuLI1SNZfVYAE2vWt+5zGpwJq3yn+00bTq+UYB7G+IXjNKVstOAbcrLtAcx07NiJN1CAaJ2+zi
7jUY0iVwI5T2Ph4poK4NgxTfnlFD+o/Ta1iqMh13ZxksXYUPoPp6N+avnh/VI7MmWvLrT3dmdt1H
FJcHOtZ24LYdr/HTkTPP2P1HCBkQiT66F7vzvZhap8kb7cfixiJRcp3ZAJCPKX5L9PC/8W3OufW/
IYPEazbAulWSrdV6h+xmz3imzMkcU2owic5M+SYG5+pK3WuNJKSdHbb2PLlrJAC9VFRVGXyaM0YJ
iggSjeDKACyQhZ1ehFAHtG3ecjydJWTeCSqsGeelNgrvrk97BnUjPdHEATcdpmn5ZMcKv64fATIN
FGTUypfUgektFqaUvDOMKMsNRxYBilV9SXNhtfQ2yhJi5Pame7se/KyRGRCH7ZhXWu1BGJj5Cz+Z
8FJH6nFFs5d4K68TNxRH8ZNRV0T/CdRlb+L3oTI/5bfcZMmHS5F+7WhCQcVXX7xn+P5mP1Ch50Rc
gZ9AH4PnSSrEr71+Rr+ZbqDb0wybhMSy1K94TCBeWsC6rEaAbYQp9TJdO0b611sMhRGcXq00niSX
K4YM0jeSFtYVsvLSDRMoUfmCYBlIxdcZBS70bbSXnc3c5lPw3iuLhgCJFBNV4iI7ZREOAGSrorYN
p9TK1dqlzblltOm+w6wTDlAIXePHzck8bku6Ig31/0x1BAlVCBFx1wEinfxy8h+LxHDwOJGoHDzQ
eytkYBWYbPVvHsWcnjPLmeUHnZbc9fmixTAPBNRhR4WaAgS9bJtCHE+N6+wdI7iVkz81kGa+AQXo
VDRrY4n1yzPvjoEh6/zvX3RP0vEGaNjPrk5DcAUHJk1WaeQQPP7ZxHrrg1mAjskc+WyKjhMM7wJu
ueNbblBHl+0TifXrz192iQlmWhrsDSfWyuxTTCO0Te1HB3QDqq2uhXKF2ceeOKt3GhvWJ8yA6GaM
W5ekgqM9gU1+V+xAJSi/7s17nJ0UN4xD+wqChAkp979LmObh2+s5SMOh8fG1I8eVupsnL9krqPV8
Nb74jhiUP2HlCWsEWY3XDxYG7b3e5/+5Cos1hoMQQhca+C3nTEEwO2ALNmCCzwbklc5LFQXbN8EL
Nb21suf4nxoa3bHq503pQvyOHo6r+24ffTeNImeYpiLFGB+8IeW+a6Ez7q3AGXyoSNOgAD2JIjNd
uHupB2YzJvCe3/sE/5Lq7KI7hUd3GXo54Bhw+EftX96BKfceO3VkuYBRf3Mu6quL1L5ViO8tIm9a
roedYmesLegHAzwp9jun7POMBGfEZqoDmNR0ADQDUK9eXPlc5FBZ1NINNMM0yAAEA3SGg5DKAcVP
kqmmwKQW4T/Pu/ifyz6HdXzA/p5XL5oaR+1SeZT/Cf6rGMrH+Vtwu4lRzJi1V8MQdbsx2n0H2urr
tLNawpqtgshw+kSgX8BxcprsovD8fXmT6r7nS5vj0U9nrKxkNzmc8VqT/CR4kabzJ7PFFUELruWp
mxn57NRsQGNIBghAveEbm8hWQJBByfExwB2xTdUz42yawbD0GN3VO9QzaiFzLsEaXnGYVT018uS7
PwO3KfOcYt9CTE+vE2ni4EtSvUUoFEtrHggPSGRfilLM/d7SIf/qhPqUQf32Q/ILKoLVOW9ivsGD
Qr4RGzjWdA8eHSS2TyERrToe5ptw11mprD5PuKXsK9yzJQJuqJyEEJm05RxLmSU55ldSxaoGv9SL
uku4vOSzyVID739wmMIf5wC1N6cGy+1bqVZWWG5JDfty8Ev22plPycvZrOY4iTK8z7wKHM2yQ57i
aE/v8OX0zDidNs6duAsr3I1nnhxDxIiJ7pdBbfWiM7kd77QI1/ltgOj175eNXWXFG6j3TiF+s6DX
Vv6d3uzqvrrCLHVkUCqsAyX0zyOem8cal5UkRSwaSjFOBvjs83k45ztP3HqLfXwObPlPojiCRD0Y
K9jVdToHE52esyt+yUdiIv/m3s724iupoSwttoA6v06oCJ0cixN4K/tJBdqKl0/snK1FuArS0ERD
MCEn8t4vuhp8o9TFu47ERrZbGnkXnXi6kZ/19uJvHB+wKnuWAY/rYNJ+7uRodeQwN0f850rpNZ9T
oBMm0MzvjaKn7peV6eA/+lMRdmmPI0vVfg/iZLu/JApYP8IxQka7w604bluuuWy9IHZbcfMTkOnd
VMp7VXcR7f+hpnbZeW/9i5UtD4O4Hm3Zpic49CkPHkkLYq/I02QnNmyBUOYs7hY0hLWTAUJAa/V/
MKzhi1kL9zLDxVqyPpO/LzzGdfnkzdhfjzJtnWCUwtGqto4OzdgCXX8soZQaFNUYJPOwzDARYI4E
8u3XrCnwl141saWCQOLyPAdJshpigj1InIMWpJ2FBJB7hIcFh8XHtcnmq7Zn2mnu2TtIcFaHOVpL
QSt27LU4iW0MEJGLWx6epL6YeyQGCQPxOscbVLjoiIWSNPIp1C9mDc/r/7JIIEw1jGXDY31bbw7Z
Cmd4lQ1v9RVJo7X0cFBXmiZmZW8yw4dvD58J0se9VMCaz/jv0QoU+NyodQjlvehGd6iXJgHRphRY
v6woIof9TzqoytrYOGCdOvsSN3uFy/mspvUt6QN+1LWXhBzgAOcRM8dTLU+Rz28nqdf6vkHw+qGm
69c/zoOLOlXIU0xLs8ykdTDfPz4isj0YsbWyBGK7JXyyXKhUD8U9r37uSN5uz//Eoa7oBg3m1kDt
dcTNtLKvyRdn9DsZshcuHQ/i1j4djaGrqdy9SlaEsVkBHgd0D9pO1TgUUtML9+fZbIrdhFFTylM8
hZp/+rosKJYaQ1yYUCdcDToWQcs3577HQDHuv/yy+vMnI/gNLJfkI4m+QldV5FFjkoLJPW61WPZB
GxkDoCulxmcRaN5uJKP8Rtsq2hogNwA6idii13u9XY8mHHzWzo+DbMD5bxAbPYaByIdqFbtq183A
gCoouceDEokflpy8rlX3zC3y8SzFbGK0vy7ARMpa1Vjzc+5nwJmexouP5wcfdvCgF73DVbxSrU3S
mM9kr+v1rsT0ILI+eu78sYaW/Y50QnoImnf8z2LtY1nTJ+nlpFTGIf1V/IDIH+udtnkB5TLHiK07
lJufnBDQYu/kXrzYhIcW6oYWZeJXT99NTCOAJwTWuCY9HHAuCAg3l9uHR5qJ7cxG+Sc2Wu7utU6D
iAtWlhnuJVmZ8b2getoLP46TzujKRXOKFoDmmVclg9IpUof7HIH0A++4fkdvHlYGLy+/0Xf6jTLC
OsGunlVSbzPHMixi0N2p/80wj8BrTV9icxmp7yXkhtPhEkvfxHc39ySo810qA4ADwSyqsI/xZhyV
2CVCE0Ujs5mii4/sr6tMpz9W+rXBBA5niNiLODore/e1AqF34lDVPU70IBfhBWTufFYVpNnt25dZ
wUWje7MqNz+85HHy56BwgjC+uZfZ/mvPszCNJAMhYGJarMhK/uOZ2TTIelcX1An/IsRdxLZmR8RP
6gmh4BJZz70bhwxVIJIfiOvF9o4cjJHL3JLkFRRc38ji8IbJhiY40J7h4+KDP8eI4Ttf759UwChL
twXg+RHCbSRMozSRPztS/3E5qfYohqN7c1FU3Hoj+AXAYpk36Vls6Bko73Tlr/41VA+akMSQ+qgH
x/asscsjDm+xlrRnJoM/WKMUOU/b9uoYj0jTXhXQhs1OxLXDRLjkgXv/239+L75XBYGMtMbYdJGd
fgegHyotWNiNGxrdWgm4jepWIMusEWqq7XdAsS5nipzo614ichaIdx8O4LHaiyBk0AQlPCkAIuFL
R0KJTPjkfqd8cZS1k7d4hOX6mxn/BCXaNeopZOOHG5jj4r/picCd85WgGX8hGYDwsZWkrWZN0wBl
f/IMWz0eWswCcRB5i5obN0KMJpJl6C2c2O02UH5z8ExFz7/YZtDSGAuQeSAxmbL/uFcbiO45NAHM
vluZ2fmGyXwKmFQYBLEUspzKeNfni53UB1dxovlLrSjBZCYV/CLDB5mTB0FgsL3Gb1x4QA3zArkO
rZgm0hEKPNFkocyap9XWOmXw9H5iXo3Y+9AX8guK4HKqVlUhlPTSf3NfwnFnyB+RY9AqAwkArBeL
SlYg+4FNpxKhqGwCVCDe8P24CGvs1F7u7a57cLJBl8i+t+ndzG3DXZtjgvfUbRcpaE8/zBCCZn7T
bk8bLYFKsIn6akAyPrnEYnUn1U+nHFR6LszYhdzCDh2OrpN4MrYCQLFKOoH7fsPlWmly8eHHZLFz
gGq6dfiTMw3qj4NZlmMFsHfXpByqhPbtFpdF2KpTr/CPb6wht7JiAGG1+5C7xM0Vq76BjOY2AooJ
8lfSSaz2eEO1d5EV8ATYZAofK6yyoSuvwuFYJrlCwCLHlhaZY6gKPUuNPhpdiE9VBTIU5zGB4N9l
SmKyemfG7CQS2Oc0YBdbwU3zoE9lh9N81vMtXvUbVXv3qbnEunDm0xseRP4Mdi5BAy5xhvG+qEVQ
4gUO1j2Ck2sl5K6t4QgxYy/0p8Ln0BYWXdRXzhxO95g1gpcXCoon6VtyLUvztKL04MN9VG6xlXhZ
UurzgWhIthHyMVVpXe7ueSVXfWQzyteu5FnzVF+EIq9JWQWD5ajL7ZXfaYMTYyMJMKXmUwA1hOGd
KefUp0rQoYVCDV+FtpWn1/uhQxU86zATR/uMdoYC67IjNfLZgTFR7a7uKw+JBYg4YkceurGKaXD4
1l+dNCTvg2gNEyhvOlT3kaFaL+GwVgSo6Pm6x0c/B6YWTCW24t4RNv/mu3tvMOtVVoq/3qjFiBUl
wn8w0a72lFkDnEHKuHPNwJapiboFhOpStZpI11utSiVS8KM3+MzhBs0eISQcP0yU0Jk1fJ8PTxSX
5lcm7DUeTMn8pPnPSRqWKsTlRCjtujQtkDXkM2jMtSD5Bpdh9TlHq2Opldfcg1OGC3WNENTVTq1k
5hE1fdPfav2FGy6IIrv5RXmDobKFNyzUcPLvKYTpnMVrCrZrIhMIiDwcedr2iSZWhA+Qm8WpMONu
lkFrr5yXZQjmaQBUjl06Z0kQ7BK75IWg3cNtc6ydeXgp+x19eSJBpBwdkXgVHXNXHrAuKlSbpdP5
Omhsy0PMFQ1DZNTrDbGD27hMJi/n5BlKBFJOpkFxn60wI5KP3oSElCwR3cLYyx48uG3H9V4vrkmg
OXCH4QY2wEejug2WbTvQ7AccPDNOurI+IYiRdrLW2UyDoh8tEvi6MxB+p96njWBMvlYzU41HJUJE
oJFD1l+jIzHmmsMk/9BYI6rRLvnnnVrnrtYS+O5dBR8Q0/5T7Z3P6ZYdfH9HiEJgkXVkXRbbBysZ
+8QPGQdYEhDIm5d0i9LuxuViSryr067x+rOTkcFjfvFtt5RjdWO4UIKiP8OQ/VXqUUtWEeNosZfS
sHcc74WlACqIDUSVHHFiruFo8rrvXbjYq+Jik4sIXgwYK1t6tJXZbV8GjL8lMH8D5OoznmntS2Jy
4FnNGjRNPJqYfQUowdry6SwTYxDCe5IfAIFLEd2M9mm3BT9Bsvlrqbw2hezbftUAPRzD8kd4wkq8
QRP1IQn+Z4ATmzHZjUQRbqoRvGCUzb7RSHlGR79FMy7a7izNzO5hN1VCOHBowGrdJrJOewj70EdQ
IZfLEJ2NW82H25x143WxFPYyQU/IfD+Q5qdVBjb9spurwGzc/DmKSSW7Urj7HLhzrHnj7TXBcFaO
TWEJyTyEwuSIxVIMcuLSMy+fSZk8efHCTH+acSpy05wUqNwiFbBvty9lUOkCbv3sMd+cPsyeiPgG
Kt7WKsgmZuQJUrP/2fIEpWEdorUY/mGEpe3Bd5jGiFmvcorJrXXz7RkLrjmAtPjSvN5kgensBNbu
/hDD4D51RV5gnXG+3Hha0PBhFYRR1RmlGuJ57XFk6SVdl9PPUyr+GdxoEXO6peSR228vC1u4v/TQ
FOKQqwXkFM238o5iUbqQ/auwtAuw8ixdgNNBDemUU1rA6qbL62ddwC38ucksrWGwYvWSvFK71B3Y
zIMoE49CyycqZI8InBF3InqTJ+Rw3dUMFIej9aGyh44rUa/IXldix4jZPKvLhRl9T+jZUujdPwIg
qNgG3K07AT28CotuljN7P+fHZQ+0ZfZ1LxUQRTGXaU6XYISl/b4baVx7ETKXysUTdOba4vVC5o8R
G1plHzp/VmtAllRgreOon4i0hHquDDX6+T7/58RIzQABTnRJQnM1FPonCEkVRky+8mda+8dU6IU1
IyQm3nPOHO6eqBs2hiBOzAvHy+9yG27VEXuIj8o3CjFERnd4qvxg/Jxc0+46noHx4QtNO686sJSk
6wZWPKOaNni93Lpyvhoym7ToNh8AvOFTfAmQSLUwjGgG4KWGcfPtscwl0J0AHdG92iUlyQLE7R3N
BlL9MwvlnTqOQgYxWntfYMni30xKZF6wwNyLIzUUYQZtRGLjXEpyr7XGTfddM/wEmrJ0pcP5B1Nn
EgOC7fWtxPZkHmuUs8Xwp8cwDBULzfc+szB7O+pr4gUlBmynJyeWSaKlua1SZ5TXruCnThQMjmzH
fc9JD+xQTIvJE2HpGTqj0GwZSbePApkuZpt1Y/lPAxsgC5aDP2ATaVtdr7X7B8wqVoa4MauZpGkB
MxJ54DkNKS21RFYVj0WNeg5AicfUq0bly9Sry3xxH+3A4iTIBf9vlE2zxwHAWqb+NTeBxHSZtsVo
KoKkZ7ASNwB8F+ufwWJ241YA8DuWZHCepJv+AAQq9/hJidr9dkDQbAT+t7uSvfiKoxXZZ0bqUo3F
stN5QdH3h7Kyd2VDvVMcPNug3Cjb4VKEP8+C2OyMwDr5tVuq7RCUzp0gJThvIp4JXzZ+9U7Y4uRr
bkjKDsd1w4DY0zYaMT1Vnnpx9mhT78jOh2k+3XuOAmkekQGPgJ9J2ss2fb788Ss2WbyrhvcB8wZS
LCaMAdzYH89WcWAKdUtILD9SLKGm9LZrxgUb+t7Dum1lsDupvTIlJ1EkCEhUvsDrT5/lJTSdzO/B
Lh6f8LGNSsqFmcqEYvyrhY93D+1r7PHTGXXQdAA9eUjpu+G+1v/Ubr6u7oXE1pX0BhKBT1vBD6Z5
q23/h48LfzQdaBu9Hgvei6zujlnNNM0TGoVsaxXRLmr4yfQu/aN4wQylVaaUuhDskAq2VCSEWNtm
nUjy7Rft7mt+5/pyOtAXSsIc7YartJH5zQ+85P2I4HZVEvGsBg9LoFK7FgZjuvv37hJRnwB7j/dA
gdJYXRhVWr8UqPmKNpsvLU055m9Iylw4tmh8J27Zmg35mjPxuWpJ64MP/4z7h7A/uuOMDuAmLPm4
A0ZB6fsUj/U8/3BOhcsWjT/7TvuKUKp73qcwLXOu3FaLEPbCGxmR+cvTZYgigyNk5mYB5vxUz3J7
B8cpJNGvb2nvBfcCDTuLKdtLnnqVlLpZ19oy3033iWIwlpqTP6e/4ge2pqjiVCS6sz4MaLBe3KmS
mLI+AFuSSVHKAmESuJoT/rsSy24S3ZKBjJdK4NeWUITsk5dOmeO4Lle++Wva7QG2Ixkfvqb2ulFc
98PT7eDMitqHpc063/j9h8iCRk1QN6iMmuetBWj5nbqSmXrVU/+3l/c+RiUMSQVH6MOWv9Jwrv/d
pzbhl9rV9zzl9uUXLqCNQNW+R3YAGp/P5lLdB7Hvf+CnlBhkknHP0MESvlVlfRWDu1G/ViiMh1ii
GjdsOz6WvMqcWVzgsXbbxpm68PuJG31MDaSfqjIa/uudEYjbIBCYBybllmCqcHVFwHBK4JVlUUE5
0dwNHVByHPAu/BHv4bVGBMfpUZIAOnrklHyB3hi/rbZ7nwwk8PW2R009xsq3FqxLkwtYq4aMOdad
B4MkB2GQs+Y9uibSUKJ47F1PZhO9RjSnC+Z6V2wZ/H42GsEde78edLdc2xhDZPnEapbjjv44riob
AkATZHxv2Epe0UzXU87j8JRCUPYl0dC58a2CH5vPbcaX81up2VTP5dxs9IJUA71SU0o3BO6GgMU4
7VyPJSFB9vtgMLI6lEsnq8rJiN+rsnNEJwNrnD8j5v9EjlRux2ZVGL4fgu9y99AO2kdJ+3mUMzsf
OvMxQ/P4d3/yHjYoeSQrh7uviwzbO8VuVSpJoJDIoQdS41zdN3LL4DBy25Xi2RAEdjunLi3KC273
Zv4cfWYBjBHBqdejKDy9uOsz8Cx8TuXe9NkQOaQySgbCu3bfZGsN1FxHgBd2ORa6BNKaX/9YA5EU
7Bz3ncguy5I6VHVn3Oux0ta7YugeecsLhCam8CtYfgbS7e/GrXSFK7zDC5jQQ9wkjF+KWv/p1W85
YJRm86nZyyDWZn8rgBDzZeTf0Fm5IwEu6uoa1NOFzZOncv1Q+bXKc4c5XWjCK8Ap8JhsYS8xPSJE
xCzdbkLmy1Cd8rjeN9040lwYzggB4bzt6fgwER/m2Fc/DcuUNTGWpT224FmloRZVe1gmZfnlfGs/
ezW/XW8MGCsnhD72fuq9W4VvYXogBUuFWRAjh+M5Bt3+dMr4PQ/jDoOSbFB5NdrG1HaeqRKVk62Q
dq83rzsPT9ZVSmpN6Urf9L+2OU4wUmfRf92VCfurOiqidqmvVn8us2Wa51cX9AuVQN1EUYcks/u8
GZSIHfuT5X2hrUbSNKigbobUT3Uqr5fSXeyiYn1dxu6dk18yV7qKLhOiIuxm77/2B5gGPLdv4X04
46XpgSltb3LzyH8xNpzvCORwoq2A92v343nuKhtqalcpNUxwHCqu9HB6mRVIvGMAs4wUbKxIMGWp
CEPG4CxW7zWrHUtyIvWTfTFrHfFJyI6VeJZK+gYgcpkfuaIzen81eW0iiqddDs6iN+Znq1nnS8sD
gm2pK2pZg3EzdNaevdJ9h6rx8wKrtANHv367Uzvrc8sNX8zhH2OgXjzhaSllmiN0kHYdWpi60rBD
MZNhMPBPTX2a42UmYtSfMD5yc6BQy3qD6gQXaKXijGZvfwY2tY1o8Zrq7czUApo7afECJP1fGniE
eZM86tI7p4QJd2b77keF1Nv6I9zEjr2gC/roQC0eeAF9rlUVvxVjPkWhFYbnrKC7l50qCDoutkez
SRaJiRhED3k1F11jsunEnwtZ+x2beaLKK5DMU10pI92SaWx92wgce6rTVenOoiTvmZmq+4vRSaz0
f763JZ+JG8inj3yX0VM6zDpNt2PwfGTtC77cQ5XrTp9kzbResDKZHXyXsKb3nSbRjcAeF7iD5QOJ
tFOj5Wh4gLB2SjM8wAheWf50cwXcNqksTItpWeKrWMpdPvfF5w1jWM8FLrqQOjIIFsxTaHXeR44S
z7x3UaMdWiULk5CIVmWP6NfwyNODsYxO5F4bd32+m/iYsoolmAPkxbsfxjaSjJos89ej8pdfcT0g
rlDpbB+7Foy01f2dVqN7mzk6GJLKWBOVqEt35gMMYiaNA3H1vmuMuyylAIfpecphb799FRNz0bCk
hkAxwxOvBZ3bNy/Exj8VlCJhCmF75jEnJLYNfJAsIjcEcIieGvpiMfmyTzZ6tamIvmXYWLWxpzz4
NEG8r7lRMIrdawjNkYlS2D0wgR0rMIYMkVFW/+oFeujpmSP9gN+NFrLfs+yxy8SR0CFrVNpV3OKY
iMnBbCsAIxXsP7zyYCe3o42Bn5rj3FS9xdaZJbrnnrYlULC680DQjtNfE0hCRUj/ZGJ9RP1cYKTJ
qDq9IJy6xiEsFeyACloYK0eZ7ozje+jCKEuc6RTSqyPcmuGhLUHg5Z7M00UjZCxUNTL84KtUnREV
9LHpa9eDhSlghdu1rvdpcsdOCvNQk4b5jkJtQn6qnzY8qV+kWmF2DBfif5ELVbycnjiKVbwHsLn5
m6CvOLBs8B3+hEyq9MHFyx4N32933UXVeCYYs/goGlWkHt9g0FXDZODKhEf7Lc3rVxzO7xMtDTAm
wSfPoRRlOzWNLxWe9gEDomBvwvDIWsCLTGnIDiHhJeB76HH9hkfRE2Lch6JDuThYVDcN246w6yRP
Fo+a4uvpkRQMSczqYW1zwFGB0sN0xzlrpn1Gp+0AO1cscJ1AurVBq6bDYk5MyaaYrTZrRitlaEbJ
wbFpFNqwD/B1xX5tB8bEZ+xsE1VWWVz6dV6fr7Y78jRZH1L60Iy2wtArv1sSKjWwNOJ2cUSmIif6
RmrJX6lPtRQm6xGTpsUoTTCTXpBeiYio5uFTduOb4WeSqWncCv8dB18B5HAeg53TT2YbRfkw3tAP
Opgo6r3jAcoS1ZPh+qYbUH2o9h6KF1T6GkEna2me4gtoZEHG4JHL08nPnqz6zhEJ6832GDTXxDA1
MtJumK6tBmNoDKsXuA3iX4+C37hgZDMb56vOedGQ/ryzIqCKDjAD7TFCm8X7SO20S5a6xtWEU5ha
hEdGv+8DFlpiReHINPbtXjg1eYaTYi8ZxLr7gR2eNmTTeH7iU2g98MprkA0JN6LyTVvGiLLgx97K
2JN5b3wdXyT6kT8MHWmeeKcDYOAWWXafTkE4913UN3p/L9mABEpRjSIIbDZaDDgJqqLGTbmN9eE8
7wHEZViBMeVNLKf2eF5g7MaGvRud9U5tPBHIDvC95On20latyJc5Tw3URe+FwhSlBYmMGt2Rav+e
V/JfdHXdHVHqBAZckR8d/cpfuTI2PCZvK3Vx+SoQLLDkGX4k81RPg9Mq7UsOIW3PGld4sz1L1gO3
yFjRQg2YuckZmXtpsomNr8OoHOMRvt7H+MfxCimx3Uh8YC7cutpdBCB+w4ZqAnso0f+MP2cqU0eu
MKspslWOiUfKZkmVNnba/ZINfuYfxlqcNCUVLg06EG2K24mme839YwngeKW/DSnj7ba8EK2qFIiZ
PR2R2tf2BDjpgA/RRD17XRGxvJjhJbNoMe2cBkZMdEj5+wtBygbx0bO/iIQ4eBNm33VBlGn7ljxf
exdtgzGiW9xLZODuQgM7gjvHcHfHAuWgXOPkxSo2La5txwWd1wuo5crs/02MDiePtK+avntAr2v/
HlielqMnxcTNz0Ia4twe09O2su24u69ZZegpUUVMP5x6K4yaHwouMIzMCigkeRvYqAreDmmjRgps
NTZz/9Sbbk+33DFhPmdPZmPpYl0xxq9XlJIWITK+egU1nARDVJ2gGTrt3Jt2CzqVlGTIPjZ6fi1B
7DoTzBTX8IJk6vKdUOmfKdr/o7Sn+mWTzwHkARaSBwbXMzfx9jq7bedV14h5+q9vmcusEGodinCC
uC0cDz4OUo0woca8fgqnSjw218I+WCr8uniY3MVbiAMJNHWLWfRs9iXxXHkISWUQQFX/CuiC7Fqb
HpY2ghMXuVJrjjCUvDaBfDtwNj7b63YpPnG8u50A1Wn+IFURAnRH+vrj9s+jZD9CTvaqAQ+3DXMM
XoEofKOLKLlDr08mSQvblXKah8i0WN5yXXQliVjtJ8Wk+bUDWeU1BMQRAaNafEXZPnMoCNiPyPpA
AhMxLQhbxmryBeFCgCsZT4azhEM39eHD7kqxJEr596Sih2dn8AzS1SNVary8l3Qcni0I/XblAbHB
rC2Gt6z2y8Yuqml+Hu8B0VszDZ1cSMaryUG78c/sKFppd4MyhObK3Ksns0eGSrO95DJ1fg+vnHbR
ffTCiFWZ/xqdCAzg1ccUvy5p3irceuFw/Qw+jgCrwetyE9N6tvcqNav9UM27v2cMpACnmiIfjdlr
Xi9XLdExGbUqbxHZNEWMYmQZjqYHqFMPFeJg3gll+UngJy1R6kekxPA4oMg+yd9/HDSa1P9jyPyp
aNoLwYcBI7ve3XNZjFp9tZx5tN4TUTqd16l4pThAhJ/pOS8IVDgZXcqY9DL/1yKH+6yiG8E0d+bT
CKP7c5qxM+AhUQgscKYZQdoBjBAUioWm3eNJz0ozLpXhiPQmQ9vfajNhUIz4zHi/e5W8Df8MKlaY
/v0oO457/bk5qM1oWVvAyZfDE4KRLYbSYm0lvcFmFYvdYhYKZu2Qv+8KcbXCdcHbM8abwXTIUWRd
bE5To3JYiK5uD8fWwFIFAd69tr3kBJgDX0cTABBQxA4T3BmCyHJ5bVVRhVFmhdg49du3MtM43Clr
qC0X2oIZHP3zGbanqEKgvGh2QeHZrBscFP7R9AI0+BHwfCwJQpMDKRwSRZE7RVrEtX9FL9XBaWvH
pBujUcNpATQj+lweXFuk1etineZ3aQHW1GFp9K7nR1gB0//91wv1SWFmLNB0akO/uzlW4TwbiY35
NF5D9cKK030t7GVHOY1KsHa+BqK+jE8bHw3l1C0jZKPBSVt2y24RCRRn+2yrErYJVS+RT3Jr3bUj
UqH7zEtP63+QsWrULpZaP8U86hfmoTRVYdT0rGD8yu0YdGFFEfWPhryQ5wU15Hbn87AJQkQtiyJa
kWgZEsqxQHz+Rf8SVTlbYXT2U87UDKqPHRs+d1kv++tK5VZq2MDqJ+zYzW6byPgbnOGWCNn9Cb+c
A7vKRLG/FiB4kOlf2Ne1DYyS+UdYb47TH550pManaGnw0XM9uo//MQdzVoLwtaQIgH2/4wAxyYc2
h5cz3v+brxSM+tbUnDiPw8+6MYJrqsAPS5DNi0DfpavRVjKbv42mU6Kj7nk59xAt8B041tp2j0bA
2oe/cJX6/T5/iGEVAeq3mQmU4Hx2XYfWeXld++wEeZaL7BeTY/byHhacBMjlDsS5Kk6y5PfFzyxK
QoGjQpfFBmmg8/4BqGBgcrGCIzR54vyHoHQZ+G7KyQ2D4VFj8fYNe2+MitlPVFztBQXEYCS6AbMF
NVPtGTtHd+o3F+isFbbHMt+5xeC9b2iYjZtMgGWVTYbi5yTkxIb3MF4qmGl8/e2ufMfkGXJeAXNd
179r29gkc6cenFQikfsjY8hPqIcb7/lxW1uIUqsVbuhq6AhoWXAXtV8aoOcO+cxmBdNCFMwlT8wZ
Rh79JqBCy0nXhIIxkYm++qCdnh6CA2UJ8bdkJfQx/0vG/n48D7NuO4b5wSF01E9GHziJWPCRJIX9
o+WIxaU7Z3hmdKEm5fL27HZ7cz4/eV0qahtaiMpBCUm3NyEmah5V7/Qkb/sfsNMtlCGRVAd5k8uj
fkBXXh41jPzQWoJsERWcLPSkp+Q8RpyHKobuo+BGV9O/A5BLycyy4MMcba4/Tm3dO4Itbv28GLxw
jvk+1xgb39IQMj3mZ24WMd3xUor7TAhs/3gbZ/MB5lhyypJe3vLo0ZZKh90cdQ8INsVF+a20En/C
zPPTnnmSX5Uu8dCIVHBKT9gMqN/eGSYh9Hp+79abSjCem4s5vK86wWnNnfI9vazb580Ia3qkrObW
0UjA15jikg2wFVhYhgh2O2XiasEpEo9bCCVsvD2hpeiApCyqmWTopFwYlcyC4a1GuYSniFrCa8H/
BXHy6GMWgCfWjegoN+c+3AVWEWQISuYmHnEzoyucj1zjiopKdAcUDVBjeBU6KY5jHajsMqns7v8e
a5LB/OSWlWtcGI8yv5EE11q/YuEjeaFE4aI6XYtH/PxwtTFEYiFKeKpGc/Ut5JgOc1Rb6VHDR1D3
DckQsssNoUaKqfrjsGO/5aZAmu1iyOGj/vJiSa+wZnjBAv2MXPVU+DEY6kEDz92vdlWRkOm1RW+Q
C6S/ngKjx0RUHOUdMBVa4qcYJi2vDSgxFtvhj+JhC9q0GVN1G75GlmNM+l7VF6PIzo9DQCILLwSW
bGcM7Y55371fBQbkj2MC3k8/rTaqJoEUhFoFzzuINu7q6B4fVZt7lMLjpp/ToDxg4YQMACgg9Jah
3+cFwBxG4ZRxvFkD+B3ChTo858KnUD+UNi3SYcCQ0TDDY7CmgnQvoY8qg4LAPXAKNqJyB7ZGqFwo
UGOZfyVgmPKG6iNf+apq89ySqEDbCCFHCkmVzLc56KkNU2A0Xn8CQ0bahjcr9obfbyuMyhmFS6/V
4U6yLP2+XZQdH1VnbLpxuPB2Y+ieiN/qJciceNLsCG9ZVa8EM3Y4WbTcwf+JILiAUWj+jx9KShjF
rw4Qgl/g0/eD7kIh+gmTG2vGYUCxwj8+2pzkIPvTb/Y1MNea7LQn9cljgqHp80suWKNwgXCJIJ+2
uySukY3dq4pxPN5Hh09E9RhK0XmUSNm3Hzzlw6SBq88MLJdzbynJ/elYV2OPxZKXyjPUYX286x+k
WvsipjOUsyb8r4zBXetRgiCK4eVnEwPb1IIilVLcxtjkIR8hKBlKQ0Fp/vpJ1ZOfRKzXjg5lLnWl
w7ruFuCq+udxWIa/t8I8FdV7eZXptW7MIG5xbnv2sTJo6KmxxIjoOuzEOs70Q89igHsbiJwXrN7E
/drZS/qeZEnqIaN5jUqSRVbeqSPko6yXAg6+PXLhxLiVmqonfXZTwOye1U53OAoR8W1cUb1Im6Gs
4zL3Tk6rAm+OGMEr/gE6pDPN9rPCyWc+ZFZ3K1UN0OPnP4mVPuzisDErN0xmm4NKVJoXN2md2LnQ
FZKAvHDG7isiq2cY+uPD7lSOoXxRY9V8QZEhxG3wC0C9/Cv3iu/p6o0p/bjKSijjYj37Uf+GaAwn
m1qNBkZ3B7SOgRXc/S/Kj0mNF3kBk2AO9PyiaoSfF8qJimaRdTU5ybYrskLrmN+l/+/hr9bma4cp
FBi7vaqTrwWaYynAtCiCm2ZrGYM/GEwDX1Ld+Zno+idkJN5HkH/eKV90F/rsJXYhHRBpUuhXIr9n
hxdtH2sp5neEaZ6RVBt41QWqQL2K59of83v5k84GGfCGild9IoqQBK/UYnQ9TtkJsgLx3NFzUEsx
9alCN7dl4sSjDrfsxwTyhOMB78p0Lyo4gkaBQj4664zYUe/BQM6E4sD+Zx7BYvQsM4vaRYHsGqms
6YQKSRTPoUpnFvFkctbqGx06RMLismv+P9FAA5IIwi62gULAr8KK0Tr0XRj3pOl57XYp91NDfJLZ
xkREdXPVn9u6fps5cxeSmL68lK6JSEkdGU8uYcV8oHG1wHF/b2va11g/MPqRkcR0tOkwhPZ+Ocf4
tjD9tthMbiY0RYDV+Mbq/Yx24yCt6i0MA8AeXU3chwI/kWIQnLe3STR9ySuRe2n3zKXUvDeepWo5
7lm+SoQOsFQbgodT9O0fZazUvKlCL1PhTDv7YCTBRQsG82mRSD4Ll0B0WYAaY7KS6a84+5YiILEL
NNHV5KKenIcuymNBFBcvp37K2c6YZoiBsI+S7Pkm9p7EygAWHuHP5cjMvapFKVZ2fXNDOeHYqMNa
0gLRV7SWfHChvhKAuPJii0ao1jWX7Bbft8FIC5laMtBpTsUfr7k9aisUA2WOjEBAl3zSllV93GOU
k+0UIfg1mqIlRs/VR/O5me0XlyFOJ8Svfm7jotvgZZ1QpXautqoGaPY+LdFqk/PeY7DofYIJFQ5q
9/MG1a6EIX6URzbxOcS5ixcdpth9LHjRgxIaAGVOS+vcZkWcldaTswKG3IXLcTL3qndGheurRNBd
7h7Kw8JZT/mzrJb+PwiFvzA05172/BSsOT+R9oKUDEVetWO2PVrYvm1Gpg65LQVV/bHh8cN2rWaM
Fa+Xa08x6BKY+CaRFyZ5kdIpaYPG3LVTEfvxkY6VVN38wveGTS6QyBcqVuAspsB2pFshGyc1WZMR
9UUubRVTvJw0njpkM2y+00vCMbHNBFPHCr6uZaigu8L9kAawmJy93v/L008s7f7tgHDSoHYryCK+
uO0TJCYWw827w3GzjA1gDYq6je1CRPa1NpLIrMY5D5EavCD6IoqEzdzjAmRNYlG6q55b2gc+pWZS
HdOhcRLQh6Cr1wLX1zbDflgSJbM00WNziwEzYsGN+AOQosVsbvVQj9vMZUYvC4WZZCVwe6PeoQNV
0EDQbqUWZ2jtXl7O+oJ53azh5hkA3wGJ4c96+Hf7/OC0YjYcXx11cgADYBNaSgWVICwi9v0Dq6TO
+EJh8AY29+NY3hqtX7o5ICGPn0TN521zTE7/vAc4P/tfBFI53duL/WdRUGv4dS8yoAbTtGaAbl4E
G0y2VUoHmRIVjZhLMbtyXw2FJs5jBSoE4TnuK0wP3USvmGyZHuI7VkSKwagu0s1m5aKzkhL+lZh3
x3pXam6dL15x+9Uqw4wYhTJ4pejl0sWIAQ5jIno2dzgszDBXSTyDG6/k4N7UoBjZuMKJTVOzVBAc
7gbheFhsMX5U6+/R3weodq+Yvs78WLbyvQcLaxZE76F4oQVWGm3pENYw7UxFyTwybloP5Pk9M9Mu
xgPQ9fpAwgb1LnByQ9TVopy8ouJ4v3KdG5BM60ll/eafveOKf7v0Rnp4QakbfaDirBFL57U8d/mb
ZVvDb3uec0FjkzsA/Y+Ipnvo5Ma0wCvZGZyuV6FNJfeQmQszg/q5prdFLr47KEoUCtxUlz/G3P98
hnShKwTWJPVYyS85hl/nk6xQu0D0AcA3Z7NL7VQrlg2qM0Q+NFHGv0mJCvbsTor7GXae5/xEzD/J
lb8aUmsEriOjaK4gdZRpWbHXItMV0KxSyRmyjalQ0TpclFeHx56TBHi+LlQjMS6D4HmcF33VJ+ZZ
9sRWp10A5y0AJQz86LWJe1aas1gmQHutPw2DusrPOTgCwVDjOVjUud2mYdkUvQrEqU0LPhQu+owg
YTRB2hJCFmZdo/aIaTViu19rwwkxhmPSdawDSgrUEDNZcBPt/Q4z2h1u5viuogAT/cpriJiXYHrb
Ll9eN7NxDR6ZdlbWKha/DAF3k8iodLUMH/Dmzb/GUDQotblQ3/gkwKQElpL6TfWjosyTqZrSglFn
bk+5mnYanIBDt1GhvGDZupcSuSvk6Wm0ZtFGHaqKc34MTerC7a84FMhOh9AoPeWOc8VXaDbE1slh
Dk2yTciP8YaqDG2K/7AKAz7Id6sWifIKt5GYN46o4Ao2ceWBNQdvqNTOQQPs+cRU+ghLfnPQEX+T
PhSI7SpDHpBgTzXs6ODebj78uvq7VFIYkAWi6VTQs5Z1HhGyABPmVW7EgHOQhZbJOkESckneknR+
ahj5NvYiHMcqr1KflOgolg7XVFniNiEaWgP7fTJKlGR5pFiWBje5OlegFjE1VPtdlRuncyoCI3mV
zNdANAdU/Rxw9st2NdzzH/RjM8qEfn4g21ZwXIZ98z/qorBuzscHDJ5BzEkLqoJ3SEQSoEthku0f
ymZFRPArTnmbRGnNYRVCZYDB+gZXvb2lAARlEcf2HF1YEZ0KYJTbVlniWqK11+/Zn8F4op1dBx15
rHDwO23mWObTzC6QU6/1s/+MpsoLnLLOCmOmTecgPT0I4eMs9aKXS/X2XwUjIrm3lDookRdXZ4vG
y/IH/ask9BEs3W7koAaxUWx3FeX0foNpHe2dcv7mGleH/bSTMuuo0GeC7qzWaDwSe9n4k6Y6INkb
t1tB4gls2Fanw+A+W2VydOukUfow0HlR/zOQqqDyLb+gdnv/YkJoxH6g7qyu8hcTjimUcOd1YBJk
lyq6E4EHGfIN715bI2gF2n2bWumz8q9kzkIxNw3U5MIYoEU2vKevWhj2KNxWH/pNLaYq5egzbq1E
HlT6juAWj0PxZIBO/GEWQjKOEZZMivy0tR89oUcTpZnpm5nZBjT/xLirABSoVUqGlQtLXDgKAIe8
NxusAWE/ljJQNTMqOBNeBQzX+fLOlM4y1a1jim5hfGeptgQRwHIk7EkCPwgckVzUKEMgkcNzn3tS
MgbvusvHRV2yRxpHSU9s3tImYjd1jURIn4nsDoW+97p/pJc3yHF8TQPrJImTGjBaJKLYark32elQ
4GIh3xCRlZJO0Wo/U0uo+UDUHzE/8S3IRRf+vGKZmAC5d/WodB8vZ/oacn321MEgpuprFVbEeUht
MHdIwd3Mk88Hb06xJN2mPCSrsACqP0+cPlibZ5N0W1XxH80g2fnfeCDDHs731OtKaPff+qtNhhmD
Z1lvlBsO9xomHt07wXrIKKtmlyIquWn02rGIGmTsOfMqqjR31jvWV1NYTnIPfRHCLJo+9TU4ZRb+
PSCRlWF6Dj0LBelTCrR1/J/7LU3bld57VFP2M1EA5Rxw/sQDQaximhEko6Ll1RGwWrFaT2fgFrvI
vyzUmSbtu79ht+78RQimUPjnWXOck1KKZ9qeTj/Tf+WrqCoSg95OSwviPmq//BGMKNLI7zF6rAvA
H5mMq80vgFZotZSiS7LtpLmTo9vCDZZtxV+xYraxs2yB9a/XWa1/d4EUNXprXIda5PnFP74MHcqD
TSFU95EjBazVcgkxA6hn+jCClr5ilJWHqrPfkX0V0zamaWJe2BT61SOSGkPEKc5N+o2m94KBP5B8
Hirn6g+YdlvMMMC0V5Do5G2A254UlE4hD5CktNg7tpB8kQ76PwZlfJQDkhB45e2l0sgXxKXSzCxu
agiqXgyoBrdMqnJcqiCb7jRmMXQZI+FAVNJbqqetAGmcQNM3EgWv+UVRPpOcPCq7Uwca4ztcW+t4
zzjNZH341IwyEMCyJ3NH4OVevgNukq0KRB+M5wa5h0rcQfjAIjqTlqC1kgQv/KPsLEIbMeP9nBGV
UPSl/WfKF4UmH/Jc4Gjz7fkPRjk0APalQYOGZ1hz4wgBq2Hm77Jme2QMSW5uEZ5ef0JIx0TN0UXa
4t5xZObAtKj/y5jEvWvQWKFQE1pmgXqgf+JnAzeE4syOzVZuIGP71Pfv4ZY0yvqenNpyXmL+sYy9
HAs2hwImkOZSHBCv59euIKvi5atN9Of5pnGvTb20r1gnf5WIdd8ao02XpH2fHJZfIGqRQLDP4DsT
CaSc+iaRf7/862uGl8pWSJm5oZKvoLpeM22BO285fcxoD/KoYLyDIAFpbssgeSsuq/6uTayvMVOW
SzZYn5u7y8VxqQFQxPTcfvg66opf4nAOXO5rEthZGPx++rtLv/t5/jrv7BjF5QpYfTdTiLLudX5V
evaNTB/7Dqa3O+chZY3trjOn7RctCFip/CIvdebF3xkKmJz07cUTNGhFHtT6uKiahwPXQs2TOyIe
IeMq+6P6m4oPcTC9bM50ddcA3aZYgafXht7nTrFU4LK1L8HC9yBHsFlgr0+1do3b+XlJCHS7X5TF
bxHGKTMDSM8PDLzYUNDq8F/RWoZhLdedbQmCTLU2L7xUSunzUuTCNMZ5Wi+DS7fTuY8U1QKwVtIz
tk9zCNwk5iUxlmSxmIBy7hiKBFk+4VGhsqldxYlvqrEWun++4C4hsbLslUBwqJ1lA0I3qzAis24c
MR8dsmfeBVnP8TyA+XEDoi28AxdWTV8YmjZB1+7lVgy0a+taZDgLs1uyhutW0+5Mm4CsEwc1jjtO
UDLR5j4yoyd5+QPbAnOyGiFwR3R2yP+2PypcxZAINLoZsGcX4QHaWWxZCed6oPB3XA1XO0sJmoRj
H9zq83MIVrMcynd79u7zmilPcR1a6fVUkx9x1V7gpkwu83l0ryYVpPXGJJqmqXjR88ec2QIKQ+tB
E3x5B6lgL1rmhW3F7OgXsF6Z1sHrdUz+Pfi9zE4TL71pmBKHmhAa4G9s7PhC5gbC70W6N3kUWVxP
L4Z+GW15GDKoRWg8wEfcj70JxH2kt8coWtWtOTusC25lGZJP+vW2Q8db8544+hRVeRv2/Osb9o0E
0yGYyHP3pLrNt0hrYnn3xapYekFkXMa+Bvt8ycuBimPPi5cuW+J+nE26m2JIphJfCLzJ9W7KNFpM
928J3LSfxMB7dad/MQFfeKTsiOqxnd+uZc6SitibtMhQvohLA0lGt8DkhzFlFHa2HXlYu70mUgwH
n5VmY9rE6Nk/NQ30e/iqusPfmkVrMOChjAgumM+pQAL0kutWJYqA/zt9QXiBxOY/9snLcfS5uaz2
+7qHNWhMsi8BNjKg9O0HpNWtceXMxUUVwbHGVX+YCRbQ7Fj40UBrQtacvBZ6dfoBD9y2ZdleZzjE
dZGLKVSxKV8Q9KWx4LueCORXrlEwqQdkSL3kNcLrB8RtU/fWQ4Iud+RQvwzDevHL+Zz5q9e9Umg/
IS2qP97z59K5iElw9IHMFKRmyQlvMc/uxJuVde/xuCFbMMteyiaJOODxrfm67vMpi1sp9K2btVxe
PalYCPCBadTRrcMZI0Yz/Ex4f0YXHmzbhaMmNHFJJqa82cQlp6Q9rhm24/RtSV82wxNMvwG9T4+I
IwT/kwkPISESCNWaI+qRVwQ5VUYXsyaVQneZhr2X/UWG/8LAL2hkVSb5RcKdt3fXjpPULYaokN4b
+uyG7bylTN1/2udaiGu2ROrXz0xJv07b5cTjN3LL/PQ6BdkNTGGBqieuSfNYiqphGXh+xK1ff80E
ngaEQo7zASTJx2B3H/28jcCO/CUuiA+ldIUmCiaDuU6OoQCWXVX0FnJ/g/twi2VqIfoKd0zO4vh3
tpUUR06mx3nqQjkJVTFQ7C3jnO5PHj3tTct294UR2s7HDt4G1fStBdNbwT5bOFdLkoLWZiSrEEww
Ig65zEsQF4v9c213nLM2yCBwvFOoDsBzhutb/vP3UTtW2qnAgjHnHwAZwsB9N2IfItcB4+090J7o
9owOMppn7vKJd93qNISULczFWxFMOBhTnD1LnhVT5d/SWGovV+563YLzHZQfefGFc6afUapnYGpb
5OvfPsVGqdAjymdBFJslK9TpubTmGr4sSzyag2ujom3JWftC9AySpwo0Wk6QNEm+b//he8cqpItD
xlVuTrkgJl+Brchmu5ob6XquGhVcILGnRCndB+8/5eD2OeRyrxJxlfyhs8RnSg/tcv+7H7rnaQBx
xrUF1gj1teVThGjGy5dO2yh+wpWiepJLmVMxEaE5MjVYyDrjmjH4EmcBxKfrlvScd+TILQ9RI9XO
w0IQrWxAdsG9Xg+ypIBG5J2lwyyyq2Ac/cCF0lphxQD+v2VyTfhNw6lIY3gJw4B8cCBQeQwi4mkA
W3Z7yXRnHGTamGnjdzYeTnBJIkzgZ2uICNBEBFZYb2fxqpP51cmnn3T7XSC+k72OpP6wiy5lfT3R
TLTes5SDHKaUkHa3Cki70fSqVrtygGSH4tIQB5245DRlHaS+aQ0O8/qLfKhwNyEFVnVoIK67pUj6
EAY/BA3B8lmwhV9gNd1J3c8804yLU8IqBSoh0xnm6aFxBNjm9JSGZNrFzBKvRyvJk7TCnz5SRbeH
rIGOMZWoLf9R2RMKM0zh5l28HPYuzNTjJPhadeGm/Rs+NGOjBHq/nWWxnFQ6lMOQKVn3IQQBUubs
5YkyTqOvuVo8QYfiWQm4q7ShQmx7536APdUkQrXuuHAU8rwCuCMmdcC9tUO0OuvPIBssgO2kOzOP
rhoAbWhz+VqY5o7EWbPYh1MosJ+0g5RuWN4d35ECg/8h8O/oSgldKScBUWU8qus5VC7ZMt9RqieD
dcYHxQ3uDHWc9LG52YCSwEMAgD0/j1cEjEmkFhjAc45gf7TDSII46FLz02RCCMMzu1igk8Ekibk8
v4tyqxlVDo6hb/2puZt6h4JnIidSKNlKQtlDPkccxdmH1CF0S9unqYVHPIEVYcJTho8A52kiTXAH
FTGuc0TIsQzNGR+gf9apZUIGuoqNsE4r99iwjyVaCVkgMXr7xR0qrAtgrndsEXFCx/eR/Umq5w3W
bZR+xhGsHnBb7AVvyYkhhanhGcby09rQqTalP5Xr1+/zbqG8I82Kf0Xaxy3/lRiiy5vHdbKQkWfK
OSBzSk5sZLkPOb4epTtCLvb9BfNWYe5C7S/zxKvCfhgpxR8mLN96RR7zG4rNEuowlmsH2AbJOMGN
Y9Zrq2kBMEfIh2S6rnkdEDlfzpKikThaT4JWeWoHe0F5+Fz57qeOf6WZeCsKh2OEFmvUCgM+yftx
JfnmXT61rcpI2YmGrG/5kHRy9vHYNEUOagKAkV8whgGJA9eUVLMk0RMjUq25Q2e/fNCtY4TjkY1H
mp3Df3et05jK63UcTkfjerhCW3Zjgk6KPD2dbfT236fpit4/GnJYY2L+0WORvU9+J3q4gVD7nmRV
y21CPkTOtnD9kLb6P7ttlUX9FaUN23hN6cme86HUDJkhK/rQNEp47eOl/RQU0Tu0s/7/CNdZJf7T
qRIatOCGRPmLp5SOVZg/IQ/7BUurhBmvXZmk0+L2Dlg4hi+xxIdbhk4IIhFXAI3wixe5fMImVEdw
6cMQqJkLE5Fh11ixuTEKp9CNOHbe/rU3fCSc+3ilGdx60mgQSCz6y2xpEIwSJ04tKV4VnjYGzinQ
z+aCxhkb8OUuzGtaBLd259srd2rn46t/HdSn3KDITOQalhBd++uUgyoGzi81mijiRVOjTzcdp1YJ
uV9Rvy6GwVq1mjlm7KWdOPL4Jid57kJGDJQjJOIB8/sKs6j+rAi0qLpHgqnVHhEw0GQzQVAvia0J
CUdKQpqKaCe92/5zEqpxtsYXlUQZAnlCAZsNDLczUdWQrwNYh79yt5J/mwimE1AIrvQuEPAmTrXv
DcsUKGYNy24A3ZffX+tqxNYMBsXTcMQ7+K52EmvR4tOdSvXPwKbRbyOQEhHE4xmv9Q5Jzsplg28F
HvA2xNZ443mMSemHjBKoEEvQSTCMq4dQcZ4fB1VrxmBc4+WyGZOB5/nTgL8UNui3+ZIPbW/enQOd
xhisHvDNtSfdDNqpo1nZ9QSRRRbC50seAid5dbO32Y/AX+96oMzgnZ0cubugaKzTtGrTPYrzfP84
Oe3//x30HLPOJTvnSHeffYVtRldPyBKvuQuFIZzPTDGT6mQ4l6M+QrH2ZYgxf14mr2LncaHZ6xPG
TN22BvV8lCb3DahoXdJNlCx1kLLJe7ENXjXGe2UnHJy+ONGaL/9G0mB+NaV4r6VBBq3Uf+txkGKo
BjhUC4LBl2uoaRk6Wpu4vicodsMRZdSM/yEh70w1qJpntb+/XYwF2qiMQW6ru+ALkIT89gk8hU+9
nsJwJKgexzuF5qxcPUVoIkc735dznMhPHfasSg/jQ19ii28ZFm2uvLytxExP081XFlLXqzSP77NY
RgpVT4HAJM5JhG4FHGER16Bk8Qn9RyQG4EBwWwj7d9TCswzgGEjyOX6vkOiaYcBAhOuM9g2lwQdO
p95zZW2X6WHzouBIHHwFOvJHNI0gkVSuI/JwXRpHxjT2NJc2uCLyLcrpbbyYBEoupH+iyr295I71
AAbj9ZSv4PcTQYs+njGNZEH8PhbT+X/reO8NrSF7Y1mEgEe6Q40sdcusRjG4Yc4fggCiodD+1wTs
gH/P0sx/imJWs/LImUH42s6gyf4OqgjKQy8T9Mol+PLuU40/MTkjrlrweBqlB0dCC4CLcXP+RZe6
Uwvm8nOH9DFO+/VFlwbMRIP800a7K/oh7gxqBmW0/QeJOlXljzTo9C1NXZ7Ig4wvxzog0nODSnrt
lzSoWcHZPDZTJ4l/t45D0Uz3MD/opAvY9YJF+VLJAIWk/Bb4HZEDFDDj7mrrenxyMwVXMpTxY2uJ
KcElhe7QmfeMU97QJ8JT58wYkAv8Ypvi7Dw4I/hyjljyJvrKks7gQgUec8TsDRR50K13v9RKDfUT
MJN6G6+zqgaZaDd+PepRcyw+2JPVJwnkK00LqemZqqWxiMvjZV5+5B5SSfRW+QgOSescmc+VhOmI
dG/iUs1vTS16GL0lKHHifwKY6+/D915M2Tyy2VFGTKYpsfCtfI2zu2x4rCeetTO5G+osUgUcEwW+
wYi80gmqvm7W1uu+JyXLt/1g47gccxIMJOetACsnLoIMqhshZoMojNfyh2ZxJfmHEsCga0qCdm8G
wIrHOYP1WqaTGrOITRn2kuSbolKJWMPsZjhSbVrS1lpQuJD3fLUXajb6/w3bA9RQJLMVAIrtYZze
SHGPikDRu6tZwBVYQ7MkGimTp3y/37IqGfIrFJTwDigpLOs0xA9++OLFHcFYBkGdGDBTb+snpIwa
paHfZPvSdKlTx96Zj33yTOmeFXNAQ7XqqUoo0VEkwgroQH9SjZMtluvGyKFqFfRP37HBwYu64M2d
v7BqhCCF43TTjp4xooc6yPLTrSDCUCXbxN0yV3Va2Pll9c90laKUNNKJ3U0cwCVxWG0VUpSR/XjH
c+y8Am1Dh2/KBtCoa3QuUtcqINpb2OB55xpXblDgYhSPkZZedNR/j3gqAU0+r+Vaan22svmT3I8W
1rpJVezNankHlb8yu+6NCQk0FYusMzWBcJcTdTkG5Frx1NG0YEgQ+NIwdWVPLSQ4v2hgv4xMEyNU
AwsMjxelByFQoYQ6DPlfweaKOql05NximXEIV/XajMGcw2J4JSymWdZ9x7IemXYUJUDWRoI1tn44
95HB367B5GDNCxVGL88g6dwo4HezZIjTdaYi+9AzQvZskd+e5CHJMbl/ZE2V1dRep8c6S2jRoub1
01HbwZmiSuzKNPnLXHv/jl70iFJIrITi6daGOxm15IFpn+qJFqWtgNOtSA1j+YqxraFBVuWEg41Y
96H2azGCJwBNljSyxGLC2DEj4zaQnmjzB2Is0wDFsghWQLLFVbTWOhGgKhNM4L+I0WgHNAUPUinn
KNMg7n4kiEMhz0vxQ1k4+fp/JW1plFZdZY7S2+vyha7TJypd0/JA7JDhgn6v9jb/Fr7fOhN6OMZw
JUOP4ZlDZ3DUWZkr53Kv8R54/R6iIUdpaYu8BfOD2W/eQroQnvm6XyAu+cllGmVdxNAyfc9MH7oF
yqGZqFIbOuxZcWG7L5bX7tf2e/lbXzb0uEFmt1CERSU6wTFZ7Ag4ds82Ez9pYcrtrjEpdqEraXK4
94VdxBCQyHBwYnVq2k31GecLWgErpmUyPJXZYaNz2OpKilngXufHNcVqg4WKf/VMaUwv8BkD5/jO
v9KSTtqL7068DgGmxaEC9jfZ/ahw4HDuoWRUc0PbWz186jyA33NsVVmOqwwnsE73vFH7RODZYLJn
bRb/C+4HdC+fzR4/zyJpStO3G1Y1vUNI7i9cXN9oDLMe9XWOUewBhraTmRe5AGRP0eWzRXQJF9bu
dg1vof24LsISVt44KzoGXR4QwxXD87J4SX5SL2EM5SnZP1OKdMI23Reu9RHP2My1vlAT88I/EJ1l
08gmf+L2JCgpYmI3CDXGrBSDf1BjB0l7DJCuUz3XjsAnpDGauyc7w6c+cPqaaxvRNkYP9hhoRKEw
iB+okg+r8OKi3tN2LnNrelTyoeBStupRR3BfJipn1gb/q/w7jI8A6J0E7viL+EEQurtu352j6s/g
XRgKboF7OMBzSCPBwfhZ/LTcOf7pg6Yh/0zQNU3ZaCiRi6mBWQUyt9r4vyqd7hom4+8McOR6/3CP
neES1X8j/vOvdWfw+d+yZ0YmmXILp6y4HR69RcpSNap4t2Ahe6xXkBSC+S4sLbvBOTWCE2mH26e9
xCEjeKvq8Moc8JksNPk9Q0h88Wxw5+rMmI4dcPp6pyQ7h53YFM5uo/hFYz15SWqhgFMPPv0nT4OK
dN4Vqk/dArWeXkRjWh3Q9/cG1LEL3EPM7Dw52Fn+fHyjn6P2BRX/KX7NRuZswQzJCVBwa95vDHnr
1z4+j1CIU2cga9pZ6qNqlEO7P7YnJ0Tk/7tcNbpf+8Je/v17NLbto1Fp440TjvkcPG/Mp1lh0PDW
AymukYcKe1ixsYaOVz/K8KMaGnZPRX3+Nj7N/wQDKzYk3/E4EnLj9A1ifeM+9vGtFUhKAp1kTvGq
eLn2q6pdmykJ1cmhEWhUMn9/JGwKDmfjfQ2FE3zJMprhQm+ZyJ2w2aQB+S9DksWX5CoUrQ9JXz4M
C24Zqhk5axAMD53dM7yqJAMHrEXgEq+81ZFAZk6LexXmpYeofAOK7aKGXvNs0dxHN5Mn5PPLcxQ6
uyCdDum9pjgFO7EBhKJ8WQtieF28K2oJ96Xm6j4WalkQ2i+H2C+xBrIzDRHbLcYfcYbGXbEJymNq
PGyaGOY6pdOlmXNpm7/20XJU+iTVNLe6sQjHaiLETX+PxSOhW6V1yCSf0zbTSAjuKz3BHwsjwchi
mUVnvQ8KD9gNDRaGnFRFPLcupAoCX7xv0KTk2vbl1JmIluCq6iDy3t+fGdupg9oy+8UYCrzeMBNI
ceczycQ6DTPXBhDKEziW3WRv2P/p2ci6lB3h8GHji9ux720w9/ivJr9bN/Z/utKtLQGEtD7vQfED
zg4OUFrukBlZWQq6qVy9rDE6vlvD1CNHvOr+FoNnPz0CfgVWBcGGLFUGCoZlDAqPPKS/uXcJs5JT
ojBAoFhMsthUwmIpauA7ymgf1XetjHpjdTQGmTcce4TtGfe31dmqPBJ57hhMw3mtg93u6S0nv2hq
HUN1eW/MKEgX+Ja5J5C4mKDV+X/cOeQMKUZc7tHOW15ZnURfzzMxxe/guBbmPsy+jwkRFsQja/Jj
NevJbQZda9K9eOPmfLYrr3MiRYmSYrPReAvdKDemMBSKuZ22TzlRs8CCulNLbYalKLgAdOcLmd+f
AxID+WGqpCQdvJaGwmsVrLxigt2rymVmGwqCjJornuo6qFTsumJrH16TpX93DPhXt/BE0InmFNWo
QFguyyZpyHjCmQUFMRrrA8/OjBlnqE0V/zC/BTA1TLv3y62nevRnCUOtS7kp+n8nX4OfA3Rbwmtw
8NSfkGiNzCCtXlHAT6GwF2nly/Wj+jcG6DWhLoHBME0cXncdbN4fqqVRNJ5yAjzhaqCmo7qcyT7F
1GGy87FQY5+34zqzbspeFmz3qUsDRrLzsdirrPtOn3fwKQkpMlCq9bP4WgyeJziPeFsbxoI7alyI
8DxDEtrpYmu21zWvBxY5Qm2JBkilFUUChXwYZ/b6Cmxn6xRrjI/nFONdVRQGC3xs4MDVxWQGXmF3
u8F6ZiAjKAI9ghqCXyhar5tgUUbXZHSlyKZf3v0vPq32NQ9npY5/NkK0mgF5hovqkfgdUWU5WwAf
pxdpM2CmChx47NENCEHa2+grb73uPA4TQHtFHI4UMYFff0m2CfoHITZI+jEM5jdKxEi29MiNFC0m
BBzrRDCIE/b2+Yo3jMtAWl5u/VRMZlIhg3j0L6LkaB45Ggfcl+j6Hxvu/2/1A+ZMbODfGBvvIRcd
MiutxjTrVQcdWIcEj3HjtC88KoJNn9Zk2/K99hS5/Mo+kgOHkaIL0asgxyWJ+YZ8vz5t1+5IpkUQ
uC3SCCpbeYgURPqhqaeiR6cJWQpGxhcnoDnbtGjVzHNcY9g7iteDeFs17gXccLdV8FyjYTZSaDPU
UBk+GpOZm7x89sRiINDF5+oYGNSh74aTGetA9TZOIkS9lWPYVUVHBUzhzTP3sOV42NjNxuvWoIbd
xWOL44iKao/U3P+SCpQnWYr2zCpKXQ6C6HnQQQoXgCK2aT3nHWn2cUT/UDIooQRSU3MDL/fNTOI8
0KzDwu9x54UY8m6iZPCo9QNWL8lbxGGHAg2LrjCZjJZOdOeNlgTSngb+9cMxxWd/JdWbuhJxULT5
VR35CUU1zi7kk5X9keRo7rfKvmgxEG4S+QrgOP0q6vxGZb0dZYVgzTQpoJJH5Y8TWHZ71Th33ofU
F1WBJ4Gympfg3zDa45arBa4p7pKw5GQ56yGprwkUI4sDdmGSVu+f3yJbW5ZITRwSt5dqLtNdJwu0
F05KfGC9F3MRoPcK9/M7dNdgBSnOJ145CTeKQIthIt13oCWpgU6nHqTN4NkhAk5uMZAmvbaduQqe
3ctGUTGR2jiVy60eNq8DySWjQcmVrDGtfeLayLa+678UvENXOehkh0EE91cmyu0grG+Z/5bjcGxu
JRh3HWc83JiqzyV0j6O95XZxnOYCUzJFcCOS/wIG8wED4Hbe+3W5e3pots+C4raRd+VO9A/GChpb
WfVM/h7FqjGvnaT2DVESc6QApRP7hyo6ObpyF9Tu6jJQsHgOgXTxU5Pbjd/pC/DpvI13RLCV906l
i2tNmKwRZ4qkywbrSJKbCDx7+QdSscdU4y5Hrqt7WN7ZYT38YWK/RtBSHE5OYqT4Jbsov/+UiHfM
jLW/IAeRfyIKFEKa4ebyK5Bh2mOKlMmqi+cmLF8yxTfoQl+BTBuy+G7vrNcWBts/kWmCBRnz11f5
tEHpN5HaSDv5qvjijZU7l+3wWOo1gWimjjJVvNqbO611jFNKDBxy9cop3z4KdxelKHJJfStXUj2B
ZscNJzahAQQG/dSTdHq+oeSIGZXI5Get8TELXCzFF6LG7/XPiAvrgzG+cTf+P1OIv+FEVWZIWui1
hnrN1Uzgcrox0Y/s1bJDesX5A+gFoRIIuz3Fo0/T0d3cOOmWFSwo3j47xwFR9bBkjGr5YxfMrXvE
SjAHsHS++P+r7ngIpYSwebw8ddMKTK4QnwXfVaKVm5PLBWo9rq8pV7LAJ6lFCIFJqYuCdbEGNvuu
AwFOwVp4rS2dhTFEqR5ygPdmqpWUyCefBQdcXkrzgWQiYAGi87EjAYCgQtsHMbvv0QJTrL6S4ZHK
8Hs1MUidQcW9dYjeEPwB8cKDyG5CJlczfyCkDonNkp5MvY6eEmR1O4LCOP4OrIgHyZOT0t2wz7fk
Ce6IDTJVwuT9Ue49zwnfYGrBWXhKCqStZqpvHQ1mIzDLpE8RDhifK6asn9bEirM6/WOf99zkuFCE
2Vr0b90UcpY8xKiOKmdXuu/YoowHJZKYyGpZJhFiWW7Eeymx/7sk1oG6UYoedUIl1losrTpGoMpC
vNG0e8Zd2AKMhJj8aODSqsiF7/QG/WE12170FWbHkj0IBn2vmSDozABS8EX0QsWHVW80mhuJsLzY
n7ORfpH0SwznWz8HEb3TTKnmEyQpa8APrmsw0qqH41V6F5HHb1ykjSBXfGgAVXHJYgzjS42cj1G1
+V0yaChA35o5WXdAHcfrx4+Cwgl/40SPJagskY1H93GGAyVkHg1Uyx8nebw+gKDZtcNLGdLpt1O4
kzKBIiZvaMCeCKBj6Fu8UW1QyQqlAqsBP6pMmaGdQy+0mDVLtOJEH33GuRo3XLkCreMET6nCTM0N
zu2sBZBZM/2dOlkN21buJ9VQn5+tJeCb7WvEs6LButYMXLAf+YKrz7usco/TFhLmLAa00LQijYdo
rKg5pFvttTciLBfmR51DQwjm16Huz8/XSCKytz4C4v+3ttwjVCG7znsTtFVVb8e0LfOkSs5d7jS1
l2Gjsqc0WeBcxBVSRekQRiUzREICuhOI/cAefBDRQcX1Ya0wrCJNWgjXzrCj2+GSRgAU4gh0u81p
Lvw4+rG5WwK/tqykEttQRHFLA6QZsjXPZxjqyWCWR2mcYluZF3DoLKIoVGO9VV0VlL09R5GhrGJV
6qySIVzHTjHvLNMgDwlWGW8+v8Dbz8Cp+2nq/ZYf00T0o87lVwKoZJx0ju1D79z0ET0eBvivx3ux
ylUQZ8biI3iEGrj7nSRmb9uu005BHaVbrrHNu0I2ZiD6pstlSEcl+BV5VUyt1STqcUQVjh5EyOXd
LRDXIcKdzKUGjOxNhvvDyop6d+0oysa73cEtPdQblGSPSGUGTzPZNjrHGbaQby18Z2qfyymAeIY8
U9FHhazRy0GBSvqzK4E2kvTMsproJNnHLpCoCUFXSgLtIYx9proEKdPMMCFRsmwYN/QSqPIFK9nv
bkxBaf2Lohv7C0qEUI8BCjPka1H1B5jKVBElT9ms8UktLTasSw49FaqRaF7biJzOL814la72pUG7
4HZ3y6cJl9lhZ6LaoCu1Pa+0UTVVfqFN82mPYLdZF0p7Zws9fXT0B+b4hM8MoIuQj+bAoTW3iPnZ
5MnDN7rZicd7ssXNweOum6R1/WBxfa4K8S8q0PUq5D9qp641tKgxrrkwFTEGGOoyvcYqpj+Xg1vh
VpujMGrhMiE5qsMku6I/Caifdp46ZVV3lKsb/VvRcAX7HgctGp4VumF8KLKUpaoAY4Zj8g/ldjha
7H/K0/6xFvudoWoMduBzUOaQ9lAxwovYnAw3qfUL21vO6aiIXSVjG1OVzFEgecfwv0z1Zm3cUhR3
9HPuMumSmbGG4ag7NBIus4iku6IcZjJXhrYAaDdL+eGv5P4LnpkZyzGBICEiMioX6HuytiUt4gey
8U0qLuQDJVRxfKEb0cy/AbI8Ex0pR8Ys447/NS86TRTd8o8ugmwsTu0Sjl9ls70Q5xtZAlWcezxz
BR0CKMo//XNUrKCeHu6El2/Ygou3J03dW0ahmb5wec5w3jo8QfWOy3QJIz2NpPGrBANf5j2DTRzI
qhlrOVtONULtqZRdyavS5QiPm3KAzBE+FAVL3otqq4zZsZJfWn2BJcYfBkB4/5MO2Yk0mMM01FZS
y9J6WCbMxUpV0RgkUeUXwFQGEwWxClFEkWrFoVpmrnVNnFlKjEecA5q6xvAbduXnh5f1jhIXinCK
n2swfbPVdaOVCSa5eQqXZ7feU0I8xRq6SAYdpX1IeHsSiG+qUiG4FLipZQqPg5nfT+iWTMuHIFbw
ncctzjqaAKa858acS18aZUaH8f2TypbW0fXXZgr4/KnUsV5E/Qgipklt1cYzTtEyIkNXFoFWZHWl
vnxzsENxUDbfcHAciLFZUc0qEM/GEKai7lCk7Fx7dJcUg4jc4R5YcvwypCx7xTL685R7X+r75Nzc
QHnkWX7TYxCuc4cIdGPHeWd363YQHoSXhcL1bcyFhQWCp1kAXpROPOcQzrDNQTqyuaDQ8a//aYxz
XmF0KFWgr1i2xW9y3Q+sIW6SIykOVit1vek5Hp3fmJojmt7qYdvtL0HQZqu/f5HGGhVRHd0kQWSs
WTHozJdhsHK724G0lbyotJ7COghh53GklVcHBZY4Vx9gZmccEtAs0eZ3pBfYca/g/4YyRXFHARBt
n+x/N96/XO7DySrbzID5X0EBfypDi2sW8AMFYCSoGI1c8BdIquZVQRFBBPpeS6/y+qWNxHqefn5N
Xt2upLnuHQBN8avD1UffShYZGKvUiyj2fxRkVTqQJmMTs4k+cjJj5gaKVy1jHQIRFNvPc90Hx6JD
jBcVZ2NiRvrALliUxf6zOgTH9M/GdkIPwSfnwC8Vp8Fh+gUy4OjNchRR26e9zzPrPVYo9mJHc+n2
2qhql0SXtvzARcRYGlEkO6ysivG1w6rj4b5CqpWvSEXyTMQHtUiQ/YmRRCT+iuPQVHdiqTgXLq7J
c/bxgvvZKdd0LYe+5LeOHgyNoD1mihAlG0qsVh/GABGDHHtHp02TxEZtspzQ3OIHpUIIZPhkB8Os
vWYgYtZGJ5zndpOYLTvvWxJwXlIRuDgmsqDYvpkus+jjC4MBotR1lHmrDcteb47XwkCKkCVbsnjn
QHmRUr6DEG1pNFoCkc6Qqp5r2G+IS5TeaKMsgV0JehD3GAUpIZaKWSsNlJEo43u5MZ1T70VCL1Ks
eA9nzst20tTjtdnXOvvpd+1LdghdnVpakhRDITSCPnutyW9KB0lFhUvECczmrnjy4fGR77jgWdD6
zYMguu94Qrw9Hr9qRrACO6txpla9stEQF0eZM/H0feaVurbSwkmR8d0lxNJgVTVswZTP0/pwDIej
riA74v5KLrQ2J/TR3Du7tzCTmd51CTgXqKXrVbmLKo3bruiK6zd6GNp6Ss5Wx5h+5yvw4oEjYS+3
B+R30BwfQHyLPufZaSPD6rVK3yYEYuI3ImSzdFepdm0JBL7BCyISMbiu4VWiv0w0N+yXoaHtHJfX
yFAvFb15kilksVjdIjH0Om4xuzldwdit7zvPWJM8cmeVDGauOSuzsCrq0d2wcZhm7BhsgkuyachM
UslvonWO7D5S8nc6Iy9C5DDm02WtKJUNnyzpLB+ZygB4jFIQJRpNNSqAuN2bal/c5sj6guRUTBj1
b7o3ckItIWRSj/1F3bseYcMATX8bkyRj3VwL0KoeJLl2BF+dhbluEEtkhdlT0DWFrrJGwK5nZK9I
zHwF70ciqP4+qGXWemumdG0GWIu43YBqTJHRnndGPiJg+RaFoyem6YpPe6mwWAnuxkpa1KoBDv9D
Oo/u+HgmolcrFjjwCZxqpDnrWQtSrbnDp4Bq+sG80MrtvCwQZER2II+rqXpVKpQWLAsb9aexm8Tv
B7Hy6gBP/673nUhJjlfG7YS1aB0O0DnbgM6T0csy2Si2XNDU/r+0aP8DP6eHORqEg5FZGqv63ULW
eYt+nB99zPThOIF7nkmjoLEOKkvyrsEp2+xvSajeMqdKC+yUtMHk8lm88na8kRkviLGqN/FXN/L3
D9JhQ/P71c2smedE+CmFWD5y4RxiS3dXZrDvUVCCkM5eQ/xB/105ml4zjMg/7V2AQE63cn89U+nz
FYx193vuo+FqkyfJpkXrJozZgH7iV+/mHf2FVdC3KFVJl5RtPN2DNPfAls+v1c4S0OdrGb7uLQeY
fVqMxHht+rjU+qdi7yg8mxwvna82fcYd1bJDrv5cbsTMyfPnn4qX7igIuvixu/8HLqCe14cLI4P5
udNQJ8TP/IjtrSgOzbLKWLguG9A3V9K/B6/vU7PuzFq6AOfIvNSp+76rPo7U9/TwORCaUN4UfuFc
GxVl+8fNdXmtCISQXI1soZ6SIY4+dRdu1018fQIdnC3GlCo2p0Xt5WvaLF44tKyVGw7UN2aE3vhp
uDalBXBtcxgGX8mKRy0NXuHFWxa1lqOYrYvich90XLnqg7eh13kyMeloKTeFFWXK4UElFKSPSOCr
Ca+uuAD9bMAxO/8BPPe59hPz2FswjJK3R8fqvIG4CcxQGk3898Le96umtqPsGSaqYshGOqXLlOVl
CZrczHgfUs/yhtXSHpipoFJSyX3u4eczY5vrr0Z/H4gpY4rk/SPAot/BXSJXOs1XpziJAOgIcJvy
tPwoGZG4LEupEOKJd6kEqgSDosYI8t5txQrnONbTjgInm1UZxspTNO7SgXczbn+7oMq7BCFwgmtz
Dh2oVF6MR3kD4W5uXroN1SWGBCc9K9MOz9Z1jiAq1jQXd+v3SnSIGW6fmv3ZBZ81okjJH8O4GrLq
5y0+37Kgnk2vJ/OSFCeNJtU0rQqsshVaLUjED8Uu4uibaAsVYsCHhCU1OBt6BOZGa0VrYSoVGNtU
zoM8zRVm9YMrKlT61jAtV9se6OtPBpHT2g/xScqJMALk4xVlZIIAZxzSYalYHM14ipjaNdEzQlzg
Izy2A2dynAUpaAVvpUudUFPTc+Nwrawe0xbhIJ1L/x+WvTE0yvGj+ZbGgjfVD0K5c/FA/5ms7Snc
HYJ9/9T7YJL1fFWlqJH0JbqbrO8jo/16ZhKbrOT46FzN3KSXGONfY/4vinq+5mzvLER6OmIt40D9
Hv7Xiqjqnnc+L9XeOIY4JUseQpBlZq3wonVOjbLlyT0R7nCIfL32TgHPFFR9OvfWxDQIIKvpAK56
FhXFaZWSBRzqt9bQ2Ug7GMGD/JTG2wv4weI13vezRotN6wbdtBCBywWTqDk5rYQSpiZrbgotk4Ve
BioMXEjA2pONYlEQnnWLnqse+TY7sPxbSyrUXLtbMeCdm27T+ja22ujBTmRKhxSa3lHOeINAmNPW
FAtPIcv2g0sQoCYcAnirFQsg+CKRYP8WwJM9HostqfZAogss07rOYxe6bDqg9C6PmmoLUlhO6oAl
NZExKzBOx4s+K+YotGJPgnQdJWXvXiI8kDrBjVihkqPTrL+LnPZcWtqT+aOt1RVktxYaoOriPvlk
ey8rMN/A9fJg69kduiMulIqJqScICNPpp7rINz+i9ooVqDNocHla8J145Hjvm+XpJEm3T3jS4GGq
IUBgS3fNlCwM60/EdgxJNeoZ5Vix5PP/wN8w51k7JJX3nZGIlfE+aYP6ffsZGqlJ1ctFmBVm8s6b
1kVuxXdsVMQK4rLCVMh46P5HZMB9vPS5glPs6jGGJyQds9gIoSmxmBzlzwdTLob4Yhw2Ot8Be8rT
dqMZHRGWXhhWOk0wgJX56q+Oa8dehw7ECvphavt/di6NWvGh+EXYJsX39V+cwp04DNT0OFlGnEdS
Ffap4XmdzmZnqGrm1tnphMF3KASK5c1Y3DyMIsmWfck+Atua8O3WwqGsyBUxC7UOBJFYZO4MElmp
HppSz9uYVCnpn/rSBiss5Z4i4UUrEeOV8xQ9N0gegO+l6qavVsa6fFJ0ZYatI/ZOsxvTXaS4UPMv
3W1mRU68qGxJSwov/wjd4uOZjrp2KFVKg4n+BxzR69eCkq1rTCmlQjJBOMQENG6adyeWDGFLVUHr
/Fwg6+AjfS4g73VSHue4IMENtX56rt9AxBp3hu+RohE2CC5q+LF2rdn0Hn/GUinl7C+vc9DAkkPP
wQbjpzJsKmTKM5JaJjp7SLobmqXZ+VLZ1/oubTnOyh+tUKNpFvtXMzzG7kDfF45hz1C08d/rJGN2
bIGiv32S8pFQrR5kaXSdE6S72azFTj6DzmJkohgHuwhMN9znhP7gXQMdnbbWX/JJzZ0tmUhBdU8N
UtGHralphIdeW/ZQaRsqf/aw9iAM5YHpZczTXMq+EVXOohEMeAMEQOnyYGHJPy9jpX4mgJ6lChMS
VCGZxGy+BY2XqcEThWQ/mmtflW+B4Yx0ky+gBzFFZ7hTlZRgeeCbkLkwuNxrHWiD+q5C8q3YfS/A
PyccvSeMqaca6RTIoI3juEAVHfsEb24N30XwvPzcvCLKZ+l4ptNV4KeKtAxoJ4wQgUWUioHUaxIk
5/9xDDaJhpL4o/q504OyCkLgBDK64PZ/Ik7fqdiJcUGyLGdjdu+9ehBVOgKLaa59OHmRSC50fh5l
dtPRKP2tarDYE1Mjv+Gt0VJTnq8XDCUOtEPJSs+a+vA2DABPM74XybO/26owWG6SA5LkG6Z9ICDo
YQCgjMLEr6RxZUsBFWDvBz6Spf3AJIJsd85VpO12HopehZ2xGTbTiQTAbtZISesnOFUiE5mvEtXv
zyuKObvKIRZyRfp6tq4wsyH528K6WwbFlb4kyg17I5NSgozGZbK+fIdbsiH/U0ghflBexKhOUt5Q
Gw6Ir4hY18wPqCbpVuswI+9itbBvOeKG+8I4E1FM+NUO75EH1HZJY8XxcL+2V0+99VwzwXOYWufe
3Pn4k7bVICppc8p9oCPGYK0EJq3u9FJL3bUUwDMHEE/n9JWV/1DPzqPKOTzKNiAd3n6rTobGVm/Z
coZ49CoxMgZJiCs3AibhNelDYv4oJngr4lAikHNqKGoj7Steyur6Sx1fN872Sfuq2oB6dabZl77o
VjROMWoldno1qpvVUn7R0mRL4oTidgsBhGWLO1BdOsk/OZjrJXqN+FN1a+FIbF2ANKIOJOoi+rKp
5Y6srkrbyD90cH2rS5Gzq23ETWZIVqGgb6TTaB5Dnrd65dDdfUQf3MeuGO/s/JG3M/D1OJKJJ/cI
Dr3KMezctAjAZ0N9plNf/j6JdKaJkI5TqgerCkXB44QqEW5+5mtrhrM7aS9ZWPePn8SMmmpD1cpj
cwB/jspYPThstRcpcO0LJLB5H3jMzFV5sXM9Yoru5tH11xuvG2uikObB//x6L2giXuZLM5ziIxRh
oIIQZFzucVVYHpIYfK+leFj6VmoRYSvjSjhgJs0YKDC/Pm10vhfr8la41x+3u6OmGBNb/8o0wluD
jvmvmuMElpQ1h1MWFE+Hi7vyXfD16Kb49pxELkSh3xCrJCIEjzVRQNyjwBW1TkawgiyIoCho/qt3
N8Rby122d5IVhg187G9uFbMJK3nseVqRR66QE1lxWnYWoJ2uKF85U/AjvfyT3IxlZVecNXgnxr/5
BeTIZbhjsQeCnYzuIrv+IwOgvIRGzwYCVQfos0waG/HqZLcOZXs3dV9cE3tCp4CbMaDOfkMiIPdg
2rMJ2NoItdbGcvIA3XwJpxl22UFNJYfa/EszRuNGATPDVMaoRD7feO7wy5J1kGGvv9Cgqkacp+KP
grMTOfOUlwuHlVOdvHdHnxTRlTUeC9ONqRDZwjFqot0OI5zhpf/XXPM6X/ylBQJiVjMb+OZ7YPvz
W9cZhKWc26rdC+5kKqWj1veyZ82rxYCKKy5WIe6qprvch8Kwor35aGYut4LbpyEBlSd2/ri3K51F
Jy2KADYeVovS6A5rjr/zF3AakdjvjVVPs1OnPLdTYXKAlpNgz9DGH55xjei2SmG4nbQZS5QOGLZF
ahiorlULY20y+4W7ftR8Hrs8abfo9Zbdvl3KYXQPj0EKuQcmQTH7m2MF51H6/+zZhA5FWm4nlVMP
Os9C/3mlE6YkAS78FkHf0uLzyHOKJkEYBsONdz3bKT/EfqjVbIeLlNCiNNoKbulvibOUyNpH1Mhy
vwxqzVk7UcE9APvha4mHl3WwSsnb6J/TSC1qOlOadsbrd73aP4iOB5VSBZTnuA+xMcdtWhzPZE36
7UA9Hy0j35dxN3s80nDyOZV3G3PYKsZV3TEiS15R3P96n0ynzfvmWDDMshxnPEm2yM7VQOnrX4+a
oUY7zd0GLeNo2HT/gzQT/vjSaW++ZpNHsv70RosMA/gdht9VmAYGq/wkrsQPrJ+ikAHS13k2NoF1
uMqInxMQrE+IL1lNAqjr1IgnoZ3BN8/vD9j3EsvY4diAhwn8lNjDw/YcR/enwOoDYDQWEv5EVQtH
TajX1Nfr3foAnaQ3xAAtaHAHopyCUnD4U+vSPEywMb0WOV4grGXRYd0LdevR8kDzKPJaGN0O/KFG
/X2YU09ydYekUOPOmFTSdogT6Kaq7TLLhnLGind2HaqMAflhgtfi8IaRdIOxbPeGgRuVJfvcX1Lx
oct91eY++a4kRr7ELWJ5/t+kNXzvWNs44qHJOTPlgrwfgQayZMmHSiuFoWDrOOKOQHEYQIXXkOBN
klmx0YgY5Vty5V0dsEe2eWFpH7PRah5GYAFZLj2MNG+9wRbOWlTsTOKVfJtroKH8h5IQECHDI5bz
EKJOIz9m2VyvUc7ITyluNB+uJySfHV6103akLTYdheMRfrRwEMc80sJ2F9WCU7jCGARPc96CFqDw
E32cL+XlC4aU6iGCbV2kONiWlgyVU/8YZyZtT0nrp70WSSE7JYGLdWugT/+W8pS2cvW5ft8jU1D2
2D40WfpIZjF6B0HSzgQEloDYb1aCBNrthsZAUv+WS3Qkb71IQ+Tac/iYd9uNkotZYgakPAX1Ya43
igPpNKqKsCV30AQ9wbgzXMYT2ifNl3z/SCF6aDCoc9HthhJYHkzopwxWOiiiqC0iqDkvFxjKeD+F
SEpzUanTlyqC5wbaN1otZt3WlxZT5yoUX6ahq0ERDQRAsUF7Rp+Ae3WRMtuDeCbC0bLWDStzFPQk
Vx7cCIUZW2Sa98qTunNOxFjf/RyLyNGe+Dp7VcxrKK0Ia9IMOi1BrKOmShMQogBPhYx3P0ep/DZf
b8DaRWMbB7MUmMrJIcPXwHcB9FIS11slkeGgws9kTdOUnKYIqwzSM2F+ccgiKH2vvbDbw9STFK7f
TLJUPB2FIakYA5IPS5VfCLIay1yo3qGQnaJeDSRXnm7VgUP/Sei2wKJ2z144r0MiRwMxP5ZnJsNK
AJdGvFegPufBkSVs7NhODriC32eGbemmHXBiJVCZ0sXyaer+AtJ2wYvlHxKh5Cs48F0xJjzEUJ9S
Qn5WgAMQ/jxrI6xNqy0FzZDtrKoxghnu0jdhLyg65nHg+EW9yTaYUAayRr5q5YUuT+2nMgybOnAb
1KO1U/RLfow5vwxBAHdxDn4s1YwVO6DdkpOeKmDN/31w8sLdbF9W2gstt//xWhe4lXfHQ8MOeuBv
kuw2UdxjKF/h5Bsmmo9KhrQEf/QelmcMTSHqPfzJvTWGGPdFB8AljObvaKPlNJvOZpTnqah90ueb
i5uaFAl/qQUHu2zDY6lTnexweGdQymBkgE9N+x0McpuEN2QPFJLLXVJtjGPLoabxFK8waYOAM0TG
vlxvZ6ri/lM+Uy95Z2eURYs3CATEnyEnc0XXxLryOQYSo1fI70m+V9xzPLvLfdEZ6wF7nCFMT8Jx
fcGfhCUxILb/vvkAaLqPOGN6qstTFbIrL7NlxPzUwQJOvs8J+hrorZ5UQaQEFu33bOAOKMrTqplA
9p13mu5p9t2MKop9hwT+Fc5dWCrPgnhY7/XESW0H0H0PaVXMCuskXXl+D5TZ0fvLTWS6GP93Qade
Cs3+JVyhNOCHMAs6YmsnJSLDS0C5NmpjwUjXecNM60GHTmHps/RPXNePiD8qc5wo+zZUWWjGRWor
w0G89yzK/gUbmM7vYri9XZ4Vf19B7i8kT93J0pdEQosbrdOeKrKpuLxRw7Gbz6GX0ftU+MApqswK
XrwKYX49UceJaXcuh+oOnkTRDvIxLrO0zZ4xOE7W64gH2wP9RvDrT7dlEVgfkMxXjY/Qa93IHHEb
e1+/N6Tj3O+FYwCw1Ct8M+h48G7lcxUk2PLH4WLNR84TX3UrIish6uMc+jaxZ5vBfiHWymGiCYBz
koQodQmhl1EwRmtI+6VhyNY50bK1uoQUZwq6frfQ9naltZK4GmsxcQi3cPFnT4URwjcw8l5SFwlS
6tB+iUuxs7fKid1+/vwWs5JJZbROHwp4kt2cSjeyrbW0EMxsKu2Pq1/ViF3S9SNV3egRaug8BIEO
FE4AJdZG+s05f+cTDy/IWBWBWkXVYkK/qYYWWfPSCY4XJBQww9ThYruIp+JFme+OOiOAK5Jb3zGV
lOiLMgcWNHURJlaXoQCE4+wwKdtUYa31xuergnxjMgXRgqJa9uK1T7yZjaYqMc2zmy93Rzw8NBxm
FPgKDX7o46M8vRpGPKHUBDO6MTAlL/TO9Ij6lYZ9riSlVr7yBw1PHZEabiZEyQ/Lyiuupe68lnd4
Ku+VBDhWKxw813Ppb669vZ1A8fZdAeI7DdLLFiXQzQyyrmUBausQUJxEXjg2A+R5tbkK5MOEat7J
WWaYsHfvQE3qSbrewXTHs17utToqtIWKqFcNtyxQ/iA9cyMhmX0JJwuWuZ5CEeqoMd6GXJwBcIRj
qKXqugoW6Pvpkis0pQaHIExbLlhXU6xeg9wlzhnUXRIlnK/o59YA0FxkGF5f87Iq2RKUh2U+vJDD
TI6Sqp/DiceXAiO5/slesCPT1+bhuUvyaQ8OKn+A/KQYkd5qkRKpJJT8jLp+QpkQs2TyglhjT1YP
W0Zktktp2q+p1DksM+3Xax2GJENiLdfM2M4MnbKpmbpZqoW6MXlZs1Efjfs6WS0aFzeps+yHPB7x
msC3Ox9nI2CqkKmvynS2NLwcRt59UvGaHtHJtGCAoWU7lJqN4ocfEUrK6f/+mVZPrUD+hUwOi3mI
IJkshDwizszV8hFFcdREwpzfwcqOljstuavTqcCXA4xI9IXPNIloJVbhmlYZgmaqFytnl3SgQ828
J1kEmal4zbwm4J9+h/uUZ2nNG5UDKKhsBkXvZkbOjtUw9aQyu7Cd8B5f82A9cFf1JsJWFxOraJx8
2cxwcg/iNFUIKtD4kyeUloRejPhSivLy0ige4CqItmm7Ynu5thXHH8CHQhIpTeP5kgjOXmnBX+ll
ttz4TKpjgngzWuLei5Ed1Fpl/zXD29gqyudSVbxpnvb89OdKrD9pH57op9VK26I1/6c/38Fgrel9
XgPQmY57VnfFlMlmsqPVnqQuy1f+9gPNaH47oT86AAV7OlqG27Dfrf7xHgfNQO/6ufqDHYGyvdDW
i0IEFnn2YzTpF7b4ihedm9T7A44S2c5OCMhz2nILo+ufVJOzup+cfY2BCNDa4XS4jpXVyJI+7f2A
6O9lG8+UVrmNnQSUYXRAqW2FjAtKozqwqWS939+pn2yuYbip8hlr3L0KDrOC9F1UzaaOjL9GmF8Z
vNdg82VqXWzLLuPnmR3RgVN79gKbzUtPpdghsIlaluWK2D79QjRnXygMZOqQlGtda1nzpL9uHtDb
8DHoEpJSavhxTKeifIbjTzsBn+OHPyhCGNa2bSfw0b7IHPYNeb6ktuPFiII+vFokLrBY43FcQDOW
Se88Ue4+zaA2mRF3iSFJJ7rL7DzhiW4rcfITaNhRzLzaiK9nvy3m82EwjMbu0HSr+agIVdA+DpQT
zuD3Ss66TqyWC4XssdORZZ/esJ48gCucdHkO7TP3BFcFsLif2VxY5u0Abc+HqKugFAIyTK7+9iRt
jQ9UQ2IH1OozLIj7ojPei0lfiJQVk1RLO60GPuulAft0XvT5v/k3y9AF85LF5/0UZ5EPp1UmJ++z
B6WBEVLCKpA7FKeqg9K6ztEswqebRJkkPj13YMdzR+fSLy0FWB0mx1n36EoFv5X/VLDZgKNPTd3z
o+/QZJAACszvThu5VAYftzqDIRwTGONupCp/Akp0VIl0S4CfZuTxX9h0y4k3B4NaRYVWUHGHGh3X
KWeuJiC62I7rHWSr7oe0WzgIAUNvRJEyHMDSRDoDeStKq7Ny5n29rpXNW+MF2p1V+pOtrVaAhuSt
T2pKphL8OmsIv0vdGVDJ8Ti3q2cTZkyHF8irzBe8rK5COuvuf3umzbp7tRkVi0LtUp8YHBAMeuT0
VGDKipRsM/v9slJHBTOw/PvquhHU+Xh7WqmArWo//jlDqv0ua/67rM0+lzTQH48fc7ANAvB9ujEw
lx8c6Mcm3jdOTMPxt82ctyL3WMPhGcaSeE2IcztfuE6mPyXFa3cR5+Cks7Pj7hOIN2dOS9Zbon7N
NKN3ENbPel1Fq4bXf0UIbI9ycpwCdMt0lGSY24qz6XlHgDxQJs+DYSXUlhRwDKn65ugv8YaT+R6P
DArH6QRB6hqK5lfOn5mbgGb6XIyF+bPVPGCqZ+Tpo8n2asbgnGvg5Uu0hrIQbj9aIda3TPmGUxx6
JqUr6n8HUxbPD/bgoOJYLNQsSqg1i3EUGoELmzBVCz0y5HBu+uC4KxRwnEY2k2Y0keIJC7yVPv/U
o7ev6nZBaZPbiyLUlC9ytYW13wjQJgSZJboR7rtrVx8vgv8SR/h2tT22C6YGwtqw+AK+y+gkygjZ
JpgvPhmJAZ0dzkuT11EBbytx2VE7yQZs6LavBgC6qwr8cF614mvSGBl2ST65F/1MRrQXCzLudQt0
3DiRqw1PCErJpT8+rcRssaxtQSLPrRtsWuZ1J/WHWb9xWukpsHyy6bkQ+chBTDIxCh0lxb6MtQaT
OUNE7PTgg+NoCeZ6FxQjn2HntCgOwz8IESZf33l8csZ3kzjuLzf/+IOweHWk/7eQwB7HYcwju6Rg
EJqV3rm9CYnsLsPr2ssnkDpBd3HV2KAsmAXVZUL29Z/dZ1cwtFLM6Ey0+4Vj0Mk740Gz6KdrYYQI
BlozLsGhxUCEYaXavpeUKgTnSwrzJNQiYCDn4CQ0agD39m4agKX3DRx+EfqzwjylHqb5QV4j12yE
cSvcPWpgPuGxkALBYJ4pGgl1X4e2Tuqgl9HT4vCrYWsp3rhlSEkyhveQyh3UnF8QWyD3YvRUG/BZ
17nZ7RELXd7BvbO+yPmkNp99Kh3t+okTYmtLXPLM/OrBDXS3ah088+yvr3k0Z3ztAHWtUI6OnEQk
A5jGGH2tOPZ7dxLXP17ygqAHH8PAAAaoP9oDa8UEbsfrB/maa4RkyUJHK3noYk9SY7aCxzNZwuCP
dyQkbN/KLZK+oiXqDDL0MweXL5a4d45pUllRBXMCATifeRwsSl7epuEtmJ+7oPdU4wHzGvDOR6u/
H5mAoqlDLzRhogHwcQZs66d9J/UdvqFb5aKR9jtI/QFp5VfIIDaUQW15M0j+bX8n9wsKNjO1NFdG
BPa3QIGKo9aGOYywJWc1sI9ByrNnzarM1l9mqJ3RUFJOF9O7keVcPxuu3UrJoPfSmIVDmwW+G0O5
GIKDlJXI7YNSCoYt1rHEwXOcBKiB3PFtrjAshpMTGHLZQpG29ZPpWqv8nO8L+GSJbNGINGCW7TMd
3bAYo2XdnVdjqs6mg9Mjpcjg2prSKVRKXqo1V/gbpveCjb9ct29AFIZnO4ioPvwm9G3DHMtjrKqJ
L5EQnlVfPdoxdaJmOSiI1lSN6XTaERDQdLK5HobytUMCQssh3c8NsdPB0FF6sFRu8Ulwi3PSl+Wx
wTfGCRiUKPj40+OITN98/ph8Q46e83dGY2YOWol1Spw4zTwJwLIVpI6C/C0pBXwO5BoVwpNgGm0t
GVl7PmSa0d2wxEAUFYvltvg9BY9af4oi3q5YBRH6mlSoT/Q6aKHcdJtOihhK5YHuSlY+sHThOhL4
ADLvF6D9Co9i5GFpN00FEOOjhHCgY5ReTNrt3zkO9I8Pc45VKGdkbQo02xPxA1W7lKjdxwHs+zR8
rhBK9B91xrJG3RRL3pTNURxGPPyLQTbcbRFYIcKVldODF0uadsVmOrvxP/g2SThzSAgWWR8d6yKJ
ZVYG8x94AR8A1qFN9MWsp42V3DZp2/uWW34AHStVg/+L0mXE23u7j1hWdg8w9SCVqcJqdsGerdou
LSs/rCx8IUb5dG3L4CH9iWD0gV/sqfn6KNFMvbBzQamS63HBv2pFkh91V+4hzlYLalgKPI5CTPJt
ZQqEgymEQspgYyf515QoSc0BU2Hmz8LkUO2SwjSXK0ux56PVuPxT4/hAlIyTedsQ4X306NJIgqCj
rN1VpRt+6XpRUIS7lA14vPV3a9CSDcWwnnzO0hPAG0TicuXK9mfgg8rZgVqETG0/einprVJeuIet
/NbaLwlbetcdmbTTNFWX8rdaPLzgw9CqGoMQ8mBREGwb+L96X4G82G1TRvahuEydJ6NaJ7CwZZXM
6zpMmId4pL74/L6gkuigaatNuetWx5cCiCP8QcZj2yTSMgkmI6EL7fphGPkjBRUHxeuJzxZDLCcb
Skq1lH6oNeK+kntm0bUUppjYgEEAcPpFK7lzk7/YyvI+ahNrXwN/sAstBae1+OBwHbu2bKfLhtoo
M29ElRDkpyn2xCo4Bn/01YjZmQ/thqJUiLzEN/h5YFkWyHW7ee82VBpj+u8n55NmjxZTXdFmdr02
05TZK6SnTrk/8bpCV0xeJiBGP9GpnmcK1VDX3W8y53yAELbLEXBRmmnk2h59p80TAliorYH7M7kT
HzHu/42vEblQKL0iKDPPVclm8KbOQJoFbUIP2niJW8V6cjHiUoIv2qNZhyFwpTBkqp24MmRQWEXA
S/RQodBsjwUqpWyIgMBfsPxpbweIPtLBxaV5/5WdrNPcIja9Tc3mt6I+NWERjuW00PbXnBx4ALlC
lWkxjQ6oPSPLQUDUdDz/f4sH0J8J/rfqNDSeY0s2zn1eWRkP3/PICQTcinBKUIAsQ8DgpwsRiFBF
SHVnTEw84tUS+EBqHnItSz5DTEQCXEN6/e3SWsDVHmQSSH9+lDYxvl3UMZvsFtRO2byJxjVEcpKX
pqI+8X1HxvUsKB+y611ofBPVrT6RlZbu3EYZLJ6Yhbuiq3Maj8l+e4bSua02xxk1JoG82qb29W+Q
PvT4USbaw0u16XWGqtvluHGefERkZvUnGZh0lCw7MdPSjt2MsbPfpT/ifKeJnnY//D0hXC+GOgpP
xX6NY18smmhJRPpILHm8LKcwjO44Q8OYqFdrEhLP4RvEovY8VFMUpCbn+1duPHrhs2XnSpgmRkJb
zF/Q+T8qEh8kgZ94PYGy0rgW+zLCcpV0MWpTn7OWuCIJq1mxQA2IPYtllXqQsJXtRWmj1dGXtD26
/Kjoa28VrT8sq3dEg4SHGcO6vS7z1CzG1Lq4UUBmb/llW5Ei25L0JkU5yOafOu4Gy/XLudpmyb4f
3G/RG6jP5w0tDjrGIashcEmPl87cYN3ZNMIzwllTqc9NkE5CkvPNNpIDngRSulwcTq4DLBXOHoUg
oqEDSTCtbox3lq6bd5ZtLsTLqM4Gq0E4Kxfm4SJNdyCCXgfer0OZvp8pmREKLvdEcVNR2GqQ66Ke
gq8gElbt5sq9VqxB2INXF/PLP7ukhx0+sjR8pcvgyiuMWxwq4hsSBlIhc7TSdOMWHcWuIK/x9CIH
AzqD0VgQHEkCDvz6Rals2+WFfijkUxnKGbBCs0DHIxrwEzKz1fHXHSRK8liaC8coeKM/1EHx9KSi
T18bLrAHeRKEJ/aeo+Xg7Jf4eANATf8YRQGNcqMsHlKcBalyxS5KU2IgiNWD+jMZYEFYKJcNsUHB
sfIVG5r7UqFKSQuM9JzhO4VCej02XkmNLSdvz72O/A0bA5HArKHOK47S/pPg5EXBjmBa4g1Srzld
xUql62mxBI3YYtLPGfCu/lvOvw4G8hMIKHp+D5XY6jFWG3s086vBcEZ9FcV445s9T8mD7Z+rDd7i
zygQicSHYfTh8VKaca6yyQVnHw1u9ynv+B/ZIq4gfNVbMYZHwD1X6tH/UOdiyBcwQc6WjBqEnG9R
4qdnZFwWM/Xq3DRi5U8Mvc5lOr5JkzolzOGN/9r+hgCRkWMuaYoz1J4C+RWzmU/ulh+zTdubFIze
bOXf9rxjADcViblwkYnHkhMX256984ymKLzg2IzWhyg8GmfUJs8JLBtRJ3f0cpDjPInmaN2qvdql
vKxVlmiJ8MdDsscF9HkiRPloet94Ln2a5AZi0XPjh3OiBB8FQqyCLTDFcVOk27Q7r4zan8LCEx7w
Me7XoazeXzcjUBj10GlaVPk4XYaiIyIki7M1smNswG8DvFXRZCPZYVey/2W2btzJJJ4WMw2kZdaZ
WvMEQ1IIV+3AT0LBgdWzSeVGib8yOtFGA/V4gZBbwwNYgfmdFxSVYKseGS/+uwRR6FoR6nPp33p5
defnNGd8WhnYepjnhGgxykCwbhMDDBEF/NrTR88B5IYiCXAC0RY8RWpAGGTxPHgXKWyR6Swd/qCe
rfx/PNO2CUuXuCq0ASsWNsP1byckpvG4NYsC+k+0e/3hz87iaI/zYPUPx8/J2sB3GcfS53XQNBGD
maU/6NopwA/FdkMRQOo8Neeo9tXlNfKHkXLuWPUt1RFYuk9ysBL/D0rkPyfwC5CQ28UC8pvmfQ3G
Fru5SxqQYk6Y9tRiLfaGBDGs/c3BJPSKwr/8bj6BGNIuuzOmQpl9Z3e2Ue0uyfzWISrlnXaGM7fX
hllvL6XXsQxA9juen/njhD5T6SOWxop3KnrxBgMAPYO++axlRJFbXwHQqulAmiVMU2XgEqOiVgJO
edFDYX0PSxxtVcy+vNGs+LNPMoC1JyoH+MWF7C5Xkx0WZvT6YirK/iVlq8ijo9S2ITpGpj6DtGIk
zWd66WQwXFw9rm+Ta3rSm6W/lfUTShvdxWDXnoS6/8ZmoiXiuNMCUZdY9VOIoBxzxMRqDwQ5UMWF
V1gIQ2WY/NUoov/AnamMgY2S7fMBuwsMZz2LrCHhVutef6Wb1XjqvBekss3idq36DY8uGxvNfIdD
u2cn6byGovjRR/k6hKBjcwEXkCGlABplvanh/V03qnvl+A3sIaybmU0BX5b7ZDv1/aHE6dlI8LRR
s3ip9xoRoYyzVOHpZDKEY3hyFA0ckBq+q++jaLTPje8BRX7LaBjxHs09ccGp7ziOujOhgtIdI42e
Xa/JYgh2XGqdmZ0IB+k8kOZKMQ4kbk48FlxIvpmMTUnjztSpTCS5Cy7+nF/9AcWNsQNt0aIxzVsE
LcHVvw9BIYf5TLT5JggG1+HPczLsQR7ds3xuo+8afW4Fj8aNC7EdvrO6sistkeXS2Wzx0eu8UjwH
qH5tI3og8CbBXvF8JEIxtB4ieODfJ/C6urj2tggGEfuz1I4wGG2JLBYB53cgDH3wY6Zp0DLwfCHB
HMzgDxDI1/4GA0Pj4JbLgiRPSz0WJBOkmnl8HB2z00IpsZuxYjd0j4rsoULCKFvy6IeilxoN0BUX
KURGfkQ1E8YnlGdCjYBVkNKRznazezuS0JzITlToZqqcFpTgUR8S7JG9hs/wC+iLud9HMl6ml9NM
eo3CTC8Xtb/Gs0oruFuFNzni+lqTSr6st1zh42CtDq9KuS/yblCL8tKLLred4Mr2pcpu2uIUpoX1
+2EsbxkulHb+KddAyzODbwwOtz4+rCam9Dmyk5N88twshEcUJuDfb4kVFXOS6i626MjLJK2KymYp
9O1ZWpvP496IoT/cVuuPpzcgaFhdLqoMrDmI/5ONTzR6zQWe+UoBFxEeQz+qun9OrzinkVV/eXWv
J4D9uvWdfVLSrhVo6Y0zsMc73tVjCNvJMXX2OQg+wsU3Urm3OPMBKBKSQzUzpFXbLiHnttly8tnK
0SlLlAvkK9ShUM2ROyxdSQjqnuZR4xEXjqvdq/fz8ShVLN0UgveKyWkdgKr8X9v5M8Rl3x2yHdgG
q51MiA3IKzFkUU1AX2KzPUAtVXih8SvWcujJd9i3qSxXgChYv8yHNyMMSxhC2CtijXcD9KzfYC3j
feqsmh6Gb+bC1DFo3wD7baDG8sWU4biVb/tG2lqfkPB8Ni932fa/h4QBN7RuPOT+QrGFTA84j2SW
u2mk1ijOryEp20b6TUka2TJa4m9XgcfrGo8HM4ikOMx3uqk5KM3QTzCpglwKhhP13VbFxlQNEmRi
FpuM2HwBJIh04ggOOK5tdGUYwXHG9bK12va2zN+WC0KrW3lMnmNqGKwJWp91y+qt5fd8kAZoCyzO
YmVorBwCwJtWmjBv/eyCbImxXMFtgs8AAPgcdP/kAWrC4IZ6uMg5A/DIgV8pT8G4ebuUVrc8Ku+6
Owx1T98sRPgRcnMJgR5tSusl1DkaOztqnvHR5O3XLzJSf8ISLgLXt6wKBTQQ3ov0vijOGDI+OeDj
fEN6oXU3/IdI4+v3gr11W0XNqBGXtHKI4/eWY+ovb9ReQkKHmC1XV8pXTc9MFZx81XNQbPKtRx7m
pr5a5H0k/jEnWVSt6mhZA8+q3SSX7aB53QMeOdU5k0CBLK4foFxnNaksM6fCwkGsn4uZT0GEO2AU
q+/eaGfRDckZ5iYLrpbOcWIUyAOvXuc5Q3DC57i0DkSv5hAyP/Q3UtXKt+2ZiLom5x9Id0WaAdk3
O50s5phQFCbWb0S3FWifpNZ8FXUVWGtXk2iDE2X+C7zTK8SNps9e+Sz0n+k7GIY4Z05dznMMkxqk
jDBa7i5AQtszoPlWpYXHIm8Q/O8wA8f0lbVHzIGuPpOnFxjsFkFmEGnWk5VeipUYB3LumFbpy+tt
OK9fLGMbHzHaPxDw5Ssk/S9NQtj31/fV9z1Iwv9e1rQoExiwdZva9hokcygi9xBCUvoTay5RZgyk
Tl0cdFBjs/Coe3d0j6nINYCp+05Mp1qZ/4CBPZPiJbcQJad4qD6b8IzG01NoEZSTIEzjJK1V9Trr
l4PmyHzW3+E37oEVLMkHig29IWkOHlmHbPpNk9q6LJm8Pag6Ul5Zu8ZJeTmjSkWGRMQydZHQ5s4e
mh39PB73Mo3rKOacgNVbsZSYV3TO3Fx4PouEMbdAAukghiSP+Mm8u6DrTvZpf8Hcsj8DlAXmZQ46
FStCgrQwSqrn9lMeah3EX/JqWhkUCH/lxZVUqp7mOnC01h9qPjgPVhFMM9x2u4E574JFAEUECzjE
b30sk52juutwkLp4+8C9E0RYtSNIv6YNJdVm5pMn+kkM9itKXPX3a+e35Xc7paarDQj5dpZ8hoxZ
PtPDUGQCm7mk/StSyhTH7MZ22OTl3rL1a0ioNT5HAKwYlXkERgfBnbNPc9N0leSNH3SYlDuWtag0
uPc7RNLSkIQqMNX16nxop02tAoo7HS3+3/XeIj/V+bUFzeaaPVL4TnpHGwUt7Ot2UiPWL9cdqrq/
7lDbg+3ksrapQi+xDkmChq8LCAj83mswryDNX4EeD6+80ofmJoL0Ja9vSq0W1ZWSewhaAM1R6Iug
iTuOeY9ZXrF1WlaRirkW9TZ29cic4b2qsuJ54lWHl4BWHweGafKXvvy8mNH9xKB+S7kFmbqjnQ3l
fbrO1NQ7YEL7JrWVgH8hnvc/zja0w63pq4chVCBl/LhXQrp+LHShfFD71dNlfh79qsTDI8r9spk3
SWwJwd+kvoYbOwTVTnPWI2hu1lgiD60QeaNJmeXNRx5bGDOFx6fj0DgsmMjdNBy2hFh5KyVSK0oo
Gfo+koc9ti9OUIpvRpPFu2pnBhUlAAAJqg6Szp6SKkGdMzPTVmSFCd9MyXTyfGwRQacVRjt84b/k
jFtJS9hl0vG01viFOhxYBTDSDxzcT5Ci3R9YA+xQRUgVpHLwzZMQUKDL7asrAGuxEDWYK4XBImRd
HUH3R4pU9TGoAqVvGwU0n1MIalgI47BWCAxBkxQTWGNR1FpCDZYmilnGSGY2FGQ2rTFw2mG71bMg
9dFwkeH2wNPMmdj/fRertsXquwDrECP5t4YJgl4L93y1acuq8LMUEIa9QKiCAYMS9LNVJFhgFRXq
B0uZwIDo+13tul7s5P3nHQ20L21yPIncGBsnzzXpcxmYWH8534QLTYylV4LnhWBuBJ0jsnGQQ7NL
49PbBtcZrA/6/5F1fh0XZq+aqGiZhSgj9rq6/IKI+pzCkPNOCP9fXVzuf6Wa8q516ectKXnAH/sQ
4D2aM3PwngWAaAJaaHDRNrQkfl1UQ77vN/9GBf2Yk0vPB43Ge6wN7hPn4n6TLZxBuOh+TMUP6b2c
0w06B+wxcY/RNPVSWGZRTiROYVuKT9AOy6zyFx8EJ+j1GaRlnkg7KND4A/l/5o/GD3VtoFpxh6rJ
1pM8uVPQYJkBd3PG7uWLI700+wKdiqaUzPGDMhZafkDSd2SfEPM+J7/c6hihWPAAfiCkbfxkf600
7b+362nBjJUwGoQ2Mim9BJwLk5sGB9zxpyUh2Mu/Vg/Qk2YoiaZBrygA6fJp9nnNynE3V5nR6/gx
DYl+pB54eYxwqVFGgcfc9tbX2LwYJFGj4aHbQLEwBTG4dHZ+85HUOBQe4pjCCnhpFnlXgTtY5EXN
CZD5XS6Uk4831PklQE7zB5FGSNMYMsKUuv19asw3h2Pp/bnQf2f+TADzKAHZKt9Ft59UPaxiunm/
ajlRkLHv3e0TyzjJU/bwSY2pdQ6mP99yxoBxfBNa/IBjMxJVWefNwd0MbmFkGORupH6de79mqMC2
E+5UnaB/ugIR7qm7o5kI+VXtph2AagUGQhECDr6OUeIDqrMoUZ7P7vZMLJa3l6kWgiM/A2Gg+g3p
nm2SeUdYc95sHDzPHRF6gFQdl0R4YCUKMrEWKrATCu71vPOQoCVSYHQi9imnQtc+NK7g/nLxCast
cKTP6Jyh0d61koPjq1lVIgpiZ146DXA/gr3rwZtcIXXvjOSNS+fwletEJTtkEOsj0ZIVxdMB5YV8
rgdV5bRz9NDLn7M6/rD0tkFz1aQrEc/O4zMRXNBDomBbDGckIicmO+8S4c24ET1cPaYWHPluCXGF
xaadBa/EO0XNUqyKHHoE8M6jJ9L4lP6YTS9S4btWfBNHsNLZUnO+xj9H4YbYaMHXflwslSAJoeW2
ZVWYYkduHas2nd+cf2tzwTBnVqDw3NDq9FtXTpJg+QC59MWD+lD+4tRg5pl8EJsPHW0Tllu/mgY/
Wd0eMcNs0V8uP+mkXr1wcl7lLlfR4cYZ4gxxnDcDQlExl3zPMBhVkFHKgL3VLXO+xp1ff35wfcAC
e9GTQeCb4aScd6/YLEPwBEnmYbHn1cb960QZEbcOA5uTxbgytDtv9VhOy847rjPviEZ68l0GK20r
knsOFzWhf4fXn6exFfn0FtXPrtfJYZcJ5GeG86ea48KdnSjgHXsrQuStwr12bwoz6rheoOZuVE3V
Xdkj1spCl2219RXMsqIMHA79jXsCk2BNIhm03U50hjL3BpCPodIjhNSS8mvlgH3uB43NaLMWgX5a
BXkVRjp//LkV2BqX4gJzmAOuERYjk98qyzOS4D5CIPaYJ4rL/EoaxOqbaezY1rq3KEARRZYak8fN
KOKlI9LBM0Fpx54ITLWbp2X8XUFQtwHSiAxXWrwMfDjJ8sdyttMsuJ6QRCbv9CAKJiARXpYXcYvx
7ZYQQhe3WZyb4wHA3jTBwONB8ncI1/kC5CvrVynggZrZIhVCntUCmrI3I7k7vnsNGZl8Fe7pS/1h
LkL5plmmJQf5aAs1cd9LuQtBwllWYGraJ161ZmpLEaddRjzBd6Yx8as2ifh/UVkw4F7hoGQ/Z9Gz
7RMgj65bltr4PuVL7eFUYe2GsHUXfV+Sa1HemPI0ZW6BjyWOIwZ3i2sSz1ArmCyLU+e8lpP3T1PS
2UCCvFzc2jrhoTLAF58PVPIruYUxs7DobWohnfG0Pa94+0RQWsANUFgbuazHEwAVhFCQUZW/CDEo
VRaKBqKt33SRpWkogHtTXzPnDsuWtL9N6Agam9L5H3Z2MY9UFD8vd2PXb0vSYCZe02DdWmL61XTX
z6eX8fHB9FMnrHVcx4qzegJBfE/3nN9WPIGE4NK63ju0/uuHyKEbOKRYDZScbd1VNZDRI7lpUxXg
ANvyutJeENffMWLjaREToD1q5FSEjE4uWE/nBF+uTrLxeuy25A7OCOsmry7meuUK4MTf/0vVqXFi
cezrfUQCA4wfUtPouhbBhIek/GhLf996+BtMgLrrjkHgiUBqbj/DQT85I1KPXZdA2hQ16XDa5fGV
5ntTGat9KSRVLh3nZUnOlGZiiBxaFKbK/uQ8Q4dwzfwS+nIHCAZyAw+LTruQwlmGTjJSbGYIH6rx
60ObFY/aJk07fy1JKXPkIXEJrS6fSJ6PgWmDU7yAgviHAOpZ0uu7eCJEfSav2mryUg4cLckvo06s
cH3Aa3eY6FJnhhGm+BLi9/gHNmOprEVWMd4lxgqtkkzov/k3P+h85qyMHNxfaLRB5lvf2Pmh+edp
uO/6eqPZ/kFo5ZZiyHQl8GKeTRugDs1EABecMO0Vgw7Ceonpoe1ZK8C5HvBPSlVKFoCvO6eAvisy
M3r0qaEzObzyQ6W4tOf4jZLtBgPd/WHLkroHAvaswMoYZDV/xczeTOPD3kL87k+v0weGLqsq6+Qo
Tzdy64EVgokbg+L5TtNi+0e+cGyC78+1ChTc1WDxRUnT8CrAuOk4THUkMKh6SSJsgiZKu6krXIHT
0YoZ01frOsOywKF+aLoXyMPX4CECIOWYuRdJbuIT2b3xBaj/ujjsfQT0TkoCd1PJdIh0fiL6eu+b
0WbrKqQeauHaoV69lL77+rnOui2eEdoRum+0pGECakuEMc5SlP6gyEotxiVheqMSfO3EXEcEOMDw
Go7s7Zh5wPXoF5cviQuQNoOr1UiTeHurwfnnjA28AEWfzvKUT1G0ijT6zl3dIpUGjLm52fW+VC00
oULQeYlBK/TR/+XrTXjvSQqLh4T+P64OFUOOmq51n1R8S6wY+ojp9vmJSJ6jmfuqe/aS007AX8YH
nmMO7mQ7E3U7C8IZSoiKFT5KskMVHgBh+inZ7l6Oy3P8IewqCGqAsXrl0UBhcoAiQwE6YVD5Keug
2RaUqIZkl3dX7YmGKuZ/RdR0oCj9TtGQ/om0+cVbjd3n3WpleRjspBBp1kLdlpi0bH63sauymntB
m0QQWlHzozPI9CFV7AVHz7pmqhkWaHqROllou+a68RtiHhluJ86WCSEr7dLcc2T2uR91uQK8wAfw
LBKjyvkxT41t8uveBiSZ2LefQYIeIgzBL4p4SMf7jo4CrdZ1AG4VbB5QiJXgcAkq3Xm/8DnOEnu7
vgQl4ea8oBfLS5jVIofrsWWSPZSSdkjdcwNxhDkipgNv1zdGvCWD76owBvNxk+CA79Gz6LMchP2o
8y30VL8RkZWhswot2op4l851d+wCZqF4qnpFIiQopQw7pQQV/IqvGNvL/f8G75RRoNgW997M1e+Q
mBcw7BebfUKmEVQPEnu5vJ1KeEzppnTlFDvICVDVvxSWkZd9vCJHKFiGn4j/bd+M11rfaXhDNIZD
cEkr+MV9dN5Zn4TqHuQ2jXUPNqfrqj5sPDslU7YeN/3lOWhWbxivp4lc4sXGM93APpETOGP6DrnP
XLPAcfnUkHaddi1BXDn/YE/CtGb8l4LFfu9ShJD5ACjI2vsn6KgZo9tB8CWOkmCxzpPUclGMCUCW
bLrt0SxaAe13JVsuKlgB6VzhROhfQc169jRT2YCUqziYNcoTom6wnj5bSH9IoOb2vkiEnmvG8zHt
we3/bF8NQBe2C83gjSJH3NS7ykQKlTJ99F/HbtGyOg8YBb/wJSvcxvgvWj6X1Rv4iUnYwIx8xFmR
pjH0ZwFJZmldBZg6T1UpBedWvUqcOI509XqnE2BbvT9Vv1wnLrgJ030pJoGFlJ8KUw/qbf2A99Ne
3g4Ueo7eK0YwaUJyi2kwg5Q7Y8pTb38gHb0OBN87VNUgz4s0nR8srHpPeTxTgnF3XGLg1Wulg3wK
bSSGLEsqu6eiZD2hHU8o3C0b6wHJ7ivjzdUYVQSz0pKZ40yGUeE9huz/VuDZGkm1xJVEX/m0no8c
0B9t9cVI34O7iVmUndzlSRaG1531OElSsRKTlt8ifVTalyEPqx8chOQVUsoUZ8Ier7Eu1/yw2inh
JFe8/fWI++ef3MOcaeXY30et6SZKsOm6tdxeHMnsuYgJKqE/A8acZ3tL3pn3xkMZiY0OzIBLEAcZ
t74BB7XPOHz5qRi/Bfs6/+yDIw8Vh2DjQbHJVW74Rud32BMEIKC2nK9xT/BoLV5W4xBv7LlKS6aQ
UrAv1PzeCgr9KVuoMULHrRDjop4vAgOGnxWz9RrpbadWAFtQcrmsn7HCKqXTc4c1/Ocq9BT6Flxb
KykquT0IIyEkTOJeCMoM6/5O6C0mewcJ46s7bG3KKHmkUa20ZPwr8wyTeOUXVOHqdXC93E5i2q0/
CB4SdSDBKybuhkIG7Zzc5BYkc7Ruwli3c2X6o6Z78QrJdvCrTetT9A+fXiznXcmPyyGXVjyl8j2+
wb5oaLsSUkNZ9KtX1UrLY8Uzri+KHCsUwmlsXqYuqhOORW6w/lRxqky5GvSCi8VGXfhfH0OdilBA
ZrESCawvKUm70s9G72zDFgDE4/blLHgPJZPbKzKSYEBH8sX9qXNxJpK/UYCi7Em8Of1RzUcDIVaR
bwgq7CiiVLmK52UFmYv5g+KlhFNtvUT1xhrIE1c/p3eQACFJQ7nwHG+6uzViWZGlVUnc6qSjm1hO
Wk64LdbHhBe6RPirQlEAIrqDzmPIVgSSUNuMJrDHBeRELMEs67M+Dp2V3lvLq2mZVima43ioWKEx
oPddYwa/FW5tER5xCJQq8YxBisWPuuccLgyTNff278nYKQK/AoKWlm4jEjlpbUHODCTFa+8txo8b
CW98BnW4EJhAuAtYTrdW6OOk4skWazrUcV7jvqQi3cHD5Hy4kjxsKg4sr45hZqY9thkcd/Ew0x0e
LUjqZoDSWD4IwYNvftmi1ZIHyPGBIBKjkvXThhhQ5DeWBRGAbnuR42uS01ZK7JTOqrOzeaw9E8qn
m3py834YDxeouTOa4rvtVpJIWfBVLISS830PZ1yLzdQ2a8ivXhdo5+VEG8SeID69mWkNm2cC+UV+
+4no2O+oKIY3Tme5uQQtbRuMivNZZLzMmBRZJSXJqCZxeAm9qsT1MWdm7dT5TGpN1vMrGtKPJAth
+jR3tfwlpTQ7Hlzg0ZKUm2ODWq1Uaerk3QvocIMhVUjjStLKhqkYHvTdeTF8fitw0v6kQ1en+oWE
WInl002HXP2ouwSeO7EQmZFj+GOO6G2CFPCpSHiEXMORSAoD3Sbp1fMrQnPBuLmRUab7N3st45q3
MHyJCLMyAvQ89hmfCaUeAa7snbwRs1eCOKUijYsqvliWlpglNRtqCf4SUumwT4/PvlDKcMGpsuiA
uvA8oAa+q/ae+1SfIydgIsZFJKwTiC9yrqf7ixNwXp6VFLXHDDbP0ekj2ilPGCF209ytUOHSsbGM
2GQRQamfpKMlwmp2H9HBbDIrEzMODFse1I/QVUpr824qbX9Z59s/dVYPekU3QMUpLv/CEicu5bkw
/TsiCjiy/gAl3G1PizZdRgeX3Nl07/tzgKcpFDuC1n9Kzv2EJ4QnmC+qa8zj6cSpoDxE+WBslUtm
cv1sRGBtWzurYogjLGBaUF67bYNGssRXenh/sjv/d55JIUVcGBhwYSsp8cEgWglNpJrZGbTh2UQo
rwr7Clvx4shIlPMw4ogq1VB0ZXERnBBJb0kDkLyRcYFq8hEcPDCdiPaNmsPY+O2PoRK3vOvu/Whk
tf/b4zPpNc702sMHxA/qbRzKZgoqov1cULclgrZu7eIyHNppkOlpLy9p6zkhZcsNY2NHGEFcVQeY
CZag1QXTyrP/Z3hXcnd7BElJjYMGozu2KkhoIbEePHyIscRqi+da4sQAViDxnGf8OOHvw9Cfex/y
yWCWwk8zPiEUzM0bto/j2hursfXmlCissvjUxxK9kBTEnuXo/mcQJNuWnfnkneBeTuwVm15+m3TF
7T2X7+W17uqYb6SJNs8/oLoKZ57xRBzwJ9/oANQZu8fh9/sULnDBjxBnIOolKPBSX/sNJsagZTSF
qrWOIz2QxoevyGNnAir0BTuVWMompGy6w/QDZZaN6ZpJsUJBabzutKzb8MWgEisUt1y8nEtP7zag
ykjcrdDBBNlRH9t/C1PL2XCjeGgpwehiSGCDEN8pnd+I5WKOxexF91jYCy9OIuXWR7ssPDece2UO
QXIYY7RVARYCzQwCsCgcc94gaxu/nVsMssHDMxBcZTNtDBJwmVESpkkGuvIPYi4vAveuf/H32kAi
Cg1E9iqY9pGpcfNQum4DTxuQAB9SemTJYouW+Eh2OXmLdcBJBN+ul34a2hGJ8ic3eH7KadiNEiS6
SrPtfELehI48TM0wMf6Pg75DpIS9IBPacmzRsumYobZ/2xwrgJl4DOU05Z2cc4mEhFcXcGCflkzu
4mwonYwhR0aklsyuuX60k0WSP4IEpRuA8trrbLMsAko3G3G+mLICih9Dp4aUEJ4NM24RHRe8G0cb
1UjZedy62h7klYXbyaVmNZrgDnF67TJJeecd/+R1EUvIEWe+yi4LWhGfK9sYDjRGJrRKbh0/32EM
bgw2ITPyVuFkWKq4/JjNlVxe1qt3tOKRHfJ2N2cfbsdA02s28DiN7J2G9CiXF14pjW2DvJUeNqFQ
OqGcsasJnXlz/XNZIRchtCrRMCYFyxvOB2jxP7L7SA2nUiMR2CEW6SVhDIWJ6KBYTlmki1UrydnA
G9x6wE3FNueopiw0d+7PwDjoz0kcRGJGKnYpAF67YPy3fJ10dNP6A7cR0amz05Ox8GQlaGpbLbM9
SeeCNv6y+iNeQQ/quawfXf2PVSqUDnBs6xSwfJEGVILR074NydmG3LEYnMoIOddqeo7OPwNFL0N1
GqW+peYPIQLNZoOL7b6YusLCC+wfPRGiHCVBzpw7UfQml1jn77w4oRbpSmjfLBd4UBA1NNKH0GpD
9YtmYRDXW49Er4joDJTrARC3Nb8p5Q3O43rm1as9IS+CuAsjSwje1Av16zuUhAKPs/TepDwGlnGg
RUmCOGRQgJbkuWDm4AO+up02+DcP+HNEkzmglQ9WKGlwXWo0beI+EZPU4UjhS3rK55EYn3XUu9xP
P1hUNgWo2yiVxysWIySX/B2dUtMsy1sFrwYe1/4CunMzL6+yCc4C/h87RfB3dulqDEGNzReikGNl
OTDytKGDMhkee3JOp5Mg6qNnJVGVg/1/+FT56c7/AG3i7GCMdghcl6LcQDYLFRhklcOdPXJAtRe7
ZhXjapz9bmMKf6RuBeq8vmzn/spw6zH6YwDheY+4Y1Vwk1Tfo83Qkywa5uGKju0/dIDacZfXNf2e
s8vW3pwgZrn/aduqL+5WcJzwX0RYmwk0ksTM1qEZ7NuFVUgN9C9h3ZzT+M7Rgm/Z2QGNuqavidDT
Jh3UOlHFdwRb7loQQEKxUJVrL16lAFzao6y0LUMftPJYJetS+G26DtYLpDpUHvtFTN9DeARhkVwz
4x9EGQpUvUvwV4vqRkJwAuH/YghpwHH+9KHuF5NTr8MVPtbB00QcHThvlYfvYgxr7rh+6+Tw0yb5
FaKKl9Qcxg3oIN0v3rXHY7zcZ4jeYEEQSLgDy+KXMK4oo033BH5RNXesnewzeHfPBkaS2S7PdokM
+2WUpx+KcN+v7erl9eZObcP+O8yW95ALMZKZMz37f3oGJ2hXa8YJxbTC98ubzvXsrhH1LIxcwS4N
wgk/anEyvFn1JAobGak1yUWjk7Jgsr0rDVmfadmgiEqlbzUeNwF8gtvTgctSFANbRlbrYNsoMjEK
GCO8h966qz51gfAct62LYn//jrTTvnlLvX7cl5A7JuCRzdAlXM8hIH/LuCSAq2ZXEiq6qKZjQyud
lav08td7AC348OS9zqTfMHRBHDZ8ITJRtWVSzBNVqL0FlMfmNpk3PHLUpuPsa/Sos/2ZLWmXR/Xv
k7SB1yWIrttx69W2QHRQqvl+uIthj0WeVfAuF3n5kAzlNLGUR1HN2owoeDxSiaX35DyixSuFVd1c
2mkqZBm63iVRJSRNdvxgEwO+FTatiOHSZA2sQrwtRtM6nJ7+kK/9rRwsiEObc+r5u5eA2Znxq53Z
jgSHhhI/86SQYVeqs839O57e8zMw+aI2hUnew5DNY/oOGNyHTtl5Mwi2TACWRr0zo2ENQFVHa90l
t+0kSA0CVkJM8W32CBQbn1SL0/Ffsqq+PLO31Xh9yzH7Oo2PpQGqpz1irWG+RZkLzTEGXMVh9cZO
/BU5W805HAJPCmhmvaBdcN1/PiH0FCFBGKi4qy0jnrWVBiBSCbyQaneVLth6AZhzOh18dpNKaLsg
LWOYtgd2NWhmSnTbLLfDpYyUde96EoZc4COnRW7LcD9kjIDa/UYgDubw2l0b1+LJM0Iel8Mxd95R
xNpUshemtMJtbfbK5fTYsc28MIaJV2dNOxbBcvIKNPDnjS7+os3muMDzLXU7sNIQ3pBIw+cMVWrf
F84x9y4CD/dIwWcftJFFS/d7nMZDih6gNXHxld2tuqCI693Ifo9eaIcvnZWmDCUBIWPWm6mkEQRv
lwG6Ae1Jj/axHhimwN02pMygHPDVarAJHvyHr+JsrC25AaHgWfqqxK5DG+I+MkMr2w2WT5zlYcNI
EzzpIIPH8YmSJkiWZSg0Z+sKkuG3zG6XIo4OSAgs2zLCkZU6I2nvuXlwyjARA9uCfjhnaB4wZwvJ
AuNOcuMlHyNT73PII7Lig+TJSQKZXKmxvBjxIQtBfkg7AWfXUeNnA9J9qA+PBuzaWX6PImZ9QHfn
0+Ebjb0oJj4UavfmanCEbvdtGrkP/uU3xkkgQGyL0ex28CiyGYyErjdqQwegx8ln7WCzqtkBWnZ5
+I+p6awQx+P7uXuxNdUC2KzjqECHQJn+E4C0J5ijOOXNsQjdW6bxs863xpegs2u22Jux9nZQcbov
6u0hGqzVgwRF+39Bmw2JJA+Rdnd2bpLAlXatMYIrEM+2pZTzp6OjST66XJKAv6jaUFXUackwlyge
0DJYZ8IFCg/C2r8YwYw4RW3iLKejqJCnGA7LDPraSCPlDXpE6RYsy4Xs4sofT5R3YpjbBUfdqowr
uoYu/DeUJCuBUWmBZIkzJFB8a1j3NSoNjWbWqEuHCuNaju+UTqAedBIX+kvjPP5Vaxx/D2NQqP+p
EB7BNb7wvH0I7Svfz+T0ch8Tsp0DTTxNm/mCEXmE3XuF3b/IuyhIPiF6fQRk0vq47q8WXEERIdSI
NxZsaVV9hyy80uu2D8LpliSym7weJqYvKsl93+68TmDNApVD3AXrj7NLUcu4Qg4YIJJxfuXT88br
WhXwYnVnR9nZIXm2h4ekP7M/YJWKS3qZAmRQCPwMC+j12smTMAhLo0bge1jOA2J4NGKbFmGC+VKy
wZXKqY/ofnxdcOhZ55c1orcAnHQLTSpwrtWbPNdbfF49dIBN99lrxL2L0zb0o/fYllj85XMm2quz
RupmbuRIa/6/C9T3RNqYu0XsH9j/TK9Yw5JuRFkOLo4NS7BGafCYm3qjwUKCHNHqx1PPDiffFQ7x
Wiol45o76F+eFVi70DF1ugM90up4cBN1PUs1TL0ZPyKJ/hG15Ii1YVwW3B2R1rr1RSQn31CzO9Jl
1rXt11EfO2lggAI0UStQ3cv3+4qI2YY4VyolV0U613b7c5SXVfDrEG/r9UGRBsqEGKHHjoCi6ukB
3v2YCOJ5Ah9NuJlVFfIrxa0xykDJSXk/qHFz+br1qLXJ3cKgfNG4qExAjXVjgMobDuwv5fEuzt7G
lWTK92hmnvKA/Cd2N5FA09nXrauQ0JaSSIUq9Tf/0fMwgaeUElehgFRm4zn40RP7aUTyyEGDuaUB
cCuRrOnhqF8ICuEuPiyMH5cHAhqM7od4FW9+Nl3DUkJxwdGlsS4J92FuMhekIcOrNiytCeOWX7I2
Yzerg3NouSafSLPIytNJmkDIrUEmRM6EoC90MBhNrcN8pEXS0/quMZPm09ysuhr+BKATPT52QByV
V0UKXkY1oS4XDFwR5qHcsv66qBud87x5BQ+STyh+TPxiqZmUjffAR+D+6ko3zk0II60/UUZMYr13
PfB7DPkB7GEvZoF+ImOzO9HKnCFj9wDlVr/wXuDGBjXJc6RJMxNNhmbmlss91aXGhWBBZYuLDpwJ
wLKeqZimlfm3oyYB0vPwa+itm/nOTUrjnBUaHBSqEdSg1qK1eiO566PCbGXv7A7y2Hxan5HEhx0l
QshrZaoR6gtBSaOlmcu/obEmwRJco3xcZeX4uegyAElVHL+MeYBx36nuY+K1oaLbockJxblt5gP/
XA1u/qUNbqzec5GzO90j6IoIrinyRMlkSiCglWMP8DuAsykqQDdaZeG/Jsz+NXNofeCZG+xLYdFI
9I/+HunPxEe71FutcuiyWdur1+D/G2rrWK2Pn/hSz9OxCGdRYsoaeYUeINKNaT0eaWDoVfWwbqFw
Wqde6Ug2YrOBwE1vkyZ5I64Wk8qLsdSzpgbCzMd7mNpOelNK4XKMvPmFLN4pc9ObT3g39PbIFqpf
CLNNsYDQXiPq7RLKJ+8/KRh3XahS+sfsOzrCCJJF+9UnoM75hTzmgI9f9WtPcjIgtFACYDKWYdXn
EifX30WUU7gNcH7j1uGCjtg9cbvvozLhO/hNoaPcBfIsRhJgF9lm1y3mdnDF9/q2jXV4ZCNudBjp
whCh01eRLEYlxMOKpEdl9tlnM9KvH9y+HG3N6OwD8xbul7IVcsTThz1+LwIJ1/Ooqb9fhbg0zF+k
iUGoyc8QxBIXlu84NJETG+dwOPOgrsXGMZR6taODxCnyZLramfrAeiLf4PrVMG6k3Yuu8nri5GTW
bxNZJ73f5gnF82t5ssRHUi/Y4RC1DoOIFQHWOcM3pfYpQJ9kt3tJ5Ud7/23gNqfM0KrP/z0lCt4c
r02IYYDknARhUG/WUIN3nS+SYiWM1eZhHokLlC7ztgRL/TtN6wtLzs00K0Yf2EStK3xBGGuDPoZN
h3t59zusICzSyfQZm91+Zvjfk0BaaK4GCX/PVIrsNai08UVhmVssiPtT8AWsyHkQ3pLneV+Pm73S
T3eKDEPHb4GH/FoUTYNgw0phriGZl8+h/JxSlyUqFrYRUDe6ErQR+faNDDJqCwwqP0INbAxc5/B8
IF0gZMxPwKKv1WW5eAYxKdP114OJ8fceh3Xpd4kBZtR99Tjsy63kDlZCWYuD5eAWTB+w5GEIqRvA
LhbvII9/OEv1Xxwih0xZmerRZ34YosCRgZSbAMQpPA6thhZNSeFJeyTrY2ZcRYMFqa3l74tcQi26
x2+/Mmq0h6JbuA2MFHGb42172Nq7FreENhS98UPy0KIaxGCv4bMjRpoFwPwNXVbil4Tokw736ctY
UhaZiwLLE4elITDK9RgsSnNXdMrmSadO07ZMBJVCE/oXsN4tkp+2PN7aA+SCKVr2oHfn/kfl0ufF
qWcgbT3Iy/dNnhpKLxhwKrzAY9qtg/Sf+aWE8jz0p5ay0/olD6pvNY8OE9sUasey6ew6XFtLMDTO
A/qCOQlQTcoGznGI4tKCxbSzNBzSny3O0osV+VYQzz58JDWEsjKmNKwCzbYIEHIdDLXdJjQWXjTZ
qdbnUPD7NWoiB0bvwRfaEwP0NcbcBL1t/oBg3OG7gUnvC6BaSRrk+N0w7ggPIDbh8arz0hLVKMjX
PZ92uaQJM5xtGPUhIoBImFP4Dtrk5cm7jZ9R263M4YDRx4mH2lcHD7Dv8GPqB+BAWQbecaar+WM+
xzPjOdHn/JkL+wMpwozDoYMXyzk1FBBUdjzgoM9PBXrsaxKL9LvTkcKsNM0gV/fdHtFm3YCQTQsv
aipZ/m7/tRY/7/ttb2SydLIse6w6tcG+w/qGzAI3PdwGWC+2Gg5obeohaTJFeP8pw9VPCqzuVPUk
ViqUy5LCgsrLOblui6cUr5lH1bLCaYfYu1hZupq/PTi4ySHLTGPKSlOmsjk3skGkeTEXfgNk/8kj
XOTWNaGOIkltBuSin5LAghyd4kw92dqbgiwcSsgStdKHSlcC/9CYcMFn7uyCupsrF9b+VpnqnNhC
eCD4y5Y93iLdYAXbc3CCrSapsJ2SMhXN9bxYa/d5AizVIv1jSrYnqYEy++9TECJMWuAFzDtJIJ5j
hVnFgPDvYFI+A1XoETpg51vSfs7MrRrK5qZWsvc95KD57UMXPTHHE8KsHKXOYWwGbo6wWYyB+ffd
So7PGDwIIzgT0SR4oEUol05HBu5cCRs9T2L0qz6+aM3YhRiJK04pjYyXbcgQwc7XDQWfpjq8zM4o
mc4//XQ4pxob5j7Gba5KWQ5r+fVrL81JPBVhooXvoKVr+fkeAtygL/IfP8/6c+L5SAnNtDgepe9K
gjAS5WnSUPInssVliixj7VMIXNKjvhBdWwEPRz6m72Fpco/g0HbXhTtpuUwInz4onieI85ZmwKGs
GpW0Par+5P/3UwVV97Qw8Ud0tt7j/FPILkm366/nNY8qbcAuuBVij2DzmZDGra5SszSgyP0F0fPi
QchK/qG95MLYR7Hg043WR6YTi2dEm5dzh7V8lAwCCkJ0GtxTD3ouzwtgeo4tSEiY1uogbi2N+0Mh
0ZoYTYMFfq6xYc4vi7EW6ChDsdQ4jzRmbipePN8gb1BofksBbvcZkcPw+jRE0WLSqMsXHRSudVFT
BraJajiQUqOlZ6yEDmGjatzOlmROqnZQfqDivhlg2pL8EkpH+hHm1vJoEKGcIBjadjN70wwkR+/+
McwSzgV8ToxaANKPXOoOPrkXyFp5qZLij7Ij/06Yz13nr92HTkp+716bvNU1dYdbg7pgiASxggCj
2QZsxkvIaGeW+crOVaF9PxB/QQqNSDenoHCrnkEOjg6DbHoulmDc3DhxewgH4zSqKMpkaO9UNFrI
qxv7LlYfTHmRp2Sx5zIKTy/Se2QCqDdfYE61R6BqNOzJxaRZLHEA563t9Z4G5QGxqf/1OYkPRVmY
erQ6KZqoPTs2/MePagQVJxoK5X7YtG5nWI1fQ/6eo7o6I2wH2Tm54nkXJCCrzuLnDQX7p+07bCZM
05LDBhb45IhVo7NWZ6oYV5ZdXx59NiJ9Gk0b27pUaEgwri/kalGYMMSQ+97SpIE3dmSmEOzKWKxl
NPZZMdCNq6wa72ijpfmlmnziCkSmUSJ48vzfXBwFdoLgQPHmbe8eFrNMKhpEp66y/5P0orDsxIuV
mEpDhT0nDyORZ9msDzhuYj/+xd/xfsiQQ4X7D9vTPRi8FHvyEnQH3jFS1O+Hss/P9VlZy4H2J+bO
ySLk175jtNb00vPuYoNf94CwCY6xQzob2Nfh2igA/qezA+0gW3KV4UpW6DBsjpiIyb2T7Ey15mf/
siazQrrMCw9goAubfymMqPzQH3E/F8VfyHngJebOQZHVHf38ocI1Cr6n1WcB/LkQCNAZ9uOXerEo
AueuKM1m0M8KkwwCiNYk+R34D/zq98SKcUl/0V6EHkcVvPZ7aVt4bQ/uNCamLInjFf9U8KZUquTC
Iiew3gKA58joK+926GCHA860LcL8ztzLJCo7rqW8WSs+NDt0diF0QGRNu/pADo7TAUvv7F1oxKu7
ccFnPFD+YyA6zTXQ8ZBGXEvi4j88QeCVNj+8juWxzNjZVuwaLbFtJtF8R5ZXuidfIgAwlt2JocSK
bFUq0zwa3y9aCkVbYVBLBW0AE5CeN7iTi+aRHLkcvfD569E0fIbb8mrTGJZX2qbB6GzEcw/6xXYy
0h/oftS5zbHJ5H70O5KSV0opv7kLATTmLTCa8c4CskZjCTy/AHl3w7GhuklXetc97mjOF72eqrFS
UwG8kZjcBqokbSBKNlREhnXeVgGO76YlHDbCLeVhDQqT5ZAHVZ6TZp0oC/Lt7ezNJ0hy9fwVVuQ/
hQs2fan17HIAW5knjNNlcHS6l1/qohQQ9HIrh7y+qPtPpDs7sXqQqnb3nqmkLW+6tMyimZv4jG7N
//MnqPAgWL25qZ94ba4wnFN0mSbOY2fYUaNuvq3zaUTPqHr/NKkNqdybKt5SAiSp4bPCOB6WxAfu
iEx/8jlwM/eNGE1dGOq2Y0QL/loRX1991mn84j80D2zg/wqpZlh73lV6kCFKeCwag48SJMXy/kU1
gw6GKig/WoBewq4hUsknVVee8CJ3mnvYEWWmIRuqdssc0SkH2MH3l1W/5nNYGSrp6wVSijJT+c+B
8yO7kX0AhLrLaIrOLPgCG3XPpBkIMPosR5Lk4PTbfiNwdO3vin/aCIf6QmlhjqM7ZQ9Ilm5v31UI
iqNDdBCdG53SM2L5nj2AlAstConhTmWFT7udNmD3vN3lrEZ5pRFodUZ5VEjxrhAUVsZ8CLJ5bzvO
5QVEvDdvGBCcbQyTYgYyXMo6UX+lsQEnA9+5gWMBGYEd0VLpg3o8Zbo1+jt+adUZf2Bdj+9XOvkC
FXSD67La+4iLmJpCnax2OtC0W8iTG9lX9FtGyRWmjilN7Jn2tjKMOgpdjABhyee9uAfwtQYaohmc
f8Y56jiKPP64bmmB4EwZ0LhdAC3jmDT//MDkAYLWQTAlr5c1+9+006P1AiQPu9UdN/ccgtF9g6af
N9JN8yz+iRf5HB6fT17mIBqOYVkK4Omdws2qGT/kV12uNEzvEayd+dIgISrVv+8KPw8BJlbDgTQz
d8BZVru+EGHq5qWA/rF22XB3H208WSwwJehI+v1JiVDPEE6+1nY6jYzs9whkAGPOW//SmU5bV7sh
WFCbYSVjkirMdH1XbuR6/Zst8UnWGYzM5CuHxVSLjdSQ7sbb2SjSyVwTmRQLfkS6ZEOK0bfRpmlw
HuUSi7dPBGttv7vQLDbLy6muQqn06BHyeDfA40z2AV4clAk4Onk/FrDeUUb3l3sjqLJ/ZOw+MU3B
DMlC8a/IsBKD6sOYtm3a8KAW6unxZG1GSPNrwR+P9vjazTtna4Ud/NbP2P4IbK1CDKH5ppCbzRVI
G3Vrvs2YI5AMNqddksuZvkmK4E3Au1SaQ1jEfYNCi48oSwWD8SKYj++4YRRx4ZxeLONNMok8oA2y
9TAAS2EBhxvPl/f9QdJa/J1CYgzRRnMoCaRaxszTi+uc7PdnjykkFVNszrNi1m89zSqywlxaQPb7
rociad9QE5HmSba+NQG4IikUjrb5OOVu7X3Wll3E/I6PZzsO22mRsoi/pkip6b20s1ase/Mr3XLw
WsVyDomjju9DjFsEnJjYgWMmfQQxzdUDXALnNLHqgWoHHiJQBS79//zNoiYLLYQvqDJAMeUXOSV1
o2qtW8VvCwxyomu9G/PaKqn7gNotop/9FbH/KQ3/9/LSidMRAbINxOIOGorRxpnpbzct31ofSw75
gJZT22vBXkVmRLiP/wG6t9Tx2rix5boAnrNGolOue3eG0FgeQl5tOEYChlUukN7YuXEelzTYeYkl
4IPth+Eshsc8zISB+naezOK35rsbQ4ILMFFES7OzqMddKr5mKXoI5Ea7PJ4tabpMi2pGC7PEjkJy
Svj66LXQEmkQgbSC3+aF06HkdqX6jYEjm8+1BYF96IRvP6oq7sZhe7c51tM7MmfpxVRlx1HJROp+
tKV6pngfDx8EJMSO/ZYePxP7A7ghEX6lW2UzmcDzT1hgFXmAv7DW1vbe4GQZDgch1uUhqckcIAvH
M/NbHpwDIpyZRLLcH5gWu3auagp633fwBRmIW7Rm0Q2IbOUdl2l6AK9xOCk/LTSpS9rwqAwyKTrf
C9Om92q85LSiGVnf1rsZWVuOwPvbDMzj/rKkGi88cYWGJ86xpJzTorfYXMK2jKeWE6xzmCbf9uMk
wM9c/74+kvOeSpfK3oCr28p7/Qf7mCmwZqgPzDrUUYLCsEs7ddTJyPgdqHCyR18lKk0wO3giMdPf
CY537h1KssPji3WoLn53TjJx6gP+6s//qsn0vxqXF8oR7t3+xy7GrFHthWCssZl5v0DQg5R4gZKY
h9HH4Ya/FSzw1Fq5gqeokzcv3i+YNPomndlTsu34gJgs8FVcbM0H1v7yHMEYeQbxh53o4WxvU3C2
VVZVzo1LRj3bDoilyAfSCjWBp4kQwuNHModZ8FS1WpQzNgTZeyD/P5DERhVsDn8VI8e7JiI73P6U
aqfR++QSVSq1L6FVXuH5KzSnbxYV5vSGjWEzDvi3DjL80cUAZHblcn1gvY8I8iJ1GGAejm8LF+t6
4wvjKzsQ9G5Pr4n6I8+yAyJSYT7vBO7mnBMqwaDAU5ePh2yMBJLESZY0gkdhjUmGMdfiPaoxl8++
hhPpwV+6vBJF2vz8F2afm060g9S13f/Ex7MB+3tq6kklVXVNJvsHzDsxy0b3cdNOkfKln7D9v/wp
iu0I1VnPHSSo80rpJh1MaNRiEW26QoGTMt90wtp+Vwu4kNCIBhHLrn01E3SmE3ZT81qGRUKvzPUj
k4931oaYrE8mhdjRDJblE540l0lE5vT6pZjOwgWrobuz5MFBCNJ60+Qkw3rpL2bO3pgEPe0+NFKz
NyoebdrYOCcmwlZR313nDUbZnfacufdn03+/uOb+JKH7/PX1eROCNGw09pJyFpuO+n/yFPIYQ0e1
+PhSOHZFTw3yjq9rtccDu3zETUEG75Cqgy36qx2Fb8jzggX9/7m9E5pDbKpMUgvkfypaLlHzY9p7
DiYAvZBmnneOWILJSORXcCOZioPNpV9XDYYFmTytMa7ZJnvYjToJ+sRCzI8OnxoJhB+196JlhzXU
J0/9MckBCT17Z33FvtALPYPSWOdoEAqpqaXrvi29fA+O0Ku0xHkicpYVBZJd+djnkXbKsJEU+XCc
KpfZSS6bsd5ljuNr1qouRLccJmPJOM+G/x/pQwB+skxIjjNf7YRRTYMxGl4KDZqaknyTv6C4SQjP
BbaD+H+gXQ1hg6X/4tdRDmkt1wOvxy+wJr3Wt/lkKaunXBXa9uiTatNjv7nRN+9OoUCxULl4EaDW
M7SHoNKtNtF8s+wZ2oUFUTFShox+pLgDHfAIzJbZHg+2faJU8ZmBpTTgh2Gf+qREAriO7RcCKea+
CTvs6tcSEd/laU//skck4iiIK7KXjfzmHrejipDJgAHKYges3YzhIZRyDD33WBtCZhguD9U+TSET
CEbyS0J1qdQT6Mloy4t07NmiR7r3FxdoLVUKw9K/aQeL97qE9GJLEMhgJv9xMnqBv2UGLMz5fj9E
2h3lsgA/iNxHAPYaIM65fYlKQcmcw4yp2CtefZ1KqYAnPpWp9qdVM2jVHtAEDBA7vyWYRv40KZ1c
XGxgG5RtPVAcSQLa4JFsLP4Ns1OCGU9nk95+MWTxvIk5BmDYFLBUEbLmzq4l6wJ/5Qd2bpC1spKI
WElqaPVU/PJ2HUhefe4e3r/cGSeA+iV8y/0cdASRsPpzXL5GvJv5oEsFI6/4858KkJkDhvxgSzez
gSYZ5/ztZCxUBd7JaNf/UiWKT2xr8vhzbwMj/QFNu44X79KHPnogDkf4iWH/1VbzISLwJdI0LUlU
B3MSxGbOtbu3c61ONB47hdiCewdGkkXZxPnAT7yilTGdjOB5wkqbIKBQJX5vXzdzLO/TxXnasKzc
GMQ4opKBeJQiv7HOzo/UbQgVwjVcr6gaKjN8hWnUmyG+VgEZ8CgSFGIHYLG8WkW57bk3DxQKRJTA
0HzAVtRn0SHypa6+Eivd1Q1y3RVAM56fqdjZZP6gSA6rPY0qBcd9jHMQVI4myYVwGTjbYZSGgkeC
rZsi+Adfs74uNMoflsSlxDuhWoBVbrltgVsewbLlrrC6kZbWxmABuKI7XmJEarMGG2Y6Z1qNE59d
9wnYbxKlYod2YKiq4OadlxuXRdsYOVLpFUDUUq9o8nG9wZsJb7FIYlBJJHFXbPnvOFhgLttdUTL5
S31kGYQE2mjJgkRSvanbIpw/A17h5nfzehHS5rr6cB8eJ68PIAVXem6igSPZ9B+HKC2axOVZtlRt
LeEZg6RpcoujY6L+YPpf+AXErrQohaaLv14V0IXR3yQyXnOLYVOkOmCOmiiFXsJlH+CfMp6IfyUp
TqPJqbSKeZ96QyP0PJ3srImT1Nv0gltsVnUFxRSiGveOzkdS3kcA91c3QEhdi6ggWpqc1zeEulum
ARaEWGeZ0hLSlxMjFIoPZQlOTObMqKOWdRQ7DV5bbdBmvEvAJjib+kAxD2e62wq4lrKpdmTgAJ2Q
7kex38u/xHiQOqoF384J1j+OpzhkQhr1EBMBtGyjjFexnPMHlOIA4qp85mdO6BLOk7wOfx6M4QJ/
rTYH9e7Fc+PLW1wJzDiKd5iw3MxhSmwtT2vbqo4cUgQALuXOtwBzQ7aImBFDq8VThROJcaBuowjN
ziBYM1YomICiH1R7S4GsbC0NFkPxOrNntR0DlND7eOQP9K6WsXTGj9WCXRhgOQ08HebXHhKOIg8a
4mzRJEXTTu4GUeBRn9hcj/wei7ebFtegYta+zrYsLCTErds7NTJGvynhKb0LY113JKuBhq5/FsxI
Qq75/4f9TcTpAPmcURK03Js06ztNB23LzGZUUlIoBjFHaV5q0GmuYQ0o7j/CZazvIyvXPjSAGD13
4rhmCtv12J39rF16KoUQr/DcTedFAIJcB/pXXWoLkoGDCpWpMNGpbvETLV+sPVVs9bsBIX7wieKH
436wGN65+plLCP1ZBXUgLAxcQIy1Ylul0TP5zXK+PyKHaExhK8VZud8cjzkabCcvAHW00B+aaDAw
FQlKak6SHYJf6UVVFLLMp7vG8vOdaVkmDcBmKrhdjbJr2vG5q93WWPJp0rKhUtrntYjnWffAVUE2
fo7ZYbKkJ34fvXomBKsV5bfN9No1wSlipkQY+pd/IE2dDXdTA8EgcuaZkYIl5NXFbIdoS6MIdjzC
XxryNft/uzEYvA+6nCfrx7BG415+HAx7/ECb3Bos1Xui5xfEoiCxECnnpvD+ok9fCra0EJV0vSfh
tkqR+9D1DJvcW3GjGChehb9aiu3WyHnJl4Mo9ZShXM+X+fcCsONiKXIDRzeR044S9P8kqs6yStjD
yCXGE71eG/VK5aI2s40EzKEF61vZYybjTuNeBoT/znNQyQoIwez5NIMMY4/Gb9XtiBpSyPkFoTv0
B6DYeMVOKbsYRzudnIU4jKrRlk8v+FSCwwpOCt8CrEBTtTELyKosJp7zwajyVUXnHxtQ/ZoPGOVS
Z0He15GH3XdnLMyXTQQUVsLTCTW8tnyfEOQ+ATFkkIrwxkyhJC73pdlFGiUG75ulPj/ePV6Kuj9Q
443T8JKNPwz+9fZfZJcazOf1j4+Zs9h7UzZ6iD0od+7qEqaEZ/rDGejbBsE8qnycBgOLDgQhm9VH
B78SKMT4gc5W4B8wIfuEBXMt27JqaHOdPObVXmP35yMfG8bJPOeX9XWxnSL/vHEJV2PVahLbwZ2H
czThZ8V7eapJZAFvirpv2BXE4/DzPJOFlLAMFc68Ki9gJsfxHO+I8w8CXh98jU6YpVe/JJTKHfDN
ZI0fPZ1uiLcb8vsH246o1dIg6s0FVyszJQMx6ORtJ8T+sgL6v1PfsgUwh9p76iTG58dHNIatHfXA
SmyHNx62trdW73H2U3PWaqYSuodXqYE1Su2Gza0dPbTCcxSZLhTMcYTqf9c8iTxns+BG7G0hLMXe
9aCd0810DfXKKGoMGlgNDm9+IN20cR1ZhrTP14pyoU/U5/bZfPHCPVa32yxtavnB2CI8kUfccUKw
2eSwTq2uJ5N5TeseVcTkR0U05hO6ES+PtkxPo4RqsnfeQTeja9E55b12Qu2JNlCq5OJeAgW5QKOM
RHwAkKORfMB52Fc0+MpWev19Y2oj8dfkj+saEkTEcGra9/CkMT52zFAot7KpovPm0ruBoxyDEUkT
9wiBfslnvDjyraa1CQ4cQoiqU5d5my6UPf7e0/g+qeK2izjJ3OG2s3VVCeR0mUCJzUBUTODmKtbQ
UfZTc/O3DoMz0YA6opC5XoLemuDI0EzAglk3FABcxbOVo8W1SL4o37sVzuj8SOsnkrsujfdsu54N
YxLJAglX4Deb8yz1UU5x+zKg9oCR2EJkc2KrSBKnXeu2tXwku1wMQRr7ROmGMW8HSWF3Sjm7UPP2
Vh9cdph1QraE2O355Wtm8T4NED67FBJCMT2rmvcOJGY4QE1mFCVy4jw53ox/xMX1zPTCuNgOjmWr
igVVjCYkaX9yIYPmtgdYBrhLm/Uo0NL0DkqQwP5Su4TekC4GPrj+xFetrM7uVFdSyClFm/zqZEzG
lAeBzdSvLaJAt+R4hxRG1RWlrUhOZ3xuv222eMAAmUFaomyphgWEK2RYLU6uVGSlMOE/6btRWS7W
JfZC3fQ4NX+qBR+CrDiJ6DufmUycXkkpl0eRDBwGSYdjNy5XADY0FgKv9XEsJ4VtsbAa4CM0wjNt
MxdQMAKXc+V7UF+z/YlxVrSSnbyEKofOudPEA+M+JIBqObM25lmAzYl2fF3n+oDOBbdHCRsZ45ir
2k9An8+tS2cfXQmmpTzpl6WtQ6VF9XOWTe3Baf0DfvodRs7HDt2a4rkgVo5H2aCBVXaM51d1C9cm
8aLD6TzSpbqPCsAmtHNjynF65zv9Mqp0Xv5K4qsAp/cQ1FMMfOdpgS2twj7ospzziv66eDlxGhud
CufjHiWuRLPxQfZcOGlHBOc7LlwQWPEoCWO8w/5/HeHOck+POS9eeHmcJ0S0SKhyqeisdeUJ8EHJ
cVe2rcUurj6BI3ub/JFCDAlM+jvSa0SO0ZyJ2FUGemXUnvG+hF/orqL+t7w6bQPSwM86IEnBDmpv
mIB4LrH+hZMYrIMQh0uXtvFiBKdF9ck+XrtMbmEGw2BMdXK7RIhSbwvB5eUJXQs63oPj65MDmprC
sz/pzCLx0yyiMUi8verNkvZ6kjJbhimvc/sgnNPu1voSISKs2ZUqVEo4PzeiCgW6dOzrCr08Z4dM
wPvh3YkCeFCmLEcOlBfDaU29tykGxM0Mm+Ae2jNmcQTwDCcRuQ9Qy+VpSe+TpG+roomAhlYdPXcK
/Gfjgcv6tquCb1x8ud6m94ATCqWcbzDs6wLtsi3t5OOq2mSunQkiqPYZvoz8dBzdgjq3ThcykK5v
HY71EXDlsVTGeGbknYzgFB89Pkz6RW8dcRqbszmIfW5v6oTD3NCu11yM0Emdl7fF3lwc5JmKbx6R
URlA/URmgnVK4yhqDT9J6RP4kFCI2PgM7PzRIcYATNGCM35ITv+ApfvHqtkWbOUK7uQTVYpqP+km
clX1oCrq8k0Xoqj7hH4qpk48zGKRYPFmomdHeTRJH2NcmblYezqSejLXNB2GOt1iWknLwlLxrt4M
gDN75z7QvHxnZ/nSoxf/Np7deQk0Mkv1QXPMhyDc5rP1DUXKIeYZtM9/Sq//oBVdrXHl7Ui/I1s7
bJMsNYh61qSseKEV+1dT2uMGpvNMQ0/5k3EwGrZkuPh7mvj8vYQUcDEKFa0oE9L2SnVSiKSfJaaX
QbnZj8vg4YBpJBhzh90CPHqOdHJEIXqvXDgSPavac1ekLZmDQVnloLJ/T8x3NdT1r9JTSX8C6GX2
GP3H+uzk2fS/WjHrnB5ccm4FyIfgorxkdFt5UwvJ1BKOfEPqYSWr6Ze/V1soL7UTUttGqn1iTXfj
qF5zVG8SAhwrDxLr8xySigldmCtP2n6x1wO0DtKDo+5hOj+7i2b+bp/XmvxjlqHBVol7uPVPRzAI
gHsuKp6K1LBUQ6oGodbBh5n5k5TTGxFnBZK0GhhqI6CUZAxJoPMjg4Y0ENZ1g2DKnwIH0OFOmlYI
a2dSmGRfuLD/CqHmU+l+JAKVhtEOWGJ3FWy6Uiz6BT2EGZHpZzcLXjCSlMrVbNHVX3CWRxPPDtL9
Isqi3z1BX8nRPUc2omoLh9RqTWdVuNQTv7MPKEjPDbAzpBSMmQIrONI90DTmyt90323ILkrNsLsh
GkXppYDVQSu6FjAMDye88P47dApyl+j15Uc9FQ/YjOvIvX6enoPdMcdBzJu03g6NQ+c852zwWYcX
xE5CuyBjpN8Xnuzb6YUF+dzKty9XbG/l7IkGnKayJnhipLBarsExRIj3bPiw8SLhVdO/MkLfUgXL
G4wSTA/aXXr/oXn5cUJpkHZfa9xH4klaXBh4rZ5G9aRpLWy6QdztD80ljE52hKkqg5giGrop2Lf3
SHJweCS2FjmcQ1/hpPKbWgeLZdy/Uh//VaxpP7rmUliNLcS6mh4lnvpLqt33Zb7rfAhhEvkIzjDJ
h7M8S3+BAGUSTvJStMOkA8oP5jZfTEm5uwWfAvZA8ww8K9BWtONdeW01W/NT7ApOyg1CZwHPYXkn
2OLsPreqY7TAurDb/JjZzT/TqduCW4hTabDUxc0uOh5HpP1KmvNDnHoMwY91kjgbA4E9SllfXVLx
E6uDO6uMzJkEyg8nSW4e4CQqeNRlQQx209yMN8EXkF+rqX3xOxZDw7VU2Bw49NygFhgABsaO4K09
yz2YLDw02peeadiBBUfdTpBDXfrc3G1Ib0PEpqe1jkG43hhKwPrxYmKkaSjZwV0IOPOpqauzkNNL
1/odOwGnPyWwMgKwxkvdOdfZ8qnKDq/K5l1vsjzswnqNKXVG9OUeE9RV4MH9mxMU8gFwi6wXaLrW
QAFSyARHEhQ6bD4F0buUOlz7ya+HRf7sQfeXGzi4BsRYCDTIL0hKKcv2br7Ct2LlwUeHAAZ7XSWo
1HJA8b5NUqSPYsqACq3Ii+cIX67PObANWo1CUhz/fI3zvSsWNInL+Mi3X/n7exrBtO+uSYcc4OoB
Apde2PT7rkHeaRYf2V/jyGJoOalE/g/rjR51zBe0eM6AlEq6qFBEAJoJnSgT6JeiOBGJTwHCIOsF
2qs2Tw+rvNZSw29fToFtpYZhYCs00uyYihse4X+O6Jy9G3XiYnCELCVqRWws5+xjGs5sOUjklYF9
TwqR3UE0swd2RyyAgnlk5FQkI3cn2t9vbp9gvsJoI2R+J3TW2dJ1sQlkudLuPWzGHKIw9uiLczN+
4zNUuJnG3m6pfS8fAkd+qboBJrgGEvQCiHmkyk72hRSa7uzunxqkzpW3rTrtE3AyYBW/GMiYrYBG
SnxB4YveI8N3eIkJj3ynv1UgJEa34AvzOCIGsulUWvsoCHCtX1HQtM41rm1Ox85WC+R5TrUIEPLR
jHfSPvwunFXa2BsCV9rwMqpfZrFT31Q2qFPSIaTJAW0iPavuAtYNAxMqcBy8gFkaCx1w0G/KEX8a
tQhz1pJR2PahLOtB2g20IgsdwOG0XiBJEMv7lA3Cua8qbxN2rAuhDOKXIM6x98bVvydzIKnPPg9/
USKKUXnImfedTJFNEux8d4pyI2al7b2o14Tp7kpq+5L3sGkG1e0DXt2Eti0wy1HRWRN00tMQkXeO
mXQi86snSMeUtQT7lRsBYjNWw5/KHfmvejtf8CUJemzMjHjfyfczMFAQIOB5Mj92ZGWhyqsU0i6J
V7AkKtWU49H/u87IGYAJHs7mxrjF3YBYNeREK1IjwLDwiHkDA14fOCe126tZeIxBrS3MAJuSC6C6
IiDfxwoK5rfwzLkM1L6ftGZNuMyaGFmDiWA0Kl+tUKJCQjhyW46UwVNgBM6Dofqpa+MNUD/ACnoI
slcZ+ghzwBtSXWuBMBvIFTfWRHnIAWM8M5RQ7MAkt/8bBFPRDj3mQ0lMmDbCM455eTtJpsLjxr7+
t08vjiBRcgSbY+D2rWM3kzTbtukAFlEzVZ33HVJiuo6m97eJIiFELY+4GExPPrwvYGCziDggH2xy
mXb71U2CV4VZt5fPuhsM9q/jddozmMiIE/FGs67BvaUBUxAdw/igNSC3YJVtGdKahRDHpLUKTxZ2
DsRYyZT3OU3VrMOC+DB5H/HgRPXdfMlNweU7kFeYPQOydft1B237Dn7EuuJPSgWP7xq8rA9HcFBj
RHx34Sn/RmC5n1mt0im76sh5bFMbW8yaKzWyBsCjpqggUe7lxgUDgpwmNORrzHa1yM9GDeRDyIw6
CCYLaRgX6cbv3tQlKI70cBoolbVSpk42C1ia3/UrOOhmDmSnOgyd4vUCex4liKi5An18uP4Sv+GM
FQ2Lc75EbhbHpVxCkSZpI/BqDXb4fFIEnkAaYEwE3pD7VqbnKrwJJEr01EwQJtVVw+uLFMXxv/an
LrAGTYCMbrMwGNNUmo/DjjtIuLvR0VXh3dOsnD5bjhpfGC25xNDmY+3XfdbYSrNDmzYAtItHrkCd
5iWIuacLSqhXyz51/JDS3ZEVtxHFSYQXqZZpUATdNPCujbGTb7lPwLP3kC9LXo642jB7darxr4f3
tMWBVv/jmIdl9ZfrhrLi6Xt3K7a8s46zK6TEG5cVM+JsfZ+Hnr5lKlmdKTxIeWaSWDbjGfK0D3O1
9QXHD0Nr/lEPk59zNTpDOYQ9K4+Jg6qz3PVaXCLKyKxetuUnrFW57ypGEbsGIyr2HfccpDweYvk3
E18r3sdsndiW5rekq96CzRacOAk6ZIE/SyMrHTbzOAM+Y4oZ2dFlQ2z6AUGt0Qm74KHLZZTPYg8m
HSZZOHf79zm3yDpfqaDm8uSrtcsKmfimGBFo6WrtyNVEz0NTLqSPxUQN6Vvm4UIyvUwhCgdhuKs3
6lwINBttuhIMVvpSDLSIjxsGj32EcHsio/R4ukp8HZu6PMj1Q0r8XAjyuWuitO5RQtMa7o3OG5rB
nP50KdVvklPLFEok5fTHH8vj9kVPdmyUU9IvGCWMWB0skalyU8ZkGg1+MeYKxu18ERpPMJ0wHQnq
laJWTrtBGgvCpxPDRCSkq8A61VPRryJRzTPC8xb7ycStWUWsHlbkMx+A0ay3uTTw27TYGDUjCamn
RsBzsu3rZf9uo4P2ctjxlqZzKeP79jwLP0Pt5xTrBeCAZVuar2l/6THWxdyXbOla0EmDbQDcPElS
Pqyvp+2ViiiABb6CoQOiIQ0GepMWa9dZvpolW1CCkuunTvGNirOaLs08IdbBLkt6bwMFNSfP+J3g
WBOBIbQMXE6CoDwi128G59aEq5WCzhZaAQicGG7kKuyqg2236jStAmLYLQklKfXkR+4INUqFwzPX
slxOV2UT926b/fKwC3WDIjNNbjbt2HXD+3/YKda/etraahcQjE17QIcX3hXOV2FFxik0arCt/q+D
j213RUNWQpf9jBRPfFDVInnlWebSwvnJBgI3498RWlLAi2RCygjco3gQ38yTkhTNJL3AV74avzjt
yhjRaukk7mkITogvOSPdZCwpPfLyjX3C9brpl8x5COYev1ZAvMFvbyfGf03CM5Ov1nxJAGfK2Tdi
OZCzqWMRyXuGNocne692om80bju5e6NCADb3+ZuhDRBtF3qWsSZrgr7LhXoCYQg5GWg3tNCmjLio
MaUhLNYTLyIjcmIuZGOeyF4caoWap41KRwi5EF8G68SkRQXzLYk5jMKBrdssAvxSfJqGKT/XvFyP
+tdqw06y1YnveHl1VAGOR1No9YcX2qDfrmNf7gdOM2Zj8BxI6ndohmP2FJsU3gV3Cyf64yuVu0F1
Dzd0Wq3JwkYJNeVOsv+AnqQZOr1jH919B706D/1XV5BOhDp729p09811uEGXuKW/vU3agULE9lO2
6QC0Ot28kTDzyBpL0loXGbQy1xmb32Hsw9drMGBwrqUhnM0QmyySWFq9vjMMoqoJPZXWgBesE4qY
iXlFF4mNhZGgY1f8BslTBkAU3+y2QjxD/2rvLDjeUtLyQ5zNOJ56CsNScdHiTz03niYET/KxyDPc
P0MFKP2LWul5GWhIdG6ibMJVW/AuIhuchw39JEu3yT3DGk1e8Rwsp5qVb7/Y46BIVlDkk7NtYR8B
G3IQy7hXhcefqX7LdL8lQ1QN1xParJZve1lJ07Qb9aa0DMPZwt3JuQzgJ6CYbiFcjU13QiEN2nVG
wqL8Ves8KhjUTHj3dqRLpW1LFvladZhAk9WEEdXLwkA6WepwZRnYbMWRiRZTB4sc803ytoTie11P
b2c5dVdIl/vqWU5SQqXcU3DQv2zV3x1vFuI3otW44pX6sJJSQnHjyWrANUsqFS2Z0aMxLi122O/T
D1TkDIZ0ZVSNWYn8zkgW9AWv2p/tCkswYu4jFcnKo9ORCB/ZC6C3YUjiQtzHEPJlW2mgA9Q+WccG
hrWcAnZH2JePDMvC7ndrWnU+aV4d29azIBTwwUZCXxvq1XPgbUG2yiwqolv7ESdXGAylQWJpOzqi
voRfl1OHIsqXDqbK/p6afQs6riMGwZRV3gJDgGgkHKsjAW/TPfaqQ4KGPcKsAS4LUz2hXkAdVc73
HebXfkWOHUrBQFjcvIdUY0ITzRO9+ZIucgXneEMHjl4GU/y8MEOoaJNM7fyek68KWwQpyRd7bT/y
IVbIHSstKSxdXdaGXyiiJIgyW+mg4j1ndBiYVBJGldztKKsoIJiuTNzaiGmL4eakRZ4YuVBX3KZz
+Whxa+goHgcxRzAtP3Q1FIZLNT6pRuA5QiWhbx9KZHfVpmED5cXCtfdckcQzwk+RgIJPrRRBQayG
ujwbBrYvvEiLQp+ieshAfBkVHMnh17SOy7upGnyhqgoAGoVCfa/mSkd0Blw1cKpSWUVathFFHP10
tVmLXu5Fq1RJyogG7nq78oFH6xX37CaTRYSaelv113uEi0B+Q0GzDE9rrXpTG4TIkb+kirNA00zX
CtfPkAiEogZqBedgyEGTiLd7t/SlUsuGjJJKUPnQ+5xmw1z7c4gTakmyxZbDPu3EP1Aa/5DA7xCr
lh5/7LS5Lks5Uh4rHTxXRyepSA16suWx8pXwFTHdcSwRiMpM36JKwD1iuZ3dTT4ofVHwMCdWuggF
FdQWEB2WOMhT0g/AWIfVxGLtWdZ2qC3/+AbXs5SsTGEG569Mror/1VAGxw5IKVafBY22rJqKN/9r
Qh81ZzXWMod4+7oSds7G0AwsDci6JtQxHKSej9O2UtJT94CROXIg7OujzmZuZKUFzYdn2IqL3vRj
Ev/edem7KaDOBeO2v0owC+8PBRw6growwH/uhghprYLC2u3KMuCYnu1+W6Sy9M2krhebpuBWhUNj
HsLsW/bSeir9WZyVa0uXZ6xB9TQzAtYthbMF9v+25XDnKZUUj2azjepTFkpBlaRhO04VCrMu5G9T
ygYoI8ltSeQRKjW2001voiBzN/OVO8kNU8+l0VYgfXLg3eyurAGQGbCSTv1xflDFGJBfINKNbVqp
vddZQjet8hsYr+sBa3p1jE2+L71JeFYWpGG54fQHhfClFIoXM6JKveW183lLlZ5eL2bgYQ5IGcHK
o4MP87ce39pR8k2sV95757TtmIke0NGj+hgO6eqDzTlu0FVJZnGnZ+P72xtYNhTzfwEjtl4jhHsP
2kg0ycIeLV3Dx2GKvI8aOlxh2idv1Ik9jrHpgNYmQ28lyzCmzxz6QO60872c/C4Pgo5B6h0gwEOR
yHxcGKusUegek0gfxCfwx3sBIIvdNx62QLDRK/hTbcoAhXhw9vS6yhX8d+ma8/qEHj9c3PpvdRsi
+MVbT9cM52YOcDiHB8Up1ozv5Yva9dCywN2VKABmTBzDWxa5aBNhQEqruhW+ZuPIsux41XKWv3Rt
3TeKCRkk0VSNpZ+4HkfsF6oNbfbkywleKhaRlIQqb0Ji3rXw7w7nraLgp/hRoTZIujyHLvHDJpRs
sBbdc47bx/A7lBGhtVs4Y9Dl+C2CTklz0Srcfzlaox6oaC5lVFrl7Duso8ZDp2a2AQqMp+mTFCl7
yZKWQhT+EUk2cXnjmN7t6+L6BrYhKYz9G8phP1rCvbVXM7vAP4DzZRriudc8+04NFdFQH7wzUEQ8
OXnLFQeTSqSUCqyz24qe3Y2eBfMEIRQYfUa7Y0lZGIs7dbwZp2ICGg/4IJwNlEQ3WDOGmSM962Kt
YlCpT48wB1ifrIS+jg5v1JHhOuCXOLYi/eDk6cRvKyCPvDd8Lj4bMCY/+sHYopbgphz0bcKV+tl9
xr2RBozI28Fcd6TBw4clRft3QDOE81RCZivzx+QF8Ex9OPxYZODMeW1tKD/7H6ZapUjp1w7jpjrL
dgG0t73afLGkbh/4fq5dk+7Q59zMyWa/HJoDrrq/1S4VEEUU62l792nR5NgZMwogU5Jcz9UT1SUW
Ok7cI9vQ2p40sgfpccdwLGITv8JqfxZjZoKmIZ7962xBzpMsAZZVGEFtHTXb097/M2ST8O9wLzvk
5TLIoeXz0EumDxj6itUvaqbi7dAAoGwU4RbMjutHfJOGmUg4whNzmZZMDgF5DErh7g/7nBVKwXSg
fzSd3mw1dAaaKjSuWCLUVhAf55bxf7s8xLu+kf/upmNiaD+9jLeNgT2CtFUPg7zWtGh6xJlRKEHt
Ay9ZK58DsGmYTHKld1kdUTeIrXiDRXTLnYkgl94dXhjBW675JnphnHQ1FN0GYiiAnkiSuNI/df1I
hve1/AFGrNN1guKoykpHHNsnJRpgvu42hksl6BGH+1hjme7difWYJRG5b1KNxit6+Ww7yfZfO0lc
7SO6pJhAO+xj7tIn87qh66qj2GLeZNPhCANXF4YJ4APS1ly+Uw7u9ssV0M/k7z2J+9xIDQUyBYJf
HN/SBkOLfDzNgp4owUwv3yVjaD717m9I+oD2Wsp2p9bm03/U1TsmIjIJY9G2ulxAz9O0icDs5+R0
YT+gIE2rCDv5ZEuH6eRsSb1lffZlg4Z5zQDxXcWqiJ7Vun3tCtdAHsL+epoCrfl0WwuPEG0oDySY
EH8dr9ZThiVRZ+ZuPRqeuB4kVL0zz0IbXJbS6qiwkbfUkkjebIgpvOCD6zixH1UIqg0X7l44I+Tq
5bpgvLpzMRsiPuAHJY9SL23wfChQpDKisH3o5TqdFV7RkhUS49bbsj1GH0zgoEc3X+Cn0DjXx4SP
xvMNwzK32bz6I7CswuQcnZDa7koZqlhRCspteqRVfqlKcbS5HUqgsvc8DqG/hF8ccAcg5sj1WkxV
rtOcn4Hv/vb6fuk92g6FHTQ4MC/9MGHrCN+bPzmWdFqngx2jyQcz+jG8/pW8flkS0tKhbFxyHeqn
7XizPLGwO+xP9kLQCeHqahltqQ/sq58NM0bIVvrbz1+YY2E2J1vw+Fwyz3xediT9gW9qonB5Cg+o
KWt2x+pFV8SPTr97aUv4+SO5iCFuT6cIsolmHQ6fPqt+nI4IeymA56Js6IhNrGJ8x5t+K7BG026F
NAyr33BWsGUxGhZKKGZTSBYoBOvN59A2r/Tm67f8omah1vpr8gIlKsz67GpdBv6fM0a8lW2P6bom
BD/6jdEMK9Sq5h6EF30U0BEf3I6eS8S3v4aO5BKUH7dvuYGfRgWM0g2sXlhq0+p0shukR4L+jw5a
JMadFFcioSr+AIllDIXdWB8et20GEkA3acp8lhN8VupMtnP2JTPkWzd4oYC2xlQfYt84t6MpyRct
W92DbhWNmZ2mPiKlL2nXbchDUGQKOt7C9YG4nv+KlJDuCdeMCPp67FxPRaBFTagvDZqnT2AwvG1G
J3lP3FE8PfMMIk10Bdw0E+i9kxcPVe0MLM4GkXPzbIC2F5axkaXWL3Shyx+CX7bKYqWuXbdexmvI
TVwdJJqonaYINSPWqcgfp1543POq3J1vBDvdo2olmJMOui1E548budrpc+vpIXeIhNmGo5o6URVO
XmwtwavlKF88FxsfQKPUBrK9a6xefxbZp+qo6KtltSAXQCisKwrvevK3qkwTFKGNzPKKNzkQ2RU6
3D8oK/XwOQsdEbGSMOi55tJj5zsm356uOPIQiprDgniV8fusbAGQOV9xY3KYYEpAFXCAZVWDTO+b
0XGawL+yrFYMfUtAiVPm4G8CyZUWd/b751FObDyJxur9fekS7Ipw7k72iKHI2r+PZRNbpsN6nv5y
5+M12aVtuLVRuh0aJDEiWh5lgml2uvHmEinWRF3IIZQkA0WZRIhMPQt9gGMLnfi0vVpnqcaEPbFO
3SLxQw7E2lI+TKbXMeYgPwNSY3lpCAJRPOswEKbIBA0argLgj7u0FkjcRxlPw88P+VWjqXvGAGkY
6GvYz5LhmXi53q3Cl/xM3+CElHWZLzs28jZypMDvPh9PjjjJz3o6S+SHEG7zLuwSsGsd9T9ekE9F
NGr79fBzY25yqywvTE6IaJJQA8EYvDThVc2thcCXibNCduUDb+QsKEdrtGLk769Eusy20k9zjfN1
VK216Rk32iNFuey33oA4QAsxGKX01LvGpSwJFsr9Gy9ODSFkwt9ThJ7h+GGx9FRnt7VGZhduA5Ys
rDFMPqguNAbfkCkZPIsGZUGQXrW+FEkoMvma1HLfImJRawno8jBPRMs3VefXDrA64p3BhQKoIoje
9VCOTIt5OV+f5YA5SKou7rlajvNgb7WHeWEo7y4rMCPN6TSuuVCVkDhaZbA1tXe1g+MIFGvDe+52
hd3OirT5+CdiQhgWXlWPPlpRd6oRIZjQFkvcJM2SfMNIpKnvT/I+P6KIFOPlwlZlhQVAnFt56+xY
ZG21zgkkKfmtd7fKfCHqrtqofvCUTx3JLI8wj8H0hbeB4jpoDSsKZRqFcsRoSoLHHgiFLv47BxYy
YTwGrhzLWSUggSXu8qqRH0NiF9lW+LoaVcJkWkw+6QzKWWykHcaxgZbBQfIxKSaQKRMv2/p5gAvh
2NXxT5pI78IN5L0S7yeksWtuZolcOh2bpHtS9wP8kOV8pQyiGZOmu9R1Ok/M2zh6kZUYJXh1nOhR
SzyelRHH/nto8rE/5kne11BLbylHzJPN2AEmW0x0P8ldZo5mtSVEEK30lTYcILzOglKCCdt98TSZ
Zg289OYr74lRoIReO+1sv0Hv8saTcUHaTdHMYicRJr5LB3mo+rMncOnSCnOgC+cbZZQWsxntKKYH
+FWtJQ1FR/lMk0LHsdgc7qH0xdmr5fvVmAyTlMraSSvGcz+4Y40+qiaweuM4oLqH49YigBOwUXFo
B5kw0hFeXs26HG9+vqOzkovB0F4i/X6sir/M9enXo11ME1wXov9z6uoEG8JDc034mpjn7JNs9wIi
GYySBjGSk1fbwLz9jTYSVrMLQO9ejBwZ1TdEvXaYY8Svzw0XDdwXKJ5Nkd1Kn3AcVGauVMl+Sjbm
QjgIcPBX4sd+Tf3xtg/mYZ+u/5vPxZ59GuYbJu2iymE4/sO/v8RUhkveXpHXCW9IzKl3NAyMcEEA
u0KERTc/lPAbQx8WiKBpInB2o3UNrQiEaYSxacCeN4w4sk6h5WzbwdGbZAs0/xbvxLrctsuE46nC
AfA4yr9vCJ3Q/MYow4TUew05Kz+i1MixzZegBentiEhAlnYkLrRCZpNawgN8weEDlbkn476OQOKJ
FDxrvU/X02FEtRyeLl+DjzOtuAnX4kcd8HwFr3rfwp6X+1/VzaI67Z10m+f/GFZEqOGT2QGyoghs
Yry2JggtuYhDNKwwr/oFdtly5RcpFVedpbTPjoWd1lcQBOa2uktf8/zqDw+isrOwMr9v1iO0SgDA
ItwtcbyEPxzhCnfElTMi57ixAnx2QMI2jM/j70Kfrrbmv5X45RmVuDMhOXwIf6bIL+0xpezAzXLN
QR/BOVtSG2OouBcb2oZogQ5cL8lXIbcZpNHdmJc/jQkruDL7CPOfOA53aFUfr/ByFd3gGBwIt9/n
IbNHKETr8Z/o1vUGQOw2NcCST16t/Xgv2V5WW1Qa/rF6Wdu7GGvqP6JTlyQ6Dixq/86OXgrQYVoq
o7Vi1D85JOxHtkyXBGrFkw1xLrNZL1qj3u5bTIIzJEF7J5Vqmo6XgoV+KKfU9KyLqhxKQl2+h5nF
BuYt3YgTNt4PoU5mh1OwA1nC+miZq1/fY7S1SzExePkBa0cnuXv5BRJ1ggpqtJQTk6CmJ8T0oz6c
AaXPOQRvp3HqpXE4+0UV9ZERZUH3rl63DJem+u7zElSYHErY5TmfhjJzVyLa4L4zw/179rd/sglK
APgde9woUaW87j7Un7j4T0Cb7xRGOzv9DVVBvjJkqcnQAK/gXk/jSjg/wp/Qc47sHGEwNpLtJWH3
Ol59Xi3dG+ttghvQ2g5kX3NxrDO2FI2dqI/H3V48+lsBW3vDR2dwc9dXQK6nECPFvEQUMkI1P9Dk
3zOh91INQxYENS1Gid+oU8fGX3KNtODGwrhTEVdChE4I9HjapmAxVZv62X2RR3xJ8UAwV5r8YY1U
Of3bnkH89ez4k6l+Hs7Dqk/wLS2N4eslaFu0z6fPugP9FNoHhrHyqM65VCtvW3uxtNPp3JQMMjCX
ZT6/CvXu2OOVgtn9exNljcOdxLTmLJnh8MrROTyxKFZWY3zBLaI2UXXKar55MM7Mdj+Q4npegBul
jnh1E6Ba0Uykw8eVWO5KmMbL7MzabJXA6a0bMwBJ0DwoIWVMHamjyfutgOfUTkkTzo+mg2AT3B6f
oyPzKuO1Q64koi8Z3zc/yEoUnw5Mo5e6lYdG6MtWR1N73+W6pTflmNydx5+thuPthKreVtsLT0W0
Gr9p1C2QRudxjKT/79mMIjtJil2weJwDQIFtm6BnFluCuCxXZGyYjZTs6UT7cNueklxTZTUoAOPZ
yhTA8fYa5Rkl87JNwe+l2CcOLCBNyby+g0iHl/vs3F66S4EXYkQaZK8jTZS4gA5yMeSj7gOZCwL4
81f9W8FlrSVfKkrxegQbkni8H+FOI2XeRmNlTul31FFdO8ReRpNUD616pFKeEvZySQziR0AWssEx
FhXdANLHWGFERbTpNcLzuZ3OIsmigeEAX3l65E06F4S0o/n5xQJ/UVzq6ynRu/5Ei6YRF7OWcbN8
uReC1Bv25P6Ebgj6V62UWyzS4C+wpocv4rhgkpg5RUFwyqdD8qucCUwQnZsDzUx+IdABTtT4KZuR
DLawLXg5LSzWpLKffhZ18hwpmqsxlprRLn6F+gUV7qg9OhEwX3hX3p45h2WgjWBqwGRmZqhVT8YS
NKRuKcyOvSmiVmdBRt4BPdp2JCF/v0EDLCo5kJU1XXElhKHHcDKCex3blQD8TNduNEqBl4yTA/HM
7X9VHuz7UePfPXKgtrj1HcV4bDABnqjKmqNzA3uXCAsHeoxbxdIeUrymFqP6eIPFR55Q+FsCgCpD
7lEW+wLGnVpMKl8Rqel8pUdKC5d0RomvSkVbZ1idb8pMD2Swx0BZY6/1Frh/xLgUcWwwjZMUTYZZ
aZqXVmBzkZZh/6+QZGd9SPfy4zZbRZkjLQd7qnweeN+tprC0uxp8j63/0jaBbFTWvXGUm5iAnJ8/
5Ci1oJZjDoEH3RlDuekG4u9mdN8PHWP7UGdcqKOg5w1ByP6EiqA9+HbaL7bamnstfpACcTGVRaQN
9YeKBpVXAj2D0Bw0wLXfLasrR9Y0KOZPD5DnKkaihrFw4fdqlUaDq+nT6E6fLIqdoFWKEg0wyhBx
lrG9W704MiTZ0raYOGoUvn119LLYdIHnkEcauOJFn03ItJzvPda2vJD5r+tzWCg4JBU2nQjYHs3N
WXJVEWIdGLoiYTNNJwh8gr5nGS5+K4YO11hyksfLzY3qk0FKGDmDsmOX2sy5MjxOtD/jbk+bfk1a
zHhwnYOARINGKZxwPDOqDUC/0n105HNFNLzKYCvqFM3UnDDZf+dEnWLy486pLZOiCM3wUANYcNy5
YpL8VJcILP6c7dS9PJdgvyv2bXODFF8cIUOTkCpB0phlJzNo2j4mKas4gP8V1P7TJ8j24yv0M1cc
6ekdpY1W7pklGfTeb7/a7WFzGXfforZHW8pWXrqNMhC183QRIxMi4fscgCa3ziLa294FyVLxUdkL
kPma/gmvm5ef9noXDGDL5GlFvws92yMcHpHHciJ47rH+bH66TUb0cw/bk2FHV0JpJ+XOawxyYlU/
OCbnbMOJ04q9uIokXI7EQf9iFjotiilhwpFmJ1PhQ312CmOL7ZkVdehrioBnSfAvmv10eOWd3XrJ
m65kdZ/D1PsncPOPPHgEA+gxMUePb6g6YAf1gba9IaEWdBvWmujWbMybJzum+4P9ZfjvHuwOcYB9
j+AG4hWMsfN5zv/bM1umdBCOfpp3z1F/EnqwzaCWJTpuO4rGcEOcSfbO8ZxA8wgbbHcgMzSlid4a
3BkvMKnd1mGADSXRbUiK72WkjqYzjtDDYRTSEujTvD2ykLKoZ3+XU6nOHZ3obA9VXzmqUwz9YiZV
vpgT/8xatNm1WljXn3OiKmAm04Z2LlwlDV/f3P+Fge+De9LEsxtF7mnFicfyRwoiQeVIUya/hp4r
4YBo+m6TrKial9wcrT1VZjZj6R+3mVNGvkZxBLD8bQSyvKBgiv+jrhC8eYIWMuriSrCgYvkMWznX
09yS4bKFVVpf4uqHrJDfys9VE3cbn1f+NRJiK4fH/+KbhYY+b6CN6c8mghAlqjb+y1ZWqEvUUEIw
BsW83yQu992T66O1kyRS6S5L4/hTAp2GvhneKjGCPek7ZEHQRbgrqmRd7uELW6vWvQTinvVMu07O
h/3h4RVy7SHQKa+TT8vqBynzVY2tURijq6OIFiFi52Mw/0byQl3uwzVZFp46wYpXPuMEAK0bPekj
poLINyxXu1kN6TRBmHIM+JTIHwc5upfq1nd+SUtFmfPXmWeHrFhhrbwUwdmlXD1EIIuuARp+NDCC
SBz63sy1wioBzb0vEFihYOxqFyW7xPC8sLUukga+gAMo1VwgT9TRz2q4cp1F7omfUVg95Rqrgbfe
DDR+nKFe1+qLf/R0Gx81NvFf3iwPcBKjmw2JtXrswHY4s8YHBwTS7yhQc9PkQzfKaOroAYyPu9nP
ZLkFekZrxJxb7HuCDwAaPvKn9WMWCRUvJ+6EWq6RT8tWI/LmnWkWcbxVInb+ok+wH222RhIWdnAV
qyvUCwzLKROf1zpM1P1zrtO4sAd0xkXuB3bQr1pKiYNg9FcTaopZXdSZCdtk1KXrhWGE4WVao0QO
YtxcIO4O+tJl5QxTniM8mmHbdnfsn+D2Dm9bNDFjhsIy4V25Q+IbJ3q0xi0lsOJmAA1srRT9L/zk
SmVFG+y9f7FbwFeeGkuFgIGJDmMCsKBXPMdbFBvHo3q8XNVN3Mt6Wit+1ba8NmbIuB9h/RwKEtIv
s8Td32DfSK+6OvMGmWgbtoWrClhGTFW2FyN26c29tSOT93jmZbvA9BnPYr/k6Lvtena/kL5aG5U+
tkWc+nXRZ/cbyLxLGaplXQs1G8y4KAo4e3Vf9bzGA1sjNI2fxeVcx4Dx309GY1PUa8KyctqNqukg
HExFLkZSyCaApExKBYey1IIRSiQlYyasDihKTSptmBjL9ZEA8XCRhksytwZBR7F/MEUKPP6x8oyv
Z7w/2Yq61ka9N+kN+66lt8cSKVrG9+i5O4CnnwVFzwrQfRpUCMEhNQo4yKIaSMb5PXNNKTOrQP7P
sp+ATSP7MZ8h5zzMbDeXvv25ljtnJXz25qy3wvO3ZRmbKNt10U+NHTojLr1kyZZezVHSHCnmQ+J0
r0+bAsEN2paGFYpeMJFYqgufZunAZvQ0q5KE45+7H6AeaqylKc8CCbRRL0gUhoHPYfuPlpqLGaEm
VeSCMCEOR3Kdjeo8M9DJPi+IPO2P8AMv7fFdZWSsEhxiqHmKVl7SMEY6yI1IaiW4h7p5pMKxH8qX
0o2XNWSj0oL465kkdY/UWlELeapsrhcdJba1mb1DPTaze+fpFwL4asN6+miTlss8WrEvr/EHG0dG
L4H2dHGaOmeko9R8w24bUQhuvzkCHDptKGqNvw0wC81Ta26eYJfgm00vUQBFa/MkufhrYD8milJd
vpiALu1ti+urIxF3RyLgVGjJHiHzPq5e4f3lmSmdCa+8x+JCI0SWjEY9SxaXnr+sMxC62D8LlImz
BSNfAOMoHm5hsGggwj5vzV60SaTlTXYQUIlQgwViPqBcoDMHTj2OHQ/Pr1OAit8EvWZPuE7epMC7
bZe0XoMCZBl97LmJayyNPxku8EY+Gp2AxBKhRFhoDjy2oc6qlrQzo0PTt5PX0DIatxuswl+f3V1b
aUKzrXY9YJDsUjGCesJpNyHG4mC8hLaW1KijoYU6mAP9ctOsWdq4OLdkwiS7nXDxEU21wD67uTFN
jkaQ4d11ofkrj9t+fiFqBTBc8SgvDDpQ+YvyuQBxOreWVB38Z0rWCifEXKuk8jXv4m4Fr8RJIuKT
WW8Fsx6Dylu7W7g/UsLU5VVt5+9rIYOsZrsnDWoTDe3YQbBiAGsyQV+BMOGU5LSsMaN7Du/RrQ4R
7Zdd8TaOXI18ZGiJz3c/Pa1YRYuTLonCIl19lpMr+yuS+6VzuEJnD3CEbZenZzLoQBeagMti4bUT
fh9lMkusIQAas5fv02fdnVnyi/1OLg5mQn25zJ0l/lJfc/bldhzavZEFKyqaOGbJw1KSfeXf9atk
2jpNXt7BrRtQ9HnT4ttkUHMqisdbBsHWXAe+JiOygubRiqfdor3s4vfJXP0C4g0jvoSxJK+LXVNu
SO3cByOWAcZcHevwMv6uQv83XmeFz1GFvVThi3Wd1YMMgekgzSIW+bpTadfrmkYXIGBerPV/jIfN
iHa6ipQaxWtJdCmCGaH0QgbfZHY4W1bqRAnQxr5GjKwLaNo5Fha1PKL70IjxkW7SwcZozzd9p0VU
D3sRqGwMMpmgrqpn3nHqevu7VbTWxewDjRcBxGu7tkDYoGLYnnocknXYrKSEx974wl/g42U6I3nX
Qjtr+iRFkXiv1t6mdMkc3BuYBJ7eAUsI9SUhDN+K7lu0NsDx8QYnWALGox9icmAlVmO0dhwHow29
I2dwz2M0FIbVRHjwvMmWPpSEagt/gDIdBQY8RmxHEThLS8ZEf72nvqHDRyoJr51T+vvG2baR1lMW
t2dHswO2xn1jRzgXRBN6aShGEnHj3BhhqtqANu+NoP7y8bk3NQF15JANMuA8uhioZds6w8mEb/9j
UGCPt4qCDnYgjjezNHArQZsLXFPh8j0wnfHax1r3oXZZXXGzJTGUz56gYnMSnYIBC6zV8SsiLXst
Fgy+mezSdnCtJURXxBCGOCGl93XBFkb/Sd1NjpjxjkO6KjekHLNHc4gZ+5I92Kx9jER6fKg7jMPA
YHJ1ULW+Zl4uGCVup8p+6T9rVVwETiaYbzaQ0bRm3e0s+/e+kkkEE9iSOH7xO9PiRjnMi/yVo7IO
2KH/ylHG/X25QnKM05nn4lVKpabMGUtXLA1pI+c40nvNo3mNHDzc7AQ8A9RaBIiuN7tokjP4B98q
DDgwe/syWsC5hR7tYYSrE7rhYs1XqwfwOsJjRvElRAD8mD8ji2PoqQC8jRSkJW0TqA0jKmjeduXp
xFfpddt5WwEKERTQ36nzfizbMYcyNAsrgDcki+2/EozimIzdjofN7hdPx9dr7cCAnHiPFzaPxQnW
oqtLA5n2H1K4hItAzo3zGrZmx3pootqlgI2EuK4pGcGOOwJbcV6xS0E1e/k14RIj2uBx9TAF6bwV
v/DuaAY+IkvdQZGA9eopkFkqwijqz96gBlXAFKXG+Iu8NclWv7rMF72k1xO3MGNSMrmhTJH5Q4yN
+HIlK3nevbxt011dkd5alR4Znyrq4MK0F+jDdNc8syd1D3ncqTlIiLVHRn7uNrPj3UmluOckXeaT
ebdfdvR28gK3zuql5/kTZtF7fLmwk28PccVyrJKxo73eK646rynVzTxp8GeFfvbPHfNuS4sVwSYV
8+yiV8MCsWZS8IM73ayXAZ/XOx0GMXeVIUum0ggOgETRw8wptKACBac9CAKXz/VUYlHQxKvdlf/E
SASHMmMKFqw+F+xAYUcdAioKZpDzfskd0M/fhh5ZIIpp24LrhbK9ibqdAmbW6EpVL/6gRnsz4ymj
YdbgD4QZUTRGmbsLf1p7Hjz5mfi3JrMvPLeOe/Sak+Tbh0xdYsa+BAWiu9BamxxXBSDpRNcSdvKC
hRYJf2ZMxSKMSJZ5twzzeQBxyz/W3ZlcZKtwZ39Jstv5H+CfAvzr5ILeQP9xYekyBlbILvzi6hU9
Kgez3cvmZkM0YfjqrnDqkwVPv0KMZ2pEm27BWeOZKuBtMJVGsQvUS89EXv/x5ESH9odLSDEh75GT
H3egq/jmv4eZ2oqNlrXR4nA6S12/0h2SSxgEbjDh50/D1MuMRe9QPNqyKsbi7WhR1vbZspBk0cYU
Lv+i9WcOCVU3U8lv2dHyQ3E28sfoJQT/yZRGIpTwF79s0g5BkcaoFmaNy7cp1Dn18ufRWK2OyYei
EVfK3kl5fa31M9uiZWwEt4NiaO6VCAGP1c7JQmmqGrNxNUdl01Dmu7OLdWGUGI58aZDg51vhGUOt
QwlcoCl3WLEA7dW2EeZsEmliCzzNYZn6myWxCv2UmRSDrMRluRA8K1gpxinXBRiG8fJJngucg/g9
oGd1LLQFnCxrb2Ez0Myr7VFn3gbcvFsdJtKC69u+25+f3UvrC2Sxhi/XZnrs/qMDSegELMfK1E7E
ja5asQnzPoEHjYMaGHew8qdC4uQBgLQwqh7cFl8qSSY8psO2vKzZAZVm3bwO3mRUxgqVGcEOKAwS
hOsXfKnFfD3a58vVGIP+jQLgyOCa7ra9S7Nxz4uQOGZPTAesqEO3xqCof2DyZR7Oc+I7lUiPYE8I
72Cs0ahDPJyKWMqQB/suDT3yKXBKoLuMLULZZdOPhUnb+xHv8qO+cWRU2sdaFh1Y9TXqfhCwzlfc
oRfNnRHuunqKCU8kGBu2N+qgV5Pu6hERbVadimhadwBQ2u/o6950or6qtABdPneI/v1cv5Cb95yV
0jgzpNifi/KJoXXx4cwkAl5O5ntmaNR/wImrXjDjRRKfUKIfTnMx4zJMvmcr4vFJEl0eb/Ifa2Im
F1vB9THZtWEIfNjctD4Sk77GK3DpgEv9Hn24/strY4zd96z+qSP3b1v6eH4OIn4MkjXMJAqc0dzx
kG2dmxkPlE0AZDzW9+G3fT9kv48uCRHtJ+agZIKZ59pCk+S2VEqUYLg98bEDg2DJLVM4uaRA1eDw
2CYGdBuB7tmMSicQSI7qVr/RTwshMAP7alHWbKpG15HaNxWR4xD7/DBN4njmeWz3VWWpsEhdx4PT
SxEYnB8ZoVtkPzqD6xTNQnonooaGOxGvtOh8IFBYm6UH3AI5rs24qtaJxEWb/0Fx1k3pTqxrdedy
yDQrwH+woPZpFb08mHcwX+37B11x6YXx1wRA+ue4bt+LdxoTjlLfaBzCgoyzek1ebDSRK9M8A/qI
xn6wCkBkZ0JpaIE7zthi+JOsKVCEFFZ3v4oBWA6OArNRZtPziH8Yx2SBg8BGyidOcLuxM3NLuiYE
mCySVpQeC9ybJMHU+XojOWQua3DOiSuW+3XW2wCKBVgR2EBCr97jlKatFlz3mJpv7iO1XBSDklZn
RH+x9mzJONlbhJqEb2OXFCAISGMpYNCnMBdVdMWIqOXCUaBrrMgZtZabTPBmuwItHEFhe/EmfU6T
VeP5VdnPZQb9sc0amsxx49rufaRrueGvekzMwTt4x72CAqAxckviQWnPkWdxYz2TnxaIlQ/br9ek
WpHRTAg9/ITUWdXf9v9Ee8GZQuSLYPP3d6fz+1oNvXIoDDHYlUrCliv1em1r0zpZp4fLelpkbCZo
jgOIc1JYqc6+Xk7UzFrjKWh0goHtmtzL/k25XsbljE6yysNVYsqRiajoJFzklyxjWA0YLcUtuB41
I2kVqui6n7irfqIcu/vH7jXIBWQmhAxPuWKWfONoU1GzM0OIcgPUKi1U/SfT/kYdINH7Fk7/AzFK
3xJmEmmOitboy/mdfpUwMeuqCnn8Zc0BCBEXORMMP4yb4tcs5Bk1rB0Rvl/Tg43FaXc8Otywrd3q
gOqlAD/LSMnjemobHUDKZIW7O/QGK/71W1IjoAPvcM9WswnXuuUpdbO9NALGqBMizZ2kXrMN4H9F
NdBumlwozZdrhBx4XlCU3B+PQaHZ7+gi/PQlik/kCJRst93W/qTfxauZ7HwTahEXKu2pAfCOeVZX
D6dJUw1kOXUZUZjwcTuz+SuN/13Gub/hseMmwP9ebci3QnLSr3hnuN/1TV9P3cOeizZTczcozMyX
vAzcTdaBZ9vySftaE7GuLNe3Sx8L800+WDjbNkjoNrHbl6bdUAuJ6cXcptijrnkmybqJK0wXzs3h
y0i+aZF/kV3S8FSp5/Ozfna8H2t7ht4gIwGi1PCB7mM84icCDCz3Qruz668m5dOzZxGgmc2YiRfP
dtbhnMvSO/MJq57A/ruT2zif9ibh3PG9o6IB4bhUj/p6ubXAzlP3pk5R4L9V0H/7EH9KTUe9OxyA
VHO0eeqFTWV6HU1lZbcihCocf7Vr/4D2nshejT4I2kagq8S5UEMrnbOdqqODZWCy62+57Jpn5qo6
QhK1ZkVf3xNkuDFN9l0NbWvgzO7sfsz7PLFBPNAq2z9g4n2SVIPp4/NJIKtdzpUMGBgMT8VDpe9o
tVoCynUzfvEVQien/uToje0w/si9S1SVWG9tKqYIZjHPDyUmtjadvQqmcIQQaji+pzjQssJu+mC1
+D3yNz7ekw4xt7fxbmYfJH73gEkVtFDnW1jrHGKSA03TXOaCGZdH8OsjwJ52bILfoE0gg6mbS2wN
Unkt3Ewlx3Qs/K9I8KtWNf9SGy8zAm9eTpFJ2Zx0bk/aexnAslonaEHTlM9VO7sRdU44HD5YABL6
iaFtXRnmnsay7BTdyd9RTDByhHmrwjbYAEvaMU0vFLti4DAdEhsaOr5Talc8iWNTECGUbQ6CXc6E
Ob7jb0yoEIUUVrzuoGAenyWj5ktR6yGOED2H/IbrzmlirlLL03Wu0qUpMjXadl0q+SZspYHLaqaY
hSxeCPwKpaEAPOHPY6hHvwz+TJFqBAR3zHoG0dTu81/XmIiQUhxR0M20Gc2HA63LSheDz7MkWqdl
O1JqFe+BxaFn4Gf6nixUGjJlM8K/0Y5JO50t+mSmPKG7/fZm9tntZyGNx19goSfsDfIHlstQ2T12
egNFzwjqyJUtmlMK2CsBuQs+hTRg+Ra6kPPWWjYcMwG6slL4Spgh33kZS0HNljK7/kGIcpOU7cYR
HWqbCPwJ9OJykIgszFfASXGeblKBMwPpmv8P4j61ZQ2kxR035uEI3IczV7E58+r71xE+Tj2qDfO0
OM6MBoDiNRfYCgnFjvxUmfVCkwm7hdjAdtiut4t1oKpbI39fYGvK4To98FYe1EAow2RMpaTXw988
BhCrwhUYo3WrABzw8FpajJs4Mo0WN1nuoyP97XTx+KzLrU3UrRTA8TAqvvwJ472Gj3Dx01AO/A52
ipwELCrx/tj5maehzhdJ3AkQ3zlulAAnPskrwis624qPBlZld+oAPzTiR4NBl4tPcNrFNzdUZUmX
VnDi5pO99UBbquEZHQPJSrSQX4QTOvUoWPvXCMMDoKtB/K7MmidLubEr4UtQR0xZhJ2L5K+QLeKv
oCQ55enRtaqL+6+YpysmmCnXrFdFoaHaJ8BLVQJounGccEzcZ1nho5Gcy7D8Dz6yFfTYbHrd92fX
O1qrgFftxh2//ZAvu1HhcNUcIbhialKofFEiDWh4/nt+0FXXqZRZGh06w5HeqwrD9N0WrFEzw/SF
GDO4G7AFSiJSpi2d/r7y5w4TTfC1eZmXYytEpfNwZgIiwoVk85yYF2c4yDWyeNBhUI3MEY8p9fRf
LPB3pz23Y6PF/sQOuVb0v+I+j+nMbuXMVvqL9oG+yhgI4KeWWYCJ/ba0up4k+Ni7bHozxDb5yCWT
Qvqu2a/CWKxExE4kvZfwtQ2jOr3QYFzf+K3GMzfzReqZmwYhWuF6VShXoSzW1XC+jFcMuZ3HN7kz
PTJi2hE2u0AW8gk9WIesisxneKgIgY3zbJXMsrwE6g0bfjBI81htXxc/SheBs1KjEZnu6tHGsIY0
aHJodunrmUdwN3eye301eV7qA57uFXj36My6ocAa04Hgmk2gKw1T2aLgbjv1IC5dYZOj8yUYBGah
98OOymVlDMyR8Cspp+SG4ytFI9ejEcjmFP4muP5PkZa2KGFKAHekCXViGn6OT4AiaEIJVRFOqEZW
whiyhfVhxC4y7QaZTQAMgb6hBHeIT6bFJ9MeHTdEl35WrxYWifwNYu2vSvRYLiD8HOWNgYSAIAPz
kiwmNsJCbVvgyiJ85jSFGFsqe+icrg/6kSuEaHgw6fjWSUr3B1Svbj3IW8TJYzsODxYSAHh0yESP
MJ6y7tAD9rdVky4VKYuWhzDyDy8/keOWeu0ip0sR80yAv3T6odTvS6G91ncGHMtoc9PYCqtwBG3Q
CIRMC9AP5QtOLNDN97bevN+xGvtDbEZGlMzlwgi9zgaW3sjEis5GzZIizF9a13zFukzCafmtZafg
VLLlx9ftjL3RomyRiFV7qP8rb/Tq9emwbKCG5iOIkHNBO9ZVQ+BIsZ03TwyUqg8rpKvyutYdc10G
49E5dP6Q+XxUv2trRmOMv1kK1aywgzBt3MUB5R0Q071pEevW9n0ogKqCnKvbuTDRRluaYx4A16in
/8hRdMp9CU04Lk4/ynYXoB18TSqDFwxNwoqpvPBFHVrtqkNmfaPaq9Xj+SSPrRdrNCXyPjGF8AhU
cUZFxHqf7edMrG3f682Ay/vOUY/3W1dCVWHP3evaezTmyUnwV/MLUmwKziapfnYD5SwAnRt39Y7k
RIWqaB2X8FMhM1bjAwTs02Q/3AyHrp29mmmZn5j/YZ72AmoVqS5hkPcN9CI9+LOSny6V0UciWEQE
fxqE7abCdmOEjcF0Mc7/DimgeseNejLUd/bEL/be0zDjCMmtlLf46GPgW4jb/fyBwva82PdmKf99
PXYfQ4FRJmSeu4qRX638rkTLDrFA1Oh29EF5TEc+VS4PWvigcIhjet1OOHr0DflxF4x7LU+Yueaz
SHiCyoXvaST8YpzOa+31d73UxCVAh4O8mPgVLhl7MXLd259BMX1T1wgRVkYRH7xESNcB6Bm6jVU2
yRSW3lOEzJ76l98y67qwUNGw7OLzzVaicM+7vEu0UCuq5FFiEQu+5tyrRzFSMVBnNScQ7aPiU9FI
eNZBK0evEQp29EXAXJ7t8SaJXaIIdi6re6XseAotQ4pDWfh1gPMbt3oIWXUbd4TsiUFxctfQpH0b
NZPrrWoPjGPSm/yds3MR7qUjOH9YXSy9MP8gbsF6Tolzyn8+O3Lb0MGbr7KN6ZD7kEbrTOqezCoq
TYgE6VNwI0DEaxdhFOm0kahuFpR1F0v9AFFVH1CCnBnu+eBfAG/a5qpb2DJRSWGc2VgjjKv9w1f7
thw8xV0xtsyZEdrhgGWbO2r3RNwnqYcxJAG2BhcCAwhTNFQ7D29GPY77FkXNp2LZZcHZ9olb5aGE
9R4xaTDNsHggeDBPTjaI17rcd8scv1Em8VrXeg33F5DcnCsYRp24qfc4wQQijKyJXHZYnXI5HXwJ
OyJKPowzAvMXxUTbYEATz5iMDHOwuhKiD5aiXrvI/Gcrr47XWBJS6+JmeDlC0iibUG2Y5vKdqr+X
SKB3wg3Z1xoZEMAZphoQULQr+7Vstb6IAr95mYTnm5JLp4o/EGrqjZWQox5DSiP11k/uVZPNRgiE
ev33D2ZNG10IHu1gcbeIHE9HH9fwzI5cwTgI2+cxN4SknArzqAV46CZu8Ol5b/DHTcAzBsfY+Uvr
eDgQjLk93w9Hz6OyJObOc2ukjTjw/Y3RrF/N2taClHlvcVX/dIOkUTebJx1z3X/elsaxQHrYpOkr
D0q7FPszgzrydtGGlCYYwW3VKPuX1n03TYmr+89HiA44vj4yDbZw2tCUAefiUoGFZjtyBPS5fstS
ayHYCidO2D60se3Lz5qw16y3cxf9uwLfWhUyb9iV5FTY8ovEpMQvelcgXP9Qz1ryYYFf19Ub+Aql
RYrMnZwqUFvfuRCC8vN/ZcFwBzeCTF2H63S8VJsHcJvm0wfJWbdtRgI4kh8lWwmV7FbEEZMF6xdn
jbjTRb+uA1feZFPO/Lptd6qfcWJQNNMm0UazvzIx4BSI1ZAHAwy48IX4TKLa+YPlOCLfYq8V1mLr
CdnTVxVWBH6FKP91u8hj9c/ILrD+848t3i67qQlkduPjjsL8wRyDslXO4feze0TvLpTbCdX6/1Qw
rz+Ctb4lqDBXPbBRyHk41Gk89kz0o3lPkzwBMQ9ZifrpjIO0JtSPFpOAjiDv5nOAlCPE2hRrRQvW
owmAKjKTcSjA/XkssMrF+SIFUU6KGQ5s3kjwyJ0HWZ795oZuIuo6Tp38RCCQzkYZ4I8mUYanqbDd
uzoUWUH7oLzl4EWFVWEV0ZAaSHJP1arvPKaPZQPDBf/2RLloJwiKybu+n6evsVZYSuktsCxxGvK4
rKvWiGEusXHOngqn/+LUwT1J4FUT8ZuDjNeYcHvTpxqIE7kZpb6dpZ/W9xB5k8aGArykjzuTGBqA
cpq+Z6vDoMh/+6Cz6hasXP8/ICwmv4ZNKtGZu+idIgAAJ4BuQuBIkodHsmzr3cisZL3QQc3hSsml
JXS7UVREvVeBO5hPx2hcl6ZpOZJmPMX+UWRL4+k6X6UFQv0dHtnXD1cuFPYJJw+teK5siVz8vA9F
/24qKmEWAuC1tOeZYIis0EB7cfgTmbmb5IlblMEPTn4xvvh1p+0OymcRK56WGazK0zYkT581F4c6
ppcuw6ClQt3ILEpRrSpwFVVRrR7PIh/8Rri3FmLXU9JTibC0aPa3RNcHybHIZmPMUvXFF2cJn+lC
n42hYmqEM3kg7MdBS65nbv3s0vSkQbL5CEu0HXjQGvfLn5yPB5/nr0Na5DB8zaeaTyG2YSzXwhlH
g1zYdfmQGv8ya3lyfAvFadc0AVxfSyjto4cpIBmj6YjfBB5awTmuUfk49ZB771E3jPGtKP4e/Mdg
ak9CWQvSXYffUNvsxt82UjKlF4m/VdTAXZikNhEPEbB6Mf7V2+ng4aEum6KdgUgl6wHNM+tnTpRZ
Qstw3DiCR6QeCeR02bh/s7nsS0LdwjOqmQU5PL4XxFKbr9eK0KCsT8G+X47iluZPQzGHxJqtA/z7
pR9E+FlprTtPuW+Zdx0bbIhMDkXpdtz82uXh1kQMbqE5rfPQQGArnqIEpZ3FDJbp6Z5g9KjiJa0F
UVquIHR6+Wm3nAxGokDsezJRTnNPl3PcWlic0XTj0Z2r5aaP3CBu0SJXoZ5RuiRUTTzsGylYXopj
5PgucyqpWCXbqQfOxGKItWZ5WlXihdONlghJooIEwbBE1sugB50mTUMFB3BNi3Glx6DYRx4yT2hl
hxQ7x7Aciplzx6Hv10O6wWtXmhYOg5sm6AEAUa6dA3r1akvTAV4puyRiz65gsv7GQOIdPaLysHVf
sx3orgeWVpm4Q8nPw74QdhpP2QG4WRwoljnrCrsm12X3j5biadzuvc0bV4vmzz1pUc0s4WY31Gkx
TFmomqQBcyqsPcHiE5zYg9aw2ahj13l3Ky8i0GbmqpqGdtQgtZ3n2drgqbXXZ3o+ne0CDHfUIUgv
fpIi8vmHwTwqJTYX+GphPsgBVWmzHCqtkXhR0YEydj+H1pWTD8wB6ZmElRBbQkUj84D2ywtt0XhE
8wuZdcwEjyrUxOk7ewtB0URD5NbQRpUGZISIvuF+mBYMHis/SYXNtj0KRi0D/bHo731LimC63v/2
m7ZkJmTExCvK4vZnGmJSjyRJXFV29VywUy12L+HuCjma/akMJ1onOnmFIxT9LCLOSuGk518gcb+R
3llohiuEcztf+iCSkEO+EHp6sN6H+CkGV/SKQpaUzRUqV5owPiJmLfmQU98buBv0SpOjGYXxfWX7
pR5jX9bEvQp2t5pMaAmq3hYfJVGVH/4QzIiCKCbnFij7Tlp47DNkpo7peZSTWMezkT/HYgqEUQC7
Si1/EYkPayMdiyhg9D50RwOkcb3o1R92TkBSyD8vUVVzzWaylBh+iVHDzCVxmTYt5yG9uA7MiRfU
dYoAnShUiFLnNeRQsjxyX13FBqktmdh6EVenXPVgXYfSeEJStbudBw7eodxIYiH6A7gtO7uqJ4Wm
nPV2hkFx531Q1r7HzvrZWg/Ozec53u76WXTDrGbYmrjYVYxAOlj4tThvLJciWXBh0JxCUizZuUH7
lkbDqSu9yfWtyZ4OTnJMTsVLEAn3uj5ua1i9UvyOGuc216uMSKftuXWhAUq21a06nfUXVDHiEJse
vQxtDTrMlFPZADkaQl1uKnDgelHwJhTNjXu5vCzTqfEDBM3SdIxWoRiAAFmMN4T6dK5vL/moZE9p
fYzZN+DEHvxPWpju1GrBhXCkjW1Iz860OC09ybaVBNWoRS7TmkTLKOxddbyvJmRVo2IlGxKjg7Nz
rixv89jU/v6lB+6vPVXmSNWF86om5Ltpq9bnkhj33fAE8QMn05RJHrt/qPzN7fiJyqwLu2TfxM2w
NkcUOn3xgD8Qk6r9KIWUpmcDvionU4B++sSCNzq+I80XByR7ghngG6FT8RveDRDKKUWyZDNFShuE
IoxRrlGFvzyaUIzJ/hFlB0Rtz2WiPfUxFMmIdNQSOYl+R1iQRGvlFVTTx2onjV7BehoKHTSZi6K/
xEHdzsULlHWg0rxckFg7LOkZvnoEgt+uB3FNFbAvfEKsKkhBETzHerCF4m0fzY1EMkbz0p8Hlg3t
l3WtUsyBlLrZfg+cwjkjaKN7EMKEh5Pd4OPUGAhd5LdVjSWZ9lcHz1nfSKlc1Z4HHCG7zdteu0YZ
0kSlPX+q6WfbBQRphitp2ywitsXGastD3s6i1hBrzZ4/RlI7YKxUfpd4qOTrVne7sume3TlSQn8+
zUorNtfDcce5mAXO/5bGRiswhq/5zBepIS2XkDbayqcMAzEG9FnXQYGSHkvUAfXvqFVmqFv40Fg7
fCM4Y8CKy027wd4y8oZPQEhPpbrw2wzUT/nHwq3WflLX9ovXbqZU3DnzeL4yMzX7nR36WOtk5zTl
/XkcHlYDBqyHmTQCOrhahCekYDeoI8tpAeqJ34S9V1PL7UREvM2UEs2VaKm04900/x+HVbym15R1
rfRNQ3olQ46RPZEgdbQYP8iDtVoVgASoITdV4+TvbADHqzTXPwduTTSCslbXY4GxyDzyuGLBw2KY
lEFMgtwerilg9A55my7lQiuwzhVl9MWLdTAAqHheMKumwgVUN1ds0e6A1F96F3YKEcxxakrMIVMm
ORGFJpjVlqBWzEOKC+wO6m10vvel81t57LAwWikgp6/JspCQto7lOJ2Pb6xpMX0DKOUvI/OUTPq4
oPVfcfP9pbAJqQgxvThmUcT9lV6yAIkWyBoIvZdBhYXkOp8GJFInYAnwVz5edMDuUToUwofv0ToX
fiiecjLwVPoi1BzQ5sAcf4ADUzLNLtWUckTo2OrlI5gVW7/3RZQ/JuF1Zut3MjkwsWhsqYngXJ5l
Z3FeF9pv3K6oAhAscwmMarV9DRRF0ybMOeDbRtmKx0LQpIQAYESwQlcWh+5J0MWreOEEdlB9+P4O
ztwypaHKU3fqw6gA3kXE2DtmjCbNRM54cXEGuahq4dzQJaV5pvXmHfH29MfCU0gBQiHSxPNYMkeN
Cex38pgUXZJgutvcH4kv6flytM66F1YQybE+mpX2chMfGo/Nq3SfMVtMIPMZToR4Blr38B2zLXpH
sokdUzq6/h4pfAVNeqW9gymB2/XTMIrVUcM7hQglPbX7oZHqheC2BV9ayuYm9Y17RuvFve/y3CgG
A82ui88M7z2xmBF+GvWwcQ7oPIC2x4ibtwmTxO4mIWdN3oXRog8YbD0nFfAc3vokzHJYBHoR/BD2
xb8eIjztT6qt4L5ZWb19hAh1RksAC3xUgfxw+t+uVQ8ZXgEJToWIqEeORdnstZzII9ILt4N3vdc1
5aLSbtH5MtG6lelWnJNcwQ0bm3tQDLWfkCWxMzLp4K03V45JVKjePEG+7N8aHPbbBsmT/KZUAC3C
ZTCWijZsAc1orm8QfUaMYzjqknMYuem45xp37lbjBsWAEM8Udqj5UdrPKzx2NcO/1rN7OfImJ3x4
7lHwn1ZmpzQ5d49wbGorKYm3xL5PQbXE6zlT0tWsT79ZSHYOQBKvSHYSUPsv0eum+WMXzU9YDBWf
xDaUgcqq88wLEKrQMzCOlq0v/3Sc7Chfzs3vRDWxZr0xhFx4TZB+NmcWFL046zL3c7eiMIf8snDc
KhQ7cwg/vyPIxqCFMjARQOK6XYHvdeP1K8QINHdP1krT39+EOLA107CNbWDg9PJfWwdqDAQ1CnQq
38qWv2Oy0axNn1aeKLuv+fi05paKAFJD3dRuh1tsbBScx92sR9WcSzhonr5gRDDOvuCNte43bpGM
9PGUdLYUSCGX1QHuQMbWwKSJ6Bz2UKFMl9Rv0jdEPwvPx2T+BsoqQXsOPEtWMMMnrIzZmUpiR0L0
k7h7FV2U/jiDiOpIwCS4BzWaGvsFaVYflW1Tv/MMN3vi3RcLQzaz72z7VCKKQpWGSrwBYyZxZ/dV
dS+i9stRzwAoHM+FzOl/WLfFslP1CE19ncpm43HODLKxmxTLMeOFegNYDDSfh0kggyWDAub/fURp
CEorffbkhWKMMN5wcztksaPGwJLpICvf6PlUmyM7TlGyxClYvhU+c1AZJ3UTYKg5B3127xq4khqg
KuIDyjAs+pwTdO087gA4Nfl5rMdz+WJwwyTN2A5yhtbwfGdZF58b+9gpngnIOTyTUYMMrXYAdQ2K
twhG8fiXBHq2zz0b/uEGXjqWjWWZd5h7OwwW/i/fhtGxeMiO0ZaLUEADMwFNRh08ShCJcwBQ28qk
7wp6TPFnhh+xW0n1HRuT3uazMtge3aySVNjgQEe2pB0GKu3DTgSbXXM+et9qxuHisrfqNT/lpFex
fzzXfa/TCYiJfk+uYNa5LfmB3HM0s9Y9JX2OSZ/FkfGx7F+sUQS8e1K29t4QolQeSeBkLquVMyzb
0Nr4hwHGb4fy5pr24XcP5EROGRUwwJhIzbsn7DA2vp/eYbu5F6+VUKUHv1RgdgQcOIjPBP3cZkKZ
XlYriBKf1P8JpfoXTS0QU8uaW/rcLlxlA7kBtjVSiuLeRtHZa6jM9wGbi0vBLPL9iV7rWWHvYrlR
xl4eGIjNFsUPL4c5gXp3bEJfYydBTyBEO1wX2BaEK9pZAtQy4C/+HJB/1fwzb0hUG46gQzGsCPmr
sDG80MjiokYU9+Zf3jav7WQuVKLgndbJcL0Weh1KpZLBA/jiH1Oh65qLTHlm8cLC9PkMcOOkcNMq
1uyx8j1bPZVtPBVeOrAfaFtZtgITjBBgOr/x3vB4bL05mueqXByB/HTqNShTPGogoSXQMFt42q7G
sjrXWbN06cvme5MHI86s2QOd0Gqbqg7Ir5fBsta4W05MG/ahn80gWhTspdM3mTFOvCF7f8gOLe2Z
P3wfAMX8RI5XZhbi9A0jUZhJmjhi9RyqGzKczadGNUn385ly5jnBl4/ESD36GTVW3zMB4Raowk1t
xRjFyTfeFyt5ZdkJxAmnzSWfmlXzl2V2rhQ3vzOYQV3Lj0/6yUkzs89Zygswy4WEAd+HqRE209gv
22MF36PlFUBM+2IgZKO5MQikj4Xo2SFYdzYJNgcsjKAtWjxD4t+i7JmKneYVrBsxL1Xx7jvuJz6E
fuYqI2OL2csxFYhiiaCnnbtYzdb1yLaeTDZwn6AG4z/XIHqImWEaYwi7W5rP730kPr5mOOjQwsYI
qtq8xVeABYPw2sWAPD/fuKWcu7v/1JcEbK+35mk5cso5DE9uvDZjn+korm9RNFWdeEChA/4G5V1i
AJLNFp4wS1msZqFINF4vsVWNOh/bn7z6UCCyfu8bae0S38QJmVKNydygcDW5z/plDJNP1Gihx8rW
aLj7RYLN+GrY/vxiwZyDCE2Nnnl/M/PKAFCnZUvA1kJQIbnROczUXlVw/5KSjrFCbbWbiMpOTBj0
7qX130tLEwlpk6KUkt0SST/k6RkTBUl62f5UbyATjtfDeB3XCXQZABPL+pnTMXoNL4ru/PLtt+3u
OtC0RytnkEUCVtUYvvNDY/LDx1+2lyB4wilx+APCwksO7tL9LuONXnZfET9QrGRwSzB2YlnIT9Nl
f5hv6SacI/5/FDZWAUx0MbwJiWTYSarYMpvFI7lquN/UDUD0BcDchkmzPFpvNWsegOqNMdAaNZCd
UXeA60gWiUr5SFy5cSSPFNNTmm3KtVDvLpn44y11fMH58Gzb+cq+2dOZHlL/cGu787UXX10h8acJ
j821jOXScCWFgpbNuCXPmhIZmHwU56BOIlx1o5JVMdeiwlvONuijd1T4meOH/ZYy8AjyKeYJ+n/a
dVjo9LjV6OFmOWbDbPgWUpVMb/iP3hy/UW7ZGu2JKVJKxVIOyOYXysBK6BuzJs0DCgp1/55xz5Un
+8RQSYWpiaUBNAN3qHvScfxS/J1qNEd9WowGvgdnOZFVeuKDynkijwjl/nuHxJm3lNwPNelj+xSx
qMYtg5Hfsee5XZHoNNTmS8qyxb1IwhTgZxplFGSvsLe4BNjYEpOdjGyHZ/VoBgH/uXkR2SkiMPF0
KkDOD0vROb+MCOUMSTVYl1eIEy9efocMsxmP7fiKN7oNgPoAS8HU2PnSnDcqNzAfqcPWJiaahlSV
RZ4TpCpOXuyBsB2gbTS10Z94Mv9xafJOr+qVy0cEXhfWF6d241CVL1mcAxqRlgpq32BSdkg9wkHM
7GzT9meS5qcn8WNYjiwnf5BQ0EVkAfsNrcO3NBAwPF1mRlFvruYijRkGJU4XWNwBNJhqNke0APaQ
ElgKscWF/MXtGPyydpf5HcQwdQNrA2y0ggOx5hBXXBPFj7aUaws17WNXSBiwKkk1/XDCgDtryMzg
m9pBFmvw02fA6LjY1mA/LbAtHxuxew6RoEDwSMSZEjq5+84hNaw2YYFe9yKDxFv6vc4lUCoaaaxt
tDODjiozQOSpfDe5bGd5piKeAT8gD+pQ9+S9yQj3K9Vq9DomdO4j/ilO2lUB+MeYUnn6NoRURnsa
OUqhiQ6LYlUBknuXWypjrMQu2R8Dr3PmLxAVFlJL4qqmhUGEsLlBFS0eseGMa46QpayC57oMqlBp
zeBX80J1fCn4xzIlKElRMuFPRqsCEOm61KC1+5r38uYLX8CD+irr0lPTPKCu1SMgB5W6mfTIOUf6
GVWAc4J4ikCG8NBW4iKqy6gHkJao9vrjPfBvXzMdftVwQGDvkl/+mr3IISVsd9+dFG0I3XMlPJcf
Bb6w04vNzf27rgdHzT646HO8aTiA6DmQq4DmL0NSfk7UbnGbVBONoj6nOdthvnBwQ5MtzxEau+4W
aF1XPWe84woOQQsIAX9e+4r2dtGX7WmTe/0wNelHeLN+Mhq8C19I+ySLw0UStrIdbBQbw6KK022P
Bd8AFQBEFq1zourwbNrXyofH42y+fxvaMrFMsS4LNtTEeDuGs6xHCl2Y0Gs7DftGK7hVRdkOaLiu
pFZ3UhnMErD2/ju/zBncW7XDmMZpW8rjewJS1MUlI+A2Fetqdw0h+kFAP3iTtj4vl2TGxBX+hobF
mt5MlI3bRz3diS163ZJU+ju5iUpXxyjZMgAbLWiCEfW7QbWCCfxnYpiBI6oR3VFfJxSBqq6Dci6X
BtFnoD0qWaty0Vi99rMawhKufpLqwl2I3HgIM4hn0zfumOf0tyyw/v+phRXi301509fAUfoOXb72
+TzMF9+oeD/z7mA/6nt6aJ2dqo/Yl/Aku+rOrk9bFlTrGi9C9ULTutqmSi5FZ4T60gmiaY0QvTkA
veGpdT9b2aBYvmcFdqm9YaQsfgVkzGkWGWE6mV3lIpVrL9fkglCTVHfbnOMXuxhyNElmNdJV+xhn
YUDL7HG8tPSts4Gtz4hC1fIQtde0NF15hJlGexYFJ9KKRUGI7SD+iMRoLkKaoYqO0Y6UPQRP+7BL
vE0sR7dbfQuLnCmyyENp0rNvTy8aQjVxBl6oLQoW7yZPgWY2xJjQAHzuUaUwQ88b5C556wg9aHtS
0ggA99KnL7hx0fheTS/70F+769w0O8Qy3tSYXvH6C1hWBbw/mS1hO4JKfgrrV68z9t3zfLyKDEPG
x37vH5Ea9YJWWD0GLZRVDQKXMjcxG9Vz0xfTEstj4hIRA/0UaTlrnEx30HFtMktRmKx73XC13t53
Ol31yUkdfHuGr16y5K6SsVJ9sUQyuHYFAU4QmNaKfZkpYkNncSvIQBYyRlZl/s1J8He4fWQ9ZBph
FhN9AVtMw2AljpHI1+vv1GcM4fW0lBVe5DF4FtIpXi7gLcN31SScb/6joRsLglnVKPIsQiSGf0u1
dIepXjBxV7b2d88wbohGGxL8XDrUgcw7KFbwQqGNXgTnt1XQraQD77momOfKZLEcqW2V/65O0Ts5
bpxUwYRkW+7kNbqHqDC1RezA7jS1FjGQtSmUtHldvdUXFicc0dcw2hdADDiqbULmv6QAIbWWS4lD
lkO3CT5IoWYMCPvFvgj5yJMYexinalDSoxObH45lUvhbBYsFAfcD/eTKK5mjZTWbL29aIOc6yurW
VaYxndGRfODfcMlWHxYS/dNQhr7Jqepvp5EqWQ1jccdCDqUfhF9c2q3O1yqAGbR+oDYQx6FDQKHf
6Rzm7bn+I9Kf0VuVnh+3o2H191t3Y3k8ZDTNIrAndY93ODQdkRgnkaEYNPkJkp1g3Jx3l/YuPL8/
DHZrqho3nwYOEOugzV8MpO/rQgaYgN1rmFBnMBnKcnfnVymkW+8d0yqeudBqKm0rGoW398/gBmEJ
11SDiwy6EY4hUokjEKglJ75d8wgrpKTOUtEUUuwkIvvQKNm79h+xrPdK+g5P0KdY8PXoKx6T3ewu
55Zdm+aR7hSLoiI80oBRVMTJogXI3WBmeDeuFEZ956KEmqUqfusfwg6Nsgs3tTteIMbJgvLTpwBO
LC58vQ2BaLOE4G2XLfbn7EVDcNfphP5e9TjmwTATQduulduWJtbb2IRUicg9xtqo5f7cRbfQxzE2
Ozc6M2g5WMc5FuSIuKZWf1S/9aKtRKt2B/SZyqMAZmCLV29Wzn0Y9iQ+SP5b33TgRFyYg431YIJ7
jTnNfKF5tHOj0nx+k7pQW1OElsISiqOGQdEUAZnLa+6s/86B1EsptoyEqxc9lREYeBWwpg45r5jO
WVWM7vI05ZI9Z/9WOF8l+OwKmczX/Pex82zd/M7UHA9b8Vis4vXLhc3xZRvi6tlPbKwECQT4AL0Z
FIUrN1MHwOMwXzMa1gqum0PCNaSmas4ZkJ59MMdfgYB9MEzcHDKmQNd/m4dQBc4uRbGyC7HF0ojj
a7GgUq4Loozd/RJLUu3mvsOelHjpZDMtbrtnQ76QoaeAYW0HXXeexDSIjRfZWdyCyTD1c6yPrm7X
4239bF8BNxS94A8BsbvmU6hfkx2hlZgREY1DbhRwv8a6V+xAdILzFFrtET3iirfP1NjVGT8LdBpP
U0B8P/dkXe5IxSwP/NNPhptMSw5C+f4zhoQdk1Jhy9AxoKECACmV4MatzPlfNEMT67zwD3oodQyZ
uSbtmsVN95r6LolrXs8TKQT5pktQhUY2PHfHOZEauew8BekoC168UK/cYstIDWOoqe5ym1bX8uVa
ApzL/zvt0vR93alDyHO0kWP5UMeMG792ej1eNg5epTiJ0Ydh/hq28s8Ktmz0smXhGOdPLx7u0Tnf
Xj1+FqO7c35oQJRGEwL7FeqYUS5kNIP5tuL32YiP22ePktrMAgpY8rP5MW7NmppS0GgTbDNloKll
6ltKHTt5D/yRuDLR1wty8gWI1Gkv0Ed8amWjdBS5ILGpSa86ZVufa5Ocr5qgOS2cOrhFGHrJRkvS
c4YMxIwsOE/9ipZBM2QtHFyLPznlI+SPSz2uCN+G57BYcl7uoHpScU6TrR5oPbuVGHhzHGsGfrmm
vu67NAwM+Ao0BwDoppbSuDd9XFVnjbWR+W2BpHdH/7MjLyeuS+kYMILEVsiClSMg56VgDFYYj3B2
p+F+RGQUbLtYR8YtMGTd7wsEYiUNSXZvu2StSxzvaduVjnPfrJcgObRcPVDXig4YMvGV2fU9vbed
Jb+hz402nDKbxG6ZsvBbx2dUxvu8Yis1faqA6RKcJGCrkINDMlCuJOE+ew35Oc4mCDXY3/aIaVS1
Ror+owYM3d1NWOBoinmTZ6fntS9K1ygb/Z63qPDXH/AYdR/BSWbcbS034zOP81vdER4EkF/c4Yew
6CidE4yFL2Oxt5R3gQVSQA9nxuZmkJEg0W+mwz3Uh1Nejky9+rp/ZhvgYvDs4Yy+pB6uSMbvh3js
CMlQihW3Zba/UFbcf2LtP5GGzAbPO+aN39s9tS04Qu3X46miZjDsXVOTjtAnMTs47tioBDb3FDQd
lPU2xxur/vpnutTecrD837xt9OagjsIrACfCedsaEYZabFrc3BC3KfLExOp3Num/MTjIL/ocqEHz
DO2iQ3W5kta1R6f1JK+0HefbA9mLCo8a8RlKa3AhwEKtL0cFHe6QjG8EcwdwqU7UXh+4oY3m0YrK
RRgMQXFc2pudNb0wmJ31RNgMHCcEyV2GESRi+dRBEcFhyARf8pcn5p083DiYy0EYi+YWQV8rI/gf
48EHNpvmfuN7wbjXfiWzatIrzY+2DXcUmBKof6NMM78DqtCD7qs0GbpbJFayPPZRSxsaA8JaZ3n7
D/mdwzKdzN5tIZ4YDKH1mPQOPE3x+19iV+WjBTqZUV96uGuIbvO1LhWzDpwAaHDJA4QA5DITDm9F
ioCGmQRcRRiEUIy/rflPg9mPXSOvVdkuHXy1SvCoqVYkX4TwF4/VZQitjwDnblPY55Q7Gs0qE4l4
qZo3xb0iSHMgtbXvBCiuZFpo3TdNP5nyvEZf6fDQ0b5zsqaOJvsNUQ5oEt32AuekkQQnR1IsKEP2
SDvfZPgBwQyLk7WIZUkXnxCLaNozczT7/YhDpRHSWq88+M4o5d3ATIOLcwcBkre8aTgYd5bxJK3F
he3QxaeuY0uhDI7QPazBNY6Lq2c/qsD8cVQD3PbVsIrF8NeLjiSr+H9+3ufiN+3eo82ClzLH6nv6
IAtRuR0lxVvfYCwTgshlhyjQ61o8pkwmezxjjU1KZccQN6DvqX/z6zBwD8+1D8Auz1AmuWzxym+7
UFP2mAmnWvU1Q6ZUKCZvFbLk7c+u5ALWHJeT3gQKo+QdnqsaCZeS8zltHqeZXS1SG9CvbOUk4Uth
Yu7b7Dpq/KYUyNK2NzjYCj3R1fkxGK1DfYvXuFM9jiCNL6htwrCB82sd1qOV2Tc3Sw1kwy2gTY/J
dnSSHgdwKVFZz0tCI1+8K4niuC/aJylPZacFW9Ga1SsdD+XzOUw8Tfa2+XOAxAAPrzbMaNqD9rDx
H8TLwcUvor61zPSAzxkXFj5Qjq9imQePh68WF/eB0rrUQujQyuHaXPEdjg8fA+GVWTLUgsPbKRho
oWJUhicTiqudkMJlWg/E19q4R5m50enioYEPYfb3kmUHZCZH7SEdGdkocUlKExwsbRUEf9odAWzy
CpMvU5h8/20CAT20Z2esPe58Mb8LfXOKoa6WJzmrU+R3BhmlqlGtj/cTAMPKaa8M2wXJ1h4gkQ/G
JCqhveN31drsrUIEqApEX0YN3v8hC5WJE4qPdgN86Z4D1wYzR7CvaKxbQRGq7ze1Tgjz/a+v2HhK
K6UiijTHgF5hnnz2YdeD2/26M2ZioNy1SPSwOYGEMFdO1Qzo7sD0Cp5sNRQkO0WgfDO9ECIPjvRj
bbSIiuPU7N3ZIkCx5GQrqBjwY/W4+MIA+G9TS0JjSjtatH7yWtWInmOQXZbFXbSXvrL7oLOBpApY
12itRTshIPtGH+fv1/bK93mhise8HDwVxsHZ+XbweSQ1DEvP7PEIN9Iv7JZ5rVTAUO8GEgADKYO+
VGi5jakeOln18VqZ9g+vxGzbo+gfbaXcoHHbzPi/cljV/kHaModVVCuxNLaVWq0udA+35sFZVk40
mwEBNFKzW57rX2RqDmfAMW/D5QNYy0qs8YQoTGb11b8p3m13lg35gxaPWKUpFmDXrmjTAef07ZP5
1HlchdgH+9q0erhujmd/3ndwBmJpSCro7Vxt9pkTtF0+68V3KSYzfbjMz6gXFNXgU+Xx2vzDtiQF
7LMfCC0G1OlH3NpQJ4d0Zkw62vp+E4S1uUNEzZX9od+oRa8bS7qNbHbm3LfiuUtzJS/KETJ/maQ9
Mva/kOdYmWz758jhMGmxAtFE/qD3njzkLcmWmZGBoUO+4mPVPsn/N9oVr9P+smHJNZtz3ZbcO8O7
8TOUA9VtRDdN0TMskoBKVcf9Gmnn9c0emZ9sp3jemPcNaDNDr76oRs8rU4xLCLekeQHthyai1d5/
sXwVFXTxZmO6+3JplACSDPr9TZFEptGrTq0fyFZ9OKih/Je3TDDf84gg4obXdh/p+V9fqcJ3R2QR
DuMrm2y6VvCYFlcENL9F6GPZ4yFPBAyhDVvKbVK0Ws1BQB8guRoi12UvDHf5JdMMQDrcFEp+Pixl
TE6odM7X5BfA1PGU5WbbirPp3wg4OM01WbUZsLrZCrmkD8qcwL0ipP68PUdAd/1Q0s14Hf8BdYwo
nhYF5FOkWh8lKop4B0JlyoMOWmXZrCLje0vZk3Jtfn3eqKASTgvQkUs6TlcYzlUH8eepeARfR190
02BxZrBT4c9qUdtoTeryNT2VmVA2eQbczqbDJ4JlCEGrr5LEapXmxktHn0I1Cd+tkkKZ7bUON462
aX1E2CDpTDByt7eD99g7EH9dtO9/n4OeaBAnUTCaZW6PaxLQD8ruPv1t/ntaOS4bgnU5DpCsfCgn
LSJ2hyDJ7921YLM59Nio+XnFiZI1FD9mxbxDYFDGicS2vfr7gpqfMhhQZqcMGk33nRV/x2jwQ8DP
JLhfAjNLx+0p/dmV3NF+VKpc0SgkGoSVnxhXZYr+7TCzPGdfWrESMtr2hoEP17V4Gj7h6lumaa+m
EUQqw359o3olKBG5ZYLQBeKu8AZ8DUp8+xqJTkd2EZVYOq0zU2541n/2B2DI+RQoZpIoVz19sHM3
3TIUlSEVVtDVV131eGvM47qrH3xJXTMdYEdDsKmPGAvYgamlFYq2ANnzpW0d2UpcuKl0HsRMWRIe
j+Lej35J7yUEbg3I8bRVpM+dFM8J8GHB4iqVKD1oPemzkhweQ7NJz8x2dkZPIeQOd2YseeQauXpF
hDDcJUQJ24Rdzj4vZGP+kCKgI9ln8ga3BVZrYxbLz1uJeloz4C/FzsAroz+degmntlO5azOdy3t7
RL++TAxIaidTmMqPAbFPvCfJhpHVqMq5c5tM6UyAV6X+iNBIV4sHNe4NVr3hOnmr53WNHDl5FfWN
j+nSnzCdHkH4YIIyxRylqUyLGCZsFoRnXBfeE0lMF6cfMqvfEb9H+eUop2Qp5HZexGBJHKjmc/lZ
y3PJQYOeJ7MWbkwz1UQWlw6qOP+iNtE4bQXIPQEMv9W6qqbQGz/tc/IaioiqTAmZbwNccpPpYIb1
rtjN4qcZn40bOKDoCsswGweFs43VwoJavG5SbayvmB2ed5jNslo/2GGoqDNClN2WAEHCCpJ1Xyq2
jW9/DFysn3nn18E61jHUBEF0VRqyUQADeJufb7X3jaJUASjvnctRF/W5hTvBFXlv7do14eik2u4W
KytkRNNSCU5tmbUMA1donB5DP5EdJblO8jb72p/yZm+VOvpQFz5tysTNWYs9QG/ZO0n7kPDMv0LT
bOGHgHZZHSagrYjTX0EJ2u4FU9lFRTR9pQHZqOVJkkXMN3pfHphvO/Ei7iL5NQACNIBcdq57Dnm5
o/XYeUuXuTnLZ+5Rd7yQ3CSbnNoGK3hClqHBvkAIh8nCtwDCwD+IegqHO/PXmqj4ZmH+RgU3IAbO
+2LNA0DEXujhFtvBhuTVOukZhydQ7QUs40lWIZtNGRGvXqXtxWcJZotiQyUBMFpZGzIjVDlaRSHr
Q3AL2MM086dBpiedyocT8yGHIz4AhE+dQNnLAKndjTqsiZgvlsAka8ZvnR2EvbYFEpOx6HteTq15
3YlCv8nvjzMk4wmbPe8XNs1pWFFwHbdrm4qMtVRoe2ZDKTDDRY8fuhV2hXkCA3anm7RqFj7/lBG8
njJ8j3u+FfAkyy+10TV4ateH3su7S/kCT9b9bd9a3q4m/VCkt7iAcW+Nk57vFUBwuOHGY4o+f2iA
Pckm0sXF54V+wXHcvF3JiWyG9D+GDjwlhtKJnAu0SKKWN08m/JSCTdF/6g2flLMSm8mqHadwkHVm
CIYEpGGs9M0G81ePSTncrKgMd9Y/7CT0G1/VC0Scyig0Z+8mBbCn7uMh4ZNFUovHWtFh0JO5HSQu
HmE4+uCjMdgNGvoeBTdzd7bxQAVCbRAY91oCMZW6X4tv/8CLkmrkUJBzWRB9IWmnL75Mu3HCWB3H
JzLV9QDFWKyGpecoo4sE/iGl3LZ0GLRgQRMPhGyACNJAVH6Adw0Dq3n9uhFEBpedWkhUiNpY7XQa
NdUsslhUlg23dWu/yzPgYWoJ+ZJUpk6AGGi4RUMpvlP17vHb3yMS0AvnpgBHfWZOMwXLFINzq4qL
uV6k+Sul2a/U9ldWbSFQMg/De0aTdoHV+6LwHYrPv7EN6SMalHisZnuV+b/mJknBCCOTDWg6ZPdE
Kmu1SwKSFDet+wX9xf3/VQo1kneQtXy4d4QgElS6PPMbsQj1G2UduMqebnubnm7t9hKYFKZgD4ib
d2zj7E5gvweMJjyI1g9rFF9eyi2b9gVpz6clhHWEhOtXaK0KZx75xyN9Vc68th3/49DotsbH60AZ
/6ksu1OMkNvYRId92VC/E3+Auqz7RsN/pV9FJ9GF6SaMjz3YNI0Z9WQ4Zp10fHWi+hQVCO8VX3K9
YUIFV9BUUN5aah3MsIUTcGn/z6WQMLu9NvK1KlkNIcgNRtsXANH1qFRWOKxhjOi8UtKHI3hOfFW/
GVtUIxIsqO2v4WtAClUolC3y+XgQ7oc1lKqsDqSnTqto4UJEX4bAz707Gulr3VD3ymITRXQpF2nj
hTFzIaPDzmkto8Stm8QTK0H/kVav8UxHyItshwIJ4wItN3QJbKrxExGs1G+9Al2HJ6TDKSpmJGZ9
Nd10p2Jgr/ceBejbq4QJpMW9QbFshW2v+A5nTy5aLiu8mhVfFZ/aktPW2QzqNOdGESr319aui7bB
ALl9onQi2ItKUfZ5P5AZD7jP9WfxSDriVflTrt/t/Q5IABI4C+6+nzB0dZQ/w3OROvyRAFN4pMdJ
a2XmXR1U91IZhjEW0pFa/1IeeJegXGVWvMlLM0uatntVJs8uU3DOP7mKEcZRzz7RgLvDNQBNycE1
dCh+7lE3pozIEXRxiuAtc2A/EUg41cbVKsXw4VYfJa1ut5w+OKZHK4ljpmKP849iTDFDQhmj+AEg
MXtJaQeJ4ZKvKq77+VAR+a39M57Qxzp7Jr6CSZhto80ZxGRM3H2TAeNKiEsEzFfoGiL728UbpAFQ
FEbU4kv2M03q8Cko+ZDVrkAfypcsceaRhDMrlpOdaDbY3XCrGraCzb7s3irStu+p6fpSc/K75DRB
MgUot5ZDaclbtiJg0MvGbk/kP27mZXR6O3ln2YvjtvFeRe34D9QXQAtNBT+N5GNRFq2fvdl+XmhS
cVjnIMTc5HGcui8GRNufuBDJkaFfKFpSPY6oTsEPpRzVG2B4IHcUrTEJpRR1EVtv9f7QCnhYiMef
BSp9NlEhNLaQc/pi2TusM22ZRfehQ3j/go/WT3ynE9azD9lQ9kw78D5pEn0xTSMj6VhREHcL29oK
cBll+9YGKcyC8aC954m63QyGuerWJtwNTH/qaPMajDDr5hbzKTUfPiQnfUU13hN5nuEWM/IqYd34
wu0+5VWo7Z/KAeMwlP8T4pJsuwWitVaKqFapgXWmWlVVpQWoE4K6+PnBg1snmJVvAYV4pQZD1+yK
ZZoAPSuz5aHnlme9Ssi0ZTlsYDx4YsG9G855I0XNnv+5gFAltTHeIEjULEsGotCLF0m9zV5uUlxE
2ffxJmW5Zt3/sOYhX2r4vtEx7AvomAreVZ0/8sYVkoJ8JcAPw4yWHJ/f7o9tK3SdBinsnTec0TcA
tH3XRZthpxv4FIxB3CG8bcaRn+/lzID55BnIZMMzsLLCveQh26d3DfpVxHwPifn/UduqX8cz5SmE
tKfbqoaLwWcT26YMvnD9686s7N+BaUy64o62bpuYDQAIGO5pBwIg49tgl2g3VTgAmkwSDJN53JhS
hC9EcH1AgTuAXHTMaqMDFlbJpteAsg2+1oN4OBhObMRhv/qCi3gvSstUNcD4X4U1bnjWstQbpGMt
GkmtFcm/f4QECkLjmuc54+ThVMhptFr2Vu+oFzBH/RSnvaWEyTpvAItY/AZ5GWu41Jvb3mtgdoKD
uvOfxHs1iE2Ew5d29/qjdiFRUT0dvoU2mGm81UWdDUZU3dIbehLd2idhTsptBcwcnxWMJLk/I0RJ
WMpb7hmnvJEf4BHAuJF++Kw6bu+/lhi+rIWXzM+VvsX0h0rAvQuk1ImJlAw67Gpmt/8m9WvWoKU0
SWLR9bTWOt5rK0YeMsyjKOaVK3lVgegX65ZaDhCSdezHV5OElbydZLOwKAvIxLnCjKojgwITgmUA
GJWgIKR6WuTEMl/IQRj/bk26xLmTEpvbuuycTFIPLilJrL57IqXgf+ScdD54xkJTfmzen236DIHg
Hd/QKUSbO2NBrPe4E16k642HITNEtVK79y8NC1MWzKQC9AxRpA0JufDyVdWvTCyNApncAxjQg6wc
+oi7LFdq1yH9HU9Z1G9UFzdIEWYkoylRrT6xjAKUTcFCZKtTjP8QXiyQGOwWj7TyUz9/S1dbt2G7
p06UJ9FwSZJTBWG+cSb6IE4+kj5jhwtOgLKaiDm96dXtG/PuynQsL05twfDOyZaCscobkYxhtm7Z
+kUHWkI21rls7xvSYMyeaVMzQ4uCIkzwaaQuKRYSLrfJq+sD0sVm6En1XIwjiTZ3nfjcg8s1VkRd
bdGGgXA8rUQ26Pb2kH3+l7H5KvVJni9wKHfuGTiV9nIeanSvxocN5BIIzzn82rPYj07C2E3HyrEe
qWc7/xoDQKqQ2OnKHDhh7BqQ8F3gMa0afFC3jMBqmwTi1sVBTLVR3Cap07APJxnbViwVcXDymDpb
yl5B2nA+9MXLRFUSNIlNHNsSfTeOxBR1rBNcs/EJpMDkTpGkDQ3kLEfsLEmwoarlGdpU2c+Px8LH
Hk5gLEfKY0SACUxiSMuns1YQRMXurvEqMZZ2uezfoR/hv8AKdukQmIb1gaonTVCtPKnpuuI8VVxx
laBo9TfY7aAX+JoDemyg5ACSKl3e9DdnBh0eBDBC7e7vZaQUHFHDFkEBMtdN+uBwfM79C92+pz6y
wv9PiKSik5N8TLLyWc3i2a+ieyfY8kkcFyf/piD+iECqz/X3xBq2L52SN769/Q2ZYEIPEKNx5mzO
x/9KEfmhARXSUYOFZnQ1s76eiOxJq9OiV6oXoEmrMLQLDHbzikylNZo12CR/wqibfVj5pit1sOvS
9P0K1ucR93zSlb23JFP09BKU8gXT8I7F9KCjeiGWe63Kzq5o/WjGTC+W8iAmTotsgEcEHHNRf7OY
RaxirGHGFdv/M3fyk38+qWegTgvdLPr5YXP2h9JW/Ums3+qsJCxdmggvy79RcLnE5CuO/bA0mQCP
dMj1C0SkFrjCmzhyZppjxDTcp3GZ8p2+GyYG0kbjryRN37cZCJ1Jx4fouMWs0DXR+rWCl/OhkAuP
JQdJP/WSuQbc9xmKj7DBWYs7cYXLveTa9DzvejziU5s5wVaXYDaDAWSh9Qbw0ABqWk2WurSTACg0
qLtLRbCk87UpYnuZ9Z8wxLBCFwwGGukPe/24F3Xu09FIxURM8ISxPku7qT5LujCSWd+CAMrnVkWF
5f8tbmEktAH0aiG9I8wS39M6p/r0Vh4yS3shCK5ye7CRDQKLyYdbavXY6LHOCsr0qmKiehfFS0Dt
agamCyif9efSwFe0BXmTj+cr8Wf/RppfVqwHAKP9nBurjOhvMg+e/lxMX+OuSz6d25iPyL45975Z
4be0WY16RWaiSzxErl1uex7LUeUnB3RTZGv3YVqGleypOZRfN+Zv+5a4hz44wI8TnUMV1N7gcjg3
T1waHFqBvemKOORAd7f7CKSd7KlinA41UQH6fk6jXeMGHENFzlBd/okHZNhU+mrJTKWkwNHnE8q4
zo6i5EtKRp79l7YTMo+plT54o3rdx2grGzet4/Ass2gg6VC+rU9AUelnzIeGYUuJ2HyvqULv60Pb
qq1Cqlm0d6Kf6MK448eB3Mb0atUQr5/fMRUlANV2dctkvRVty4SR69VB5ynXp13e8hO4Y/J6NhsQ
WPUpiUeawuYchiNxDk/2Qm1LNoW+wXVVxi+eAReTOvMfEeUIlZMYxY+qx8qM4SIStfRe82LYxAiJ
fbz2/LAn7eZbLytLJP2I/Yyz6DZBmDiCwH82ZtzHtf9nqAmCNggqyV4zz/0uiKtZ6EJcHZfYStpJ
l0V3l01cJvkDE9SZ+vD+i8DucYbnrqH/15yA7MuXMh+qU1Wg2PV3h64jbZ5SolDFbnMF2B4GVln3
jVw3ZvQ+y96Io76CXWhNYuaC/MGATRZLFGTpO8WAxI8xIgR8TwaRNhCWZcXUuDw2wwnV+/k3oG/T
6ZMJu7MCs8hCPTEc63D7Cpj76WpVfai/iiaPXS/h5U57fB7bp9xMGl13t3reocGwWFsfwSYkGkPe
PFDHRvlOttngjLQJ8WziO2N2fTRmg5Ydxb8eHDzr+BWnMkr1b/0YI5x3fofZR7VifkwBO6tK4ZWM
dvXGL5Kac/5jKDARTU4ULuwJ893vxzbEJSw063K+E+2cmL7mBcRoNYkvt6jrJw/Xy6w4VfDrGFPH
Ocu4DkQjEf9bhCjnZYZc47Yb02dv+kCaand1Za87r2yuTZ1c/NXm8M/DKGalobr7bolaj13LxmMc
o/RsN3MmLuY67uIm2k0SzcDKk4PLe9I0SWTdgYaE7bCfeS/a/0PCZ7Jzlx80PyxwO64QjWVEVA/G
8w4gMUK41jbLMdyLd4rIyZstt4Sj7QJPYvjEn9z6AdE6HbpjJqHXejgBLyLxO9AcU7d8TqP1T3jd
oYe48h8h5pz9dtqTejL1pg/XJMY3RhnmCwmjfcgjjru4i2qYSZAXZ6adaKFdSvRmg6o2iA7rpNvS
yzQcQrYb/anauijaZ6Gq0LG8C7ZWxPFiV+PLWQ7SQmFG2+a7wiGIHZWbPMf4ecqrvlYgAkaZojEV
GT2hy5pfC2qPespN8mEWNYLxyr2qBhqLut6dkHaAmSSak+XTV9J8v/KV9mxXWzG+T0uO7vOyFi+C
uJ3WmSyVxcCgzdmb6u9bXVvZdph6tDXhfsnDwXz6L279Xc0ZsFVLnR87Ca7G+mkXT6TJbeDnLIDW
FucU2UftP1eFflJLiXOJzLwRR/oSXFJNHAAF5feQUzq/ZBeYF53JRP1XpLNk5HbkI2j1T4zkBA7F
DBER1YRmK9B9e68txRKw/erIGTubnVLtjGhgoyWPadYJj0agbH2cC0Q/Qrd1Ebul7Ied9lF6pzeh
FXqU0jlOZWifaBph6zu1LGDZUnMIbKmKv8jWfHuSmZq7Z0MJlDXlck2h5nOSOObxG/JpUUZssioc
+W8PY6YJlHVfZPnyJHrFCc5mtQsCRd55vGFFklhNHFWvwNR4urmD5eDmdc/kkG85RuyJNF6pWoC/
ftvVeXnYrmQHk2dhJlJXscx7RJ/uFiZ9jd4QUj3FNC7bLC/bdjVIgrE2ttugVGOLFMyX/iQrEYfv
wcWRChVw9warSplJJXid4wmehu5yqO/mC+eOlJi0m+0zowqyCecIjm7d97s7rU6kXXS6zri7XsDx
87NwaF+BiodI/LDo5UPDIEg+ffn/9W+pfC1CtUfrdridAsqRbS+vQZJGnbWozYrV80bR/kjNR537
PLxK7eDe7qxPFS4ZCCE9Lc+c9g1GvTvdmMPzOJoGkvI3V8PWpsi2s+AhUPKV8DMlBT61eV/7dXAl
Z5IyuaJSC9uBPLFYujNrW78Fcmm95+IVGQok/5mv1Sk+0InlvmLje9YOHCvuFiJy8DYeHGZlbP3u
H5WCTJFfJ/uv8RFgACEFl4QkDXMX1aDUzcrtHyNJ8uAO4ajPw4stJm3SeOQvXcM/7u8pfYvkzfSL
Wc5SauBuU6pnsqRwbjSVe0EnETdS6f10yaKxIUQl/e3ZxHJGsELLIwKbiD4YRuw/9JsvmDOEuc/G
7yD4j03e+IWZxXyw+ipHFePn0tok1mZvoAW1A3hOZYIz9IOHS0I+1OP+dl592YDejNfAs54vkTuJ
xlrebCM93B1T9PT51ccfpA8ysxV90Ln0cSlL/u3OqqCpotzMYie5aWfKSWlT/8AhnSbcLZ5/+D4k
0YEtxBOCzGqOfzssOWRZqeMgN7BAZefwypHUTDwefLNPl87aYzR/NtOFSlbV2WwZVHaHXDbcTOhE
qfd5B2aG6fEjpVHiRI4PUqIgIVxY/8AX0PzFGFIy9MLB1iZUK6y/j4zbptqO4U22Zd/8bgCvTrPk
i2GNpwdFcPkLJoyVAIIdcob9E4KkecZZKhUSuDGAybU31CDCy9MH15nNzJb4JL34Bw3cJnlsDs/F
VZUS8MxFZVtDE8wYQDqvbRaOcCjI3iyIysIhC+Hxl69o9ISIr29+0xf6b/rvxC+VwHBJ9pji5KiR
b4dqFhkbGOT+c3gaazYTtvYUPpNs+u3GROFfz1MOf1J37tNLvGsm3S7X+crlT/I68I3zp6TXb59b
t61q6umqmzQ2WisIXgu3hr/MxB4LW+kxJplXh4h0IoeUBlCjL87PqOZZt5/Z2CnbmY2UzxcqtsRl
zM4weRe8Bj+B5IbzsDFlY86rKbBmc567NtZa9Diz97JBnv8IiMTs88QPYK3XuyPWbkFGZ6SCAbpB
qezGeD+OFWdojqrz2AfCVITGcVt0CNnRShhdjoqU3u2zERiifICpkaJiCh34r4UPY78UnbSb1Q9z
2MqE/w7eitQb8sGabkvbq05isa7hgpbtK8kob6Ndh/uSaRyQSvAGWbY2mzLTUSJovImZc1Gm96qI
I27x//bnsFYcUFb6Jwy5cSMUnkJfwh2i9jtyOW1zXGh5+lmGyY7yjjLStf3kCOS1BxjgNsSj4ec1
9nrY2t2rBjFWuyvecC+S22XQophtnD9V+7hpTrDl7g3xULTQt6BAywt0mi5c8PTm++9U3E65caIX
HU3xffc9r50ojvIrG2AbLHjphLC1mIsQN1DJOo1XbK9b46rOJiQaDfLqdwZSnFvCP3j7opmflz07
lojjmGxVMivzJqziw/B+nK4IA6Yy6R5LENtm+sVQcevR98DoPuyoTKVgOlvjLmKhq7WNn0SwAlba
9UhOneHteINB4Xuxu/lWVN3avq8NVk7rdEsaVKY5Ma6R2gXwIyva506ybTQcpHRWhTwlWORagLkF
6VKmB8QwrnZC4JkHpoNJsEyA0WkARFTQSNZ8XoSLJkhVLJAa/07/MNfXzlVhvfjjOOprN+wx4IuF
ou6tTdIEjOPtHu4v+wLKhQYsKMFgcvhceRMxFYS4d2HR5ycpVh5KWdamp3MpxsXMDShhJ5tOjaXL
72520eDQlRFoAFcWEGMdNmqLGZnCpjL1GqnN/KrcKQ3dxFlCMx/6hdUj928YneNuFZxAeOn++l6v
lgqb3R8gwepBe8zccLqtyF3ywom9kknUaxLxQONTsRx4bNaCv33MIeLNGKsOw9uPygylzCWs6tHb
rt6c3uYwrKD4CA7ZbgAslGCH+dCJ+sDVUMU72DiQTshJw2dS/b9BWi6JTjk4+MmUTox7TJTR3FNa
3KHGE7oXKloJg5b/8jEh2Z+3Qt6YwQHwEsqWZJUb5iiubgMf+utcJgQJHwT3m3vAblnYY7gRbpKW
wota1Nz13NUqBAfDYYQwlb+2Cg/rPnVfZbqOUx1mnA8C5M0yoyZfwy7x3fU24HSXJfHuiTHpfAAR
7ECpKede5SoKq/V4DbTrNa0zD2+SfAbhPqEz45lcHAje3JQ7yYIZ7p5C3Z4AcKrl8h0QJFRze3l5
QvM9p4PcsJTnqofRsThv30sppbgrUwWjOuUtz/diyNi41TJxWz4f9o8KrZl0eHHbsEc4fwsB0aDq
T4EuIHMRGnlIsoWEX2pGk0bhvDUcHc/osg3VC9m+pwct0YfrGZ2wyj/iS6r7LytxNfG8qPmfNSKN
yma4MAhKZ5Y31UjiYQX3K7vPgHDln+UVdV5BrDmv+FFFwS1f5+xBYQmfhf3zVXyf2P5CKTIFqvMV
RdotPhl+07PijfZvdYntdQ5VcDCROTD0gLvzyT0MDBQ3GRqNvWSeufL2mkNyOREqmeSmRWMzW+Fu
r+kgp1piMxH+stDploT3solzPg+yhbwRbJB1GiYXYB+vw925lEN6662yp3BETmlTQHLRevWgN7xE
SSTbDg1YH550TB9zeiy2hTAxW7mbfuTyJmTlaHR6UxrwMhkiqUICwMSMIqepf/FWoBZb3p6a69ER
NQ8wan1I6mli7gUEd1NBHaaMqsKT0p3HPX/k+ZRd9Z2TdgJMzRY+xH5bqnxgm4VPgIHhdlJ8/2qU
xsIs0ncdl3l00vpODOZjA8VvdlbEYsAwqE8AsCN46qVB19KMw3dL1j6cGvdFpMU3rJd4ShGGdnyc
gPIcgt2hSZl9QDAEspdKKOdMgkiNr523WS+LsTMEiqc1DH1psnm+ZZpcjr9U6+yrs6MX8x2i3bLk
So01/XvGmpA3LvD2z6eKmZg/2IqfF4JdylV8dEMaGrjk2yjtrAwzGq1lvq0rNbuPdWLtKUR17YXA
lMWDGb8Fwt9T8uyAJXNkqkWCtTsqJZqi38kYv45+voAIj3XqM+/zG6Xgk+F/dBHBELIpjeVh3nzl
NCE2UToBpM+gvNuUVns9dhG4X8a0lzejA4mQI3h4ESWSEwK7mJDIurmUNA/KBlMgagnp61mAwOpP
20ehSii0/tXYw2nml2M529Jd8PezKTQ9HdZ1EaZvLcZMxLYXdon80VyqcqeB1y99WKq4AVnnfxbU
ZGptZ6zMsfC0apNFXZuzvyOZsxpq+q4RvQzSg2jMTNla9jsxtm+KheDZ01R6/7PaaYoRHnMUqY0f
n0EZOMTQe4rdVKRIS/Y7FC2Uaf5bPZkMZF1cjBDGIDMnwr+/zJvHUlMKSrSMdsCo1k/IlW/cuK+L
Cid3A0y1iMmOejXg/zPg98lO8TGBlLfVCQNfwMLyi3lRw1fRnAkhRSYWdHuGN8c+5RmxasbAhakJ
j3nFgJrR++cx6bT858ZKUK1stbnyCry8x8o0o4INNZi/OJJoZqgtClgXQCKQdNUDg706U2Z9HSXJ
jmXDWdnaTRUAQHoG2BecHpeOYvty1psEvq/8VLl91LsFtXDElPhtZb+9uoA1p7icOlyQs0jSy5Vu
RnWHF+q+hhQ5hrvRCRjvYg1PjdLCPaEgz9L1oIE7dr7jaHKV2UBWtmtWokHA/2KLNXwe0voe7mn/
ec5nUFd2GqdwQae7VCpa5KJDpcVRPT6U1X8QpuwRg2nITelXXZIjgDogtrFGGzQC2yx11gVM4S3V
Y63ZYSGjZDsoMqpGKghQXP01Wr9X3SEF5BYEoehTvzFGM4sMMWvcCbh3Fw5m5g0uw+JYUU7w4t+2
8/KJ6qjX7dRI/rk7ofPUYMonGrOpC9w8h2alXNMR7KH7L2iGhP2EMpRyAD+615ZxhFvJmLaE21NB
5sm/p+7+qg6U4TX1TSe4FqNOmEDZWNuR/yR0EzQHFOT94lgWpFmnse1MlLc2ARQv/pxAg4O0CSrP
Sx8PsPXg0FCtSF7TIKEAVOLRmKH4yzjI9rFy6KRshuHErfkM2FKB3gcogRHDZQ3kvDC7b/2ng4Wg
iPL1o16ciKD0oLKcUf0YPz+kFq3lqK48E5DQ1HP/LxwOiyZqAK7X9/JgUwZUfN+ylx4fXKa+4x/L
dRedRjGWK8cn2hVuBW99nnE9o0a8ZidDUR/Zt5fof7Zol9J2klU7iWd8BOsvcXZV/feAhKFOxDSA
GMW4V/nvg9V0k5tRF20wlNFRjOvfsD02y1RkKTXXxBbxTYtHB63JpTVAUA7rgqH3RsrP4nfP2ur1
pVqWVjOQ4UVndUNOjBLdyI8wiy6wek6s87aBv9pfqzNwpfv7dkSZAL5mO/zLXDeZNI3dLTBEAvMx
dz8GmNKH0t7Lp+oWHcDiKxG4xlX5UTMxwgiW2orETuIbEz50BGAoSdxpb4zGqi+Du4LHPZCTDnas
hzxmd0mBQYtjyJke8Yip0Kbr40ArtgAVos8GPZYwgkSmB1tFgOs42UjdgZMFJ0DphzPTxWoRRh1O
LAPika5kOHHNh9M7uCwTskG5j3SYJVeoamXQVbkt2fsS7qgD0pyMDI3KfAO5PkWq80lqmr7vLxFQ
G9zcuDV7lG+7lkomg1AKE2+qUFkSGJJdkX4Uc09z4kdvT1rkEqy2kjq/INxqXWXp/K7jCqbNnWWy
Aquj1IpfbWwgo70q0KM0q5F1PEe/JHIftKDw5cqglhBzDbuEVqHudkKuNKbVyu+rjJK/fW9HBH+n
0gfr5JrmSLk+TaIRqW9smvWs1bGD7EU6U2caDvjp2T/dmlxd/m+pMDycx3iI7TgbEBWjYxFK2cyx
MJpgt38WH6V5zmqoJvDrB/8HrFP68I8bCSWd7vKEx93K2Cj4f24f4Tnyq6s73i+tcq7oDC/3QobV
ljCLpGBjiuxl8nXTGaBZJpej/5zfRnwJh4RQCTFEJfvyd3NYb2VaCTFDoO58o2gotlaux6O8evkp
N2iaMaCWE002FiNMpqRKZ0uVwSTf6W3+i87+vmXdMH7+Kp0DL/SUhcSHhzOW8CufCFfepjjhb0Co
xXpNil88LUT4APsc3Zx6DgwLad5CW1fnwWkfivUq+LcQEW7dhuwb3bpOnvpLramLxnd6EKoXUe4T
4/UIldq/oPn899kIbYcvNzJkiVawammJAWo+UkQJKc6sAQPQQ3hn5VNQonmBZ/e/Idl4q6kyAfmv
pZf/IYcA6tG0l4qp1CNL4yMlf6A9rN0ig+Xt4P0mu9/g1Lmhmrn3mHUFzTRIScT10i+3+2pVKsBO
Z8sRNyqmx4WvsbWHnSbJHjnM+OkU69AsYlFTkKl7cHWdZ1KqFoMFtn2vnCQ76KOUjZ0GhumO8d4t
zZJU2IsIBr8XSfjdJPSM+bQvSobqMQrHUmMusnMEu9R00ZQZMMr6JZgR9yEn3ULkGfeufWQ9Pjku
hTnsCvghHP70c1hj6U7l1y91XUEIwES0orlq3z+q03aYXS/0HyEfaFsPcU/LSUNT06quKDn7ktkd
cDu4WzdprWVyK9jQ3TKHcu3o01OAlKcnBAzjWzEgXcJJS3wA1pNjO6yUmv/BpKEONO5kKb6LwXUc
XLJkrL+o32Bc7UW8cC0i7+Whgrey276S5VgGLlityFEDKfoRo2QRPJ01tffRwPpBvenOz/Z6lO15
giPDQ+SGMMeB+56kP5U0CIOs0rLgIkmdS2mtDbUqrxvpUuTxe7n8jbmLvtKRg9ktlCCqPXKCA8tg
B0T5mG2yjia/e5+Sg4eoQCQ1jrVc6Nj167zEAL2WCwKtoBGWglWbI+rHF6G2Q4+we/DSSeNTjP+h
kEjuwpwHWzARS1/YFIh1nHg1loXI3BLUHD5OXsNsn/bzne5XNImJYDnksaXR4syLHJ9zTkDRuDHp
GlTMNRfPepk8Jz46t9zs6OV41anls5tKizKsKa7OYOf+1GVRBIyuAh2tbuww6B0qnQ4x5XAnitf2
XWQ01P0xu3SYZq+FMKB8xYGAjMtm5/x5oYMQC6PGaEECkPosYFgzD/LIXsETtUvF/P5c6EbOa1GM
GsvRtx6VcxDBjVf2GHFmIJAFXmvwbLw/033Vr2C31h9KjrCRcPqoflMSxRPxZa0sLU0z0O9gdVaW
NKzFc8yW+B5rybbUgzt5MgTmUPYtrC7S3M8jrY1NMdVUarVMTWGiOWW+fMrDN3c+rxcUZEaeXWo6
HXYKcU2uX+NTA6Y8mhbP5PtBYcZ5NEeFqs7KM/XkLm9cYN4XDdrWb93tfvl4DCvJL0rdm13qnk2s
CjKmqkIdLmxfWuqwfUzg4cbeUGXNxXXxkb3e9NzgfKwBQVBXeTw2nbMlAV8j+S4mIrBz78P+8zV7
HidSaSeMkg4kZ05UoHstSI/zT6tqc0+nzIdJSqtK3pT162UGU3qY8Om8ZOvxbIxUMI7aE4VLZngc
A4LGrnLQaUK7LaNvKWuQjFZGSTsJAQ9iNJqrOThnUun1sNPRu6QvTMPgipjsidQU7VFYGITjiDvQ
TeZVn3XD+FcaI6h67bo3gG1j6qGJQpVHfjZ61G5o0VD2SZcH1HQxtD7DYcGUc+WJ4G1xaePf/Atr
jN2SHLo4XFbSPJQ4s4CAXb9HpIgd0BCu7mvRlWEVyIxN6YDkZogz6O8vQO+m0jrJT9aESkPeCfeX
vSPnL7Q/DIW9gTvgHg8sPwJpWJgqj/H3gF4iDo47q/5qXHAhTWlBFnbkcakawTMMVEP/IY5nh4Gi
8aI6Rfy582P2ojTypmGQIMNTaAcZne+vxHRO5/iWlmOggc3q4ytiG7UAGxYDiMaXWOIdOHc84OoA
YnExJNx/A49wOoaBjviHIVuoLxjJIxrUeYQQIMSZ8f1BlMH5NE9zO6bOXkZYbuVVrXa9aZ/cgpyW
07+v6qsw/uP0kAibQRLL3ZC5Fs32StP28d1TiagFvvjrCUaW0uuLOJiqZZlOlHxQymQdH5qomMoW
a57qtQz36UZ+3AosX+qVRoO0R20zczWvQjdGrBdwnndpD9ycweV+UMnynPfdC0UZk//IA9lZeB5c
aRpTGBcHC1cg53xDGTOXD+mLbyoBwKXvluwf4dPD2RxlTx4gFMZAW3X0Zb471Vcgol/UrGksvaG5
EiT2fBuLgaZy5aJCEmd78XK1LGmt+RBKxjD7CALZQiV6ct/mfh2bB0s2T6C0VHbELWUBuWImwj32
/aEU52mWYvT9QYlTBbdHxOzRQ4i6jM9G4HS7YkQprPWyr6zFbq4Kj/y1+dOX7fDsG88IPp8/OUcQ
/wFdzvCNK+vVLWVC0snf8N3DY5fYwNXzw5VXUoRduBA+twxzNLACVoNT209MGXo0SovR7VFEg8x3
TgKzm0CfsqgPPb14qsQFX+ZcTvZs/OjUZwwyHtrFb7kX1p1tvyQIKIop3We/ZjqZVpSbw9hmz2ML
E2omhN1cbNz95uBNsMonzp3DW8r3bX7Q+cCDWWbWi5JwM18fG4iJvP2Q/Oq6A4VgYysKL6rSSF4I
7QbAIlZ8LAq19c0CQht6uaFu8z3hAwqjFucYW59pZpdWbxM4rHciWqTpad2gK+WIPu5T//0sji0d
SCwykQe8q2VGrSCWMLczRbdAPgvz1WDLzVImclyYdesTWyC8/J0XpE0pBrVwivex3mZpco6RHW8f
0sorS/bLs587hVtZL3gupgehdMM3U4vKp7BfcPw5UL9HhhZCCjROI0TCSHrSjbkfcRqc3xHbhldB
ysVlJcVg/XIasKdHDNELy1y2kPu+WIoO8hz4v6WH7G371oBIWYWDHBBA9ggJHa1Ke4FADUzY6eak
ZjVcrdd/azapIRZe9/Cuxd1rUJFdd+u7qjZ4fskPzxPJZ2mdRnSUoYhgsbgU3aaTMuiof21TQ38g
ujxpnqTXBkg0gG3Ga86tCXLeDZzfqnS7rC3fqYIuTthZLC9ruwKc+oyhg/XAsRWDPz3UweHKOdIR
bt41mjpAbfiNqHlmSCVKGskMOErr3hNTtYL6vB+duJzfzclWEsF00ZE3w0ohfqCxA1MjL2LvURTV
h0+dHuLvqrsU1PD5Sib+dGAnbGctaM1EjtF64X+YuJb0V5fRrGXL6izPgeHTt4KrDaJsgYLPp4il
JBtWMShFQ7wblhdRMY3JrOQTbt0YxSIs4FudGumSffSg4eiOzH8/f+gDWvdiWVJuBeuVZlwlw4Ow
IOy1Y0z+4DZChfD6zhsmiFhC8oEl/efnwR18b/cmb1dwJiVL1KSzSep7S2t9WiPoa0MKC503jpUa
J2v5yEL6da/4K+fDFfsS1Jg7xXQvTdrEVnNsbkSdeMcnXnq/ayG6uYiTJQqzcbYnGjhKP9HqpXE7
tJB8c0OZFj6sLqz/M5cL+dEQ5LQug2xGCZqTNs8PE9pQOXYCkCTR88O795TxqEUeFynjr4zVvLU3
cAXexP283jCteto7zcLKGe2R6Ydg/4NhQ+RYcVRliOBNxZFkY6J4uKkQBRI6Kxo6mYVkoZeZnvOd
kHv+bAJ4z98ofzjNO5TTGA6TugY1XNlIN9gNaY+k/QtiYPT2/d1ZTlTe67FA5Fi9CKbALqZLHm3t
V06UgdfCEzoyZCK2NLyE44i7dIC1CmDOoc0N0C2GQFkIuTVHKILxBQzVLcuu0IFAUREcZM/eNvZm
KVUb+JLmSYGIjm1DKbSKOI0Ns+yumhH0Vx3i2C7cASZK8qQ9xNGLUW9imT6ZGKt9NYyNC2TO/rD3
iayNOID+ue1WbkFkD2mp9kOxItsfA0AMK3VyfnzD8JeElk7m0NRX+yrCztBBbXgQPwqZGSsmFJoe
aGXAZLdffw29mDoG4sbukKyh/L2Vnvy5F+VM2yImUfqcyMsWohSOqDp2rsUAFy+v4QD252hMhhOU
X0beMIhqQYA9HRjmjAAgMJ052/MPy11Jr/n14vXniwEcgGXi7I4kuQ4BQ48wkDFrhSeI65UxVkkT
k/Bgi4sPN9S6w4bMWoem+ZCsqPcRAIuW02kX0jCk5E+v50iuk8pO7LArpQ/joqWh4xjAW5dhed4O
Z6nXo7MDp+t5lTHu/SOlDTRBOYdo4dftjrZX/YT7tflYg9d0fomXxDponZ71wNK36Or4obc4/KLA
2fHp0/l3R5dmVsFn4ynZUYf6LIx6s3fLn4lvjIgUmcR5Lp9aFrvfLfLzUw7kBrQqwjvEUwsbWOMH
BMIasqX6x50EAUUtu5HS21/vZIo1Y/mM5JHTlPI5DL6d4OQ0HfEMIPoy68ebY51v0OMPNrftsBUI
ucoaP6hp1R7ahrtedSQqaH7KZr7ggrLqtpTK1EmuNMy1kknHhtQFyl9h3SKykKRbuKrDU7rNc/A4
NRc9vNvbam/mRYH2L93kuAptBlqOos4lKfZrgDpuYddhc9KsdTa/pznxZzgsYmN5fgSCzJeHEWTF
uHONScKkK8cpUaqFbMQlw9virYUEXDHsRXGYSEKCCQfhzG0JO7RZtaiCJ+TtSYSft5OhoA3JNuRM
Ja5mDz9KA+cnuZzPvCwPAoDk+/M9f94XforhZyTYHtBeueb13jMGy0uRgssJUz9aMtjI9ye0JfQe
wyEmuLrU2ePk4W1xgGOhA3wiupJ+j5NjPxhen19lR1clU9rv89yU11z1bRHy0hRq3znisMimzj36
fdYsBikFCBEBEew+prMrjboJDtWLN0zGjlimvXgu/h0z8qCXqzG0Cob0DMNVaHiKGfN78W31dsOs
+3SG8NvuN3hUF+l7myZwkYHoHDXDqqsLORG87Ef6StDcBgHOeVZ5bqzCIGmk62+Mk6fpGDfLK1px
MNmCAx6T2jveZT2mH2vzoF67N4qTKSSowhvGrfVPuck/GRPk+68fJUhnPobVdrB/C8FROGu1FqZb
Y2C82hm5YsvLdKojCfILfA4uG6elwY87BMz5uc2U3KiKbLL6M8Tsgs8Gp9nvHr931tjN5FWEp7D6
/Wy0+SPP8N+CumopE8nD1jirFaW6eLFvW+57+isqnPcRs9cFhF92pguja0qjKZAo8Z3uPc/3gBsY
m+BausHR1JjsyWazyTuuYwuwn9fPTkHq0Hiv0uJv5KGghg6wBOCiuwPRYw9ADs/F2MOp2NMIWrRM
MxdRwUR9+G3vZV8VwdFZsceizupHzT8R9OlJKPZnWgkfQA4voA0uf0avDsOJ9ung04x1SBD+VY9/
/v+yt/JnzStnUgLDgEoLEIY6CZX5rxTWLglHo9ryBi+IOBbxwUO9v6cuOJk9ZBWO8Le2hw24g3fm
EKub/jNAqApsoW+U316xOAcO5j/NRh6ZlAuvZwuoVt/kGRGYCm2ma3DoaWBaNzcW3BE511ZD8QJ7
9Gud0XHTup/Ta/eMcCKxPe6ufzwyuC6sgvWEJAZ5CVV1Y361/cDhmkRP3Hs/iR3JKTTV7cLUxeDx
CnlaK4fHNU9AoBLPNIFJgq+CBXjEwm/fthsbo6HKuKzdgoPpw/RqztdiCkoEOjOgVEW9ZEEy9Xqh
RfYjUest4nVPctyxCKBnBbpyQmUDRkqAxkm9xzXDzX7HGH5522FDJC0744Glsvb8Hu3OQte011jA
gPgalTPOOpX7+x3OGcFaAUJfVGxM5AERbpTAn63wRAJNlm95bd3NuIJSGhBypVdPUhprqbexX9os
+3tztFf7GEskVVyxW1U9LNfLhik8KswLDn0IIq5rJL5qbrNP8JtjT61YQjfK947dgciUHMbMBAqr
oILb+/V39QpszfY8cSV8/AnXr5k6m9feVaSwkp0n5PBgHUFptyNqamD45mpsl6asMp/CVtyLOOQU
jm0GDpoQvKuxF4lb57ltKNCWKn1gqO48w3StyunGCX9Ck+JEvYdtd3hsMGwJ63+d8kmVL37VEtuj
tVB6JVAL2H2djw/UZIRcJYtQ3dtRXCLZZq7s+RyqiGQI3UPApwFY50JM1in2MD4SoYwNBKRfStkX
Km9c4W/51z7z2DHnS6JgqEd9My1FH2x4s8NSdfnaUER1MIGx3kO4IsKiCJpZC/5icsj/VrpLCQ/7
yK4SeEnggRV7BpLUetQdkPSPwK28SsEfeKnulXqgpQ7Uw9cATMmFmInJcalLbX7Q5myN8jyS+mSB
v1YdWpb2MwZKTBYdYdQTYGe/l+5gIZKvERSUUtXRAgu4Ek1vvkFA7Ch64wHfGb3qiMH9w5xQ1rfO
spqu83H7SoT9H9qP0XSFOHslM2ieRUvbyV3JmGlihxtZTjzZkIpV+4ZtAXWjAmgXDWSJpqVjcmp5
akPOZWoHdTWj1MiCtuuY6y1k08EdR2Y+M5aPmsuV5ZANr2ZtQPLqF0vGHh+9voLPuFtYY8pR0o1V
HkARh5/BQi3UbbmfT00IvLAvzx9QieX2z/0VcPn/TlFXIW8eq+cRcy0WRcD+K5WI4dqmUhjKNcRc
aClM3Ji0iZJ141IZhE944zs/A9hS61Lkowp8Awm32hUPNQNNghih3p6QG/fdMmeiWXdPde5NVlMj
+Demm8MjIVA6Yn/CwfvyHFlDv9NSLbvC4cpiz8xB11aI54Zzhou+haWeZs8zQvsg3hUHq8YK6zUO
8IsDpppDY4aqwoBKcOWW2PVYk+Dt82+T8khNxlW+N+WdAfnn5I39kyYGxbPqhrTDlx5B2esZF7+W
NNS8uug+5bYz+aJi2TyVxSOX9zXtBbBWfU/3dGWh0V0ac7ujLIOSJhagtPUM1XdrvSrMjkts4tUy
v7j5XQ/Vzvxpn/kAMtycMjPBAsYi5VtsYY25XxuLQ0ucWiweipXAo5atEudxiSIN9lWljTtRfo26
r2sN7AhLOVpb4KR9QCuBrS5+Mp6eSbbvNcXhp2cu6LoLbdYadpRchfWnbcioiwdTwMqfZl4xt3Ze
9I/lvDBfFQE0onD9rFrXKOqxKwAzssTf13xfshaxrxdFuQkjN7nMORy7WxkPG29v4lF2eqtr8Xiq
FsnLbzQynPjLyIq6gT6QeBEfO7KJjYf2lfyh8DgDNT/u1P3oc5mHG0SVnr05rsrgVaNbbTsS1u84
QXkaSaEjl/y3btERJlMwAkDjbys622PBCmYv8/XFtYxMScIaVMUI1rH6Llg46N7AK5MEbLhONgZU
AuWmRJbqNlhPS/zrtMHdspIWlFpenc2ZvOu0TOTGPItBiGDgGMRoEib3eMej26trjddsofoqOcMH
DFRUwKnuWRV/h0bXnqZwAYGj4RKJuyo6L1V5S+0wmFKeedzMUsoSogQn/hGYzm9J4QvwwXGaR3gT
kfy/OyUKQLrsAwU9yvrtg0Myqs4QxQwVFxiL6kXUquCOUmS64dn+8iwP6nVYCFSLwi40ONWP5JLW
4AMXZNa3L4J6Fjvb2eu2I44Ub6+msvBWIg2WXOJaM9rUM6XOxjWOgDfdogpBkGeMA38riMLp55W9
HJbD+haOfa92hx2eg3rVHoCHB8AtPJZ2SFQescfSOU4H0rUXnPa5I1swk1OYAkcumADxHvptMdXQ
Gh3dnHhF9vxZHgkxzWdb5vCP99lRyx8QhujsxwpVR5OyYstDt7iZ96T4gd0WlWLmw7e+gCzX3SHe
a1BXwbbRHjR3B8fuJVD4zKs70rSTI9Zrp3vZcXpEDZG0oiF0RLSfm2qnJW7Pv6jGlZq/miWQVP7G
ecovYPuWgmvmGs+ExrB2m2cRVkU4EhOtlMSwMHHEue8+ZZRi1TgKUAthiwt/Zar8hqsnNVTN0Ca1
h8EyE3PJsVcUNTG6p+qvgqEsNmlFw7EuZi8QHBcQnLcWOhceHhwA1Wxz37mYnotbp6GQkC8oEVga
k8UFRSpGtoh5gt9da7o8osVQnaa2K1eHoRQKvx5Aov4fOEIUStY9+gEoQPD1oFoNdorvSpN1Ihg0
7VE0eaE58inricYlYdWs5dcFelbdbpxW2BI+WW/av5Oejg/z6dg9bPC4XH98wKv1Odeq+z0z6u7t
+YmLjaTea1emQoLFgUQE25Z0S3yLxRHRdnjWVOMI0VIkPy9tsMZ88qzDl8GaGQmcKcPy0AMKtaJg
2CRosvDq2SLA+QleEDYa+OQIxKyYZZ6Hu3vS2US0bgNUi1kWwHMWmY1KgJkgm4/EuWSjhqzcuTNU
Ud53twrGIaE9rWeC8uQR/Q5Swnb7ZnEgDCZRFkgSPWeVcqsTSKxYiultO82n9Ces0rlxsycxU2oL
jl2PdCAHF5QEtbqVpOFfh8O8Tws9+geu7JrnjwGiujLCp8TuxIblI3zRCVBFmI/r4m8rTGV5y5kW
PBMSv+TbliWeSNlnNCawXKONZlyxmrDUcwkzElRPxaonbdAPPw3an6dUW1C5PJptkCpUHpJJkYZd
CadhANSBdN/i6Q/w0qOhElTnqo6mQe18oGdrgYtktcBuJRHgVIftaluypuka8aEv6AK9Lqz689Eh
49I95sdrcScxwg/XyyFkZdM3i249h81tNiv2czaGGz1ZGFlUcrv/crAob40fw/TAY5qqS3aZ7vBy
GqjrYu7tY70qHlQeWekJfv4CuyyKHrIZ4EM0bhVgbKtjfiRbG9cWTBjBgoNvHkov0ApQDNxakuV0
DwZoobrbJhx+8yk3uWjXl2fgX3Gnvbv5NDH/E+s498sWfwlRZckDDrOsD7uVzGz/I4fPxVG5BX/r
q1j7YOkjz6HxWlgjxOs50aMvbFKQrMUEY2TvtHB9MO9XDFTZXiIGv/sEYvp5/gbZUrWp40KZEmoI
DhANCotPCmOejl0ASCwSgUIT+d4QGMgZWu0bXZm6+xVwf4GikOBSksR6CjmhtNzh6jR05cKG+t22
X+JBJLLG8cDrs8wQYL5RxLujcPelwe9e0t9Omyu48W8UEO/kYpxd72X/F7eaNQl8KCIkmuSK6Qbt
Rmbyl5ZWLbUKygJ8j2ayBbTvPtDILF4Y3epg5PZPn7kyTGtk58zyYE7jJ54eZ5gVq3pG8IIVVGMA
LdrUHqA7sEuOpwFrq8APKsJquy31MqNipVzjcO5ohyzoFdp2E1mEkfFYubSs07FUJnVka5HwO3e+
qe9q19gkgDDupGu3t9kOdcrZPDJJ2FeZnuzRTOl+eX1SYzD4yIvAj5N/uYcjQxkkyVAtqQBGGwi1
DnWja6IrRD+Uc59Ecku+qrsfHh53s+3743OFcS+UvA6Dd3nHCLRcpt9HPNkdaGDNi3Uo5bjTJTuL
UhGekevNY2uQcOWuM2+e4KF+L/tmOTV8qasznOj8wRGnSyJ1mRTOvGQZ1oa5tUQCISnDy009wG6N
z7vNwz2+G4wQ89tXY/jjjjUGAmf3yR6JrWyPWgW3pdeUdxdhJCv/B4VLGRznfqOhFz/dZkpZGB25
EVq4xCXKsEBqeMQGjIm6o30V2ZulKRsbwr0LOUEQ3tGcutVDzW996fNT6qpScsWmLAYrHaIqq4H1
LRApMi4pRs5cXGbvimYPfnGWzDutbrvpRHY6EzdpEL2up6oratzruSml80Ha/UIY3hml7LdPhNs2
schrFnEeBpppNjuY90cZ/hBvbfj8gqA1j6X/Xj/hMDULDxZoCWVpk37jEk7gm7rr6rpAla1XIe49
uALae+bn997UyIQfG5BpHJSddS4M7gCBz51binvJjCEIEXjKYlL/ZioF+uTZoTyQ0dGOQndS1dnO
7+zXBpmebXIXoBd857x9bb2V8+Sqn0E+bXb4krEH9E+ffF2XnL7wbVgMCdUNlfgS2Thj35YohOQe
wjWSubbSog7rmadrvjlVV8hf5ThSyqwTkGxXMYQBAzjbBYiG2ahz7bV/6Vo5RzkUS2cceq4QKFvj
umRON/9Lp4VRsmUzsaITUuM3jrcG2Oc5AfQg7gKwhOr74q/bDkpC/obCApeTjUynbpcI94A3NWJq
s+z8DctR7SRJvcJwAqQrBvr0B0/G6R1H9EMkmHUW/CC/ifuVctlkl9HGReu363HpfxtDfDRKG/Ft
QKoe4dFrmTxzzz4hUCwIt2A9F8DDgWusKLAJoGAEJFsXNKsF6t1vE0DD7H1a+ZFxzxJfnmL/+QvN
VprjZN2JEU7LudGGWcemExfJrk78QbgrbmiWjSTTC0DlTm3qUOgXMSikE+Upttvp2MaDCux8dX3a
15Oma/JS8ZSpZzwoJUvaigGxio54UdHQ1bHj0OuGaXwZbAHh2a6oIDDXEPiGEs+nO5qXVUYzefyg
ZS3PImuRwiSQsVQrYj+yTldMVkhtJdsVvs3PhhV/McRcimjWtKcDatRUqakORwLT6qzP1OZGnJ/w
1EFcrCvL73NIF4QlMF6ATJxAc40BxCdIe0syq+5QMOFW1WXezXbg6E/77nkGfjN7P8OReLfqa43o
4sWbZpYrByH0Kp+YlXGACR9Laj8VnlCH/xB8YSjZtGTuQE8g4ESY4ANQfoNZKcy5Z553GX7sNcJ7
QjFZg3Zj5cQk/zHIZhOpx1aK2bAoQOhd4hjHo/ZOrA9oCUg/hbeY+Z61zRchfwzl/L9NdHpCHx44
R9wMk0U9uU+xMzz9uh5Hxxev5pZ5sf1WJZZdH+eFcM9Dba+WWL5ac+tWSdakVEleUjJAbeFGljR1
fumeCRLO9lbHT9hnzUe32FI7YWMOaJ7U16PV4QNsu6vRu152YRuJseVuwH0rZk4QmrB53g/1i97J
q4Dfh+1tGZj6dvV0nxLfOqBwCVaswWNYuFL6JM/ypEmWD3LnrwUYcNo4jRsF1lHF71ZRdp1tJd5j
xKibd/iiyntvNGDxI0q97YO+uM7zrtfKzCa1mbd/lncg7ruckdg/IlnuvOUIr2hWSJR+SGYaW//4
tS/Uzp09X0KfnAW/n9aa6mcA23PeAxuxSer97/R11aBJ+ll+JoTu3bCjmIoVFu3lklrDu3BQ6xRd
HYoxS9Oy4/E8O6ytVdLLnyJLJI29b2JqSKMBqh4VDF9mFgbPUpHaFKnRhilb2dgT1drWv+TsMwOz
HIFjOdhZo8eqWLnqmbnEOCSRP/QeDAm/VEeSCfXCEkf1kPRa3QzoxQRFAcRFyFSVnjTp87//pLof
EWZPRKEMuzjm2MhlgLnaKYFDi1vvzlkgZwDJSkvV/M924Ptpf6ujhmazGBb4CPYAlZsbNcuB4EmP
Q5w1GIItXkkU4mPVafotdTSbnhV2cz09ePqn7k0qLvKut46i1E6Qf377vCsrdo9BaMgGsgoeqCDx
/ome1ISamk9qYb2RBK209xlOlTlMdYD1s+KOz07o0OMPA8rN+al9RYjJfj9LbbhYPD4k147Gsi45
e1k0crFJKa4CN6zEXnpr2W+aPxj/r9VvR0tVNAYS1xj3J7aJkU33oBUXMNHDQhcc6dRDpHpwjZeB
xOO8MQpL6oPVny/Eves9KGzR+3XHU+wRpADlfFpR8aWZ7APXB4EZgBVlE2KVoEg7dJ7RExX+3iQX
PnoFd0PQqwhgXmswN+l4sZ5mNPSf7sjU/ntTWrDgxqQKQjDBj63dCAtE+n2ZLTaxntGH7H2kWivY
Zls5okZ9ycFJga184lPriNLFDwx+Dpx5TVkdpIoENW3imZFCDaGgsZFIWhNwJILAMb8JwKeX0H5N
S4Kzy9JbeF1F+euJRDZqeXxMhOqGj3xLjTQJtExNta+mxXVNVTspZNEim5wWVUtiXwg8bB1jL1QK
0nf5CFXhVEwWH/tjpHOCUlxSlguCPd2dCCWQ8gjUWYBPqoIUsVvW8f35+5noDD6B0dYTI1C8sUeL
ki41YpvXvjw8NRvFBV3cY7vjjEf6RZHjbYsCzxQG72HBJkNyCXedKf+yNbhza1nbBprRUwDqpN36
0+33beNVk0re6WAfdFNA0m5k2/Gkj5iOWA8mTRqP1qjBcc8OD7nUAL/CoyfO+FO8Fhqyn3y8pWeS
JZR4zIzvu3fZNBvoHGFcAxxjp7HxLbTTqlhrTJ13TucSDHVESLZgvOusDvCngcfS9+ewN5gDAUEW
Vk5DfZ9IlBdBGtdi+912AsSYGK6niGTIsYVa7Rf/3Cj4y5w+DePz8qz7odILqo06GqBNj52rWJKi
9TRTjdxFOCGMp3fep9xIrfRKeGEeEha4juRc84S/UkOleQagIhgqt+FVGk+vXskji+WTNRjOGywK
Ti9oAITLIwWj1keYaHDW6YEwP0CEJhZoP0YkzrJ06Ag02Oyu5DblR6YUsGMcyu4F+leiG6q2+eIq
KTTy0cgeqiORqqZG+B7LHjtmjmC4Gizo8IdT2hssEr9wslYlNxYLCpMpviJp3BeSVsc3hNrLmfwz
mEMo4ugCXj8tAqRqqsxrj6ECGTuc4K1q4mRILzFB6maJ1d+vvlIYytjvRaa7MujJSuDdWj/ooGcy
Lg7mBk9j7H4DLmklWtvP/iY9wL4wxFeYK+bzteWFMV8lxLT0m4ZWOE5cnQ4gcQYAoCA8CqqeDZMf
lUZoLrjdXmKR6LkY0Nk7WMx6Dhw/ZH3iAewrnQ4KFp6KPi/wcfNJtVJUqmQvEk4SPNZTWufqsdZd
Fua4ZdxjV1QgtAuehQHR5BnJ1xX0wWCziwQNsEcZVWHk8Ya7UglRyqBx9exZMOsUhp7k4zkJdcmF
tZvqhI8YHd4+z4xP7TiUIVO6wiYYOEgh0F3uYtdWK3U02pUhBYCSddf7RSt5Yxmrol8hkkCNKMpG
9pbtGyHOBUlOa0DfpnA7N/D9JWBUpY6EMYMLi1E5QDQqZNlYLqNJFC5gXhOiSF5etKFPmpPLRhGi
vp7HQD28Q2DNT1wLh0aZTwsVZh/0BnflpHLd9bRaZSF5mdkfD/DlfELzTUAuBt6e0PcYbHKpcPVH
PkhdkmWtwlNCO8QXQkVofOqqeBL6Rs+WPCwp2gr1gcg/NpEzFxelD5J5U6jCSctQexu1PaTGYpvf
lRJcKA5U+GjRgWbnqujFdeNtQh6mxXdWRL/hOpEeW1Up163CzYeK+ZwmoMrqCL/e7tHAzIC4ndlr
RrStLpOvwdRHhl9bnlqlsDm76kttyyIBVJQ2jkjJ4QIyIoRIeVKhb+FDt+vwmNsiSiOn+nEwU87O
6bRSdADSzK0rit0S6CxpXeDSDpPkCraoRHrEHfFhVkZRjdI7s6zPXu+K/larb7+tQDVHuSU+dvzx
kGjpTl2yqlphThO1H2kFdEBd6hORirVAEAamJBWVAHVg3+PB9RHKo16CIFhM3sEiazF/YXGTC7bp
TGvSSq88WAi6p4QCjrwTE30eu2meb6DH9vj3NP24iKs4sQw9DEFPqyns9ZguVJkdJ+kOi48DYVBs
DQVp0n9WhmmOeFVV9msg2JyGQaRNcwm2rD3qcNLQbfH7FoTFBeNJgQvEhpOFDxLolHRZts3pSLHu
iumWtWjHU8/WyQ0suM+RoS4L1o6CLvNBJUuGbH1o7o2QVDk+w4CuwWPZAP9o59BqpAneucIy58Zm
CAHaVkzu8Oi0weZGG280oo0oS+9+AeyU3dh0Td4JsiI/zs7HpBIC5VEvP3dWbvNUekORimW9bgpz
btcUysf9jwJCclSq/DkEz9H0f5lURQBhytRWTFbouqEstT8/TGHPRrCLTVxjkqRcLvKvqXuJCskq
XE2nR1q9hhoWwJIkXYI9kHMpYkzXnqSKeT4u/qbUVa/j56vbrwTkuu6A5DGrF1DWXzBS4KiuvlBP
51FzMax27OgnrcgNmVv1oxpvkPGfQ1aVF/ReJIg5gh5dJNNe10fpOFpQZhjp4ocWFo8SRc/rWkE1
qc6zjzZzlPc2bVLbxpEgfjqxpntYcwYEpLga/FSUhwtSXkMasCnOK2aW0neq1Rnta5VCT47Pc1Os
W3vcnVu/jJ3WRp3RcJT2JgwBeO1SA8yemDZvyWiz3qTnUQXY51A4KUjgkUk5jSAN8rRQbRYhqELj
5diGbgnvjeiMGr1cU511ko6zlfmldbTcAS5eLpkBetdGruBnejbBy5TEqCr8oBK7+rjgWQG/edmP
2RlJf/OsSeDiEHzNpM5Z6aYP/39GqXevEz/in9dr7QiVsWxT6J540HZuT08eU+yUSwqgE3PqEyGR
FKElrYRfqlKwvHsRb0e5zC3kEcpaBXe3WYNT2uhiJ6WOHL7zUHDstNZFwIvSMmQhF8PHkOGoWeJH
BiaSRt37PwP+kiWeV1l5y7s9N+l/szYnxEXfZ+z9vZNUm2GOKjA4KBte4G5rcHTSwqOuHcFarSUV
/5OVXdWoJDqJhgaZYULeXRowz86a4mCyOZP734O1jOzluKdg8L21ldfXKsICienDfXduKYNRg9zf
R5GETMoZd94c1IThlGkVSYSsBD/Tt6uHeYC4YWGPU0tG+GMbuXlGBzpdwr9+JyeawuBhZI4QZqNb
v4kfkzONnVEW2QtNyvhS44n5df189ejE55P41XPwBq03UaLQixZCcsbw5IyRyQcWtqGuUAfd7q1z
TFtgfIEaDEXpygDn6aXY4NIYc4xXVHBXePAeUvScwtNj5+71k8Ed9/aGeCDaKvCU3RW+8qkTp08P
L3M32x0iEdXIfHNn1zWgUB/FD5uPzkd3SQPf5NGHsmus+hskMmsQ594jeTo0S1KyRym/qqmMElRn
+7HTjblAThRoua98dmiW6WxlUd9y9mdvy7kDPaPN1KF12mx2j9K15jy+3ANfJoDYuKe6CRqlWeBG
pKeWuJvCtrL5Ga6XYjnjSizVuJvQW5RYiJvFlhtuWBOunJzyycb3X4ZSm7AIt+ZrppbA9pNR0EQQ
D+kR2GQnRmAQox084lNVT2cgKfRjqw4+lsPPdYgaXD3QvXTaXetcQkM2WC/Jb+fIVZVcfpGZ2BBW
GQsBB5Gcz1xd4ZBCla/N2PgZDYy1ar/dz9fJm3fJc6muMp1NYSTLBWSHutTcp4/GjDv555UmG0ph
o8wn+RlC09wyly4HICcefdM/7Hm3/oiAHlFS1SfY0wLXobBGzzKRUSo1h+hsBoXsJ98n4PvhCe3n
xYeBXN7txsUrzrqxtrEOFmyJ0b3j2QAYzssvJI41VMrYAjRxp0umDyewFJyv6gC/wEAaY/bFJKCX
9RmZeRzBAq7bagHGpUA5YZJ4PbMR3Ol8zfqmcfMERvXupHZqM/5UKdopM6DA6E7m1aCucbnSJ0Cc
821tI4MKwoKvMXdQbtgzD1aSHOqvXtD4+41AQt1Jb/UVaHpT1pLXScW1pi1WnqAKM1ADuREAPpGD
dnJZArhYtELTNeBvB3LSmkL2mLq5Mz08yzy4fqkKre6w11w9mqwCsOI8y8tTlEUzo2fRUg72Zikk
6j5FViE8zwMk09ZIW34MGGDtuzM9Dom3L/0yIIjCccL7CB1mX/E5WufHP3Wi19RBLrYC4uvTx6Wj
U8UFDJMrlZlNJYyPGvFxvEQdnr/64JSLryA3nALl8jDXAq1ta/w0FwM7ll5AX1ykKaYlZCCAQESa
nhSJMr9iSKETm58T+BJEfkUXaZMQwNx+yCbyvvyRCpoQo78AzapRxZvq2Q0vFQKsh0GVO3cCsDDt
2T1gSB1mhe2dm6C36WE661k1p4rjIukp02cLDNWjqhJfq3Vu2YlqfITkdbPGOyRZP/xVMh1Fni2f
YZnD6Nss4Sp/moG5FcjSIMhU4nSw0VMvfYJsgwqY1qhg7Hx1UtHYb4eeMvDwcY0msGdf8/EHVPhh
vjuv3eLqpx7WqQ7IdDxRIyFQPHqHSyuSu7WrkiqBfCe86ON2jiMdAuKPaWt524wFG8lnPD0av4n5
ZIwS/JFc/hoEwWk9Ier6Y4ALM6fa88G9hL3EWz3RiW0YaDiOhd7qN1rZDEH7zMJurJJAwE1VgxtP
PXvGt+VAhQkx3rciOpNIk0HCajB5JvS+TMN6VA/0h7ghtosdAai+D9kieS40EFKx8OcBbiyOzT2S
5V2eIJ7j+7+YOTt/X95BYLI+PinQhnS/TJ2rsbI76xkjVe083ZPt406QUt2rJVKs4CxrhbeK+JY/
4ordk279Q2wf8xjZjeRiw7CGDCHG/IC2dRQIlmC0w8cZyror2s+JGUUmIkibKrGUT2ms79yFH6Xw
H63M4HddPcpNnEIVYf9kVPT4VpYnucchDrXilnEF0RQlm5E0SFv6iuvn7mooF2XU2agBSLOnHbwl
0+8hhzl90JwPXlxrWEIwwLuMbkUSf2VgZumasFMd5KFEqV3TuBiR8sczcjOf+ndLIvc3Al7nlH0p
Qwkh4RxJyfU6vsfb2inVOkpKkuBcZJ+3chEaRm1tQsRkQKAuaLkNg7JuwCZH/p5nv5OuLc7onaut
xBNrPh327rp6Q1W8HpnqLS1CgXt2hzWpjND07ErNFzK0Bm5QY8U90cWESePYYEK831++4Kd4Azo2
sVpqYrGM7OFN6RsFf/8Ht/696tpVvNbx2CXBuVpfduClXSXZTZJLQkeX0DtB2Nn2lfXkiR0fZj6B
VfoU94Hc6eXznG4uFSXgOL4jHnlM9U2krDRqY8HJQKyVolLjsC9VQIxRZS2VQjXs0OZaLAhsV35w
6oH7zH6EhyfuFZyNbVn7XpPmBrKZFIaVb1vSBpIk+jjMl77LbrMhBEegPbkwtzMR7kxMOCsrioxc
gpzwfDrQ15SEiSvCqFL0bPvEEIa+bvFugjSItkG+FYNZs2mxKT5mNwe4T++c/IjNaqCQQU7K+Wrp
iSuG8DUM4rVhd9xhLVvNUNv0tN8op+yGZTtp/eAUpsM9xY4pKYqh2caOjl1Vm6H0pcJSwdLgY1+1
xbs76DnJfSGy7ONXk604gKgyE8blIT6XHl+yJZpyt90HO+X2mp2vsdOFVXAGBPc40jIOzRRH/3g0
Kwe0Ugvd/YX/+tsCGovRSNPjH3Y1EaADc/3xZ5U14pNy4vl9rv/T7K0lAYNT5VXpjlULBUOHTqPA
pRVXIVWWsa1UeaOt3VOsVhmgbaghMKiufQ1gfkcNn/CUNFuq3Qa2538S/UumOU7awfZCHsRm4yqi
lM+OfFvmkgoa3W2GH+/4H604GQ06EOApyCC92bYxIX+2FhfHCddok7N40YhiLBetR946yuzrVNkZ
6YUABV2F7VFepM750tiXWeezzz6uvvfMeznVzYXbA8z6R98IQr2b4yhFhrfbQ7RwhOaIyQPxGUZX
UPgrCi1luFpyXjExJmR+vmRu5C1mb7pzEfhuh6v8QKAVoSawKT3aP8VWav01Jibo2z5EHXvZJeIV
2Ios4rOCwaqb15+mNxnrseDHPI6VtxhpmsTBvAoRGw9xyBqkUyBQwS2Wxo2jSfdd4FM8dXlqTqSc
f8btYTktKCPDlK2YI5zWMGNtjIirz2vhFPupOIWwiE5kAlZ0QHQSzm0b9fS4rEo5QrG8BPEoo3fE
B3DvtuzkB3Dz6UDKSnQP/TklePoksKX6q7JJxoPr7UeoZ4MM+qlk+KJNuvTD9We0hWnllrHsamJb
lmk/dWuj94Hf8ktGf9vzEY6AElWad2iAxMwdYK75SpAdJqjEwzDn9g3GWT7K3FUr5f6VyR0qmXW2
p6UnvwMWE3VasXdceYC7y9JOeLuQmM+J7RbVqMOoq9plt9L70JuYd19u+zeakvPArX9Qf4D1D56S
KX//+MZgwF36wQ4mEdz+IAnplmDn0CIHNMLnFT7qAdu7i9PATtZDH9QbL59GGH181gjS/YsrwdE5
MmwpqtZCKwA5kZTOne8TNSz35Sbl3TIbN1q1U+1s5RjTvSefYYiGgTlE/MiN5jboFauQNppLOGNI
OFSME4X8fdo4Xe0RrJEkKNb2N4eU0NziDelCKQ49VtcpLJoVtd9lEG2xqnczTBcFRGmzmTZDYuwU
AclMIiZMr5n3kl0JOXp5io1x4e3fSoiNRQtoIQg/Z8PbtfCeM9eS988DUkqlw1yTJkck2xTKBQft
pXfnL2FsjTE+ZFHIF2SrCn69USbIfcxdn9+iI+Dy5K2XUoc20Uj/hRw+lc/ugz5QrJ4tyngw9wOE
ueqzqBODCcBa905E2TeCgYEGFGXaKZ3NmNS3EEBf7ptkrHybmKreOZnIp4uTu8x1c5nHgABqmU0H
q9dW18rXQzse5HyYhp3DKgX9f/39o3jQnwsNmHUI1eZkDMbcT4RsGI8keo7EFi81oQbCysX4qiGw
Nc5H6bjD0lV3Tr2DmQ2niVietYicvlXPP+GuiNcZimo7F08s9VEXKBU0qXdvi0lh91WuEZgh27Ka
eVcg2SEHr2q3aKAEe/25gEbKw/HUXIJVgNccWB5cSV+mksNeF1T5v3By3MR/PNL3TcDo8HjetPzV
96rxxdHne+uufX74go7fGa5z6ZYu6RVGU5hI7H4wKpIxh4FgrDg2+EgEsK4lX37IiZ+0kRbCHn3p
VV8iIr0RrfLJUN0Xd4udlvzbB0f7xJ6p5NU9o8FXcbDhaZjjKruexWtGmqsKpeCQSDQwhDIY4zol
Ep36uDhncTzAETLKuXPwLcWGWh5HJDlC5FRKWkZo4jACb2uqLKs6UKG2wpkJyAsrV6ImquY+2LbL
bxUO9d/q/CAbSRX1XCUj71D3vNKkpWFM8UvpIXzoM46NbwQD+UKTvPC7VLJ//6TIexSwyneZ57Bz
FugKzXzNTcRO7lSwYUSyUqIk1x0ACoXJpA3XjLbyuyrmi+7q/DUP9aUsqx9YTCFOphYgYHjOdjEP
T3l6MT9b7eKEmYOzX1Hse2cex6xK6u6xTZf/7g/LEqD78xma/CyEZ51QXV1N6GxFdp4sFRl5Aq6z
W3XDnwPngG2vjVgwTNrLADididtqJQoHgawPX7Pq5DXdBrOMm3xFb6mcs+USWNbkQCqIpVC2hX+G
8qnBFWCSYNiItPfQNuyTHcNfMBCCSbay93RVnDOJNFCwkGeCqdEvXvCAY7eyihcCGs7VL4HvLy8G
8BM28z4z6bSfpnrKdxKr2tW2m1BM2HCgI1pTEVVkCXax16G6cgHIVUJazLnrjk3R2hFgZF8zeoZ6
2z+hz09lhvO8H4xsU3Xq/yIp41X0VdJd3N6etq9CfyepmFGAJphDoUR0gE6yRtQlzxUKuNOL+EMC
hr3KdR822DtBxHHEsaxjJc5Sx0adjHj1Zc5E/tjOJTkgr26sFNLkK/EiBurD2HvyKu9Ct223U7GN
Ty6o1H0HCy9joKMsf98Kls+dPnpcB5d7dQ5vrTlF+zgCS7WH6CWW8d9OpsDZtXvDQTF2a3qumVV6
NF6eilUzA0W/D7Wg9U8bZYTUfc5JutoHQDcbiRRWJ9b1NhABPwwycg3VhSugtL/IkA3KL5qshG+1
EG/nUBjjJ6L/nG8N7IBgj5iclQ5kDoYWtpHt4b5l3AJ4pbbIydA2D7YgpzXOn6yCGjO6wQQ03w+k
WI2JcvrAisTski1c5ESGfHrYqpJv3fbuQsJhFGrzlsRownyw8xN46g7UizTr+C9jDw+ZdNVhm6Ua
A4UMxuO6BahOeNvsGABBqEDRck+0yzjoyFAq4WJS8J2b96PsentulclWWacQfDakj9etCUBaffzx
JtzSgd1jrApWckUGdUSBKulnXj3TvUKfkj21B2CF0cEou6rebxUDOJbivumqCmfD6UT5ViSg5APH
G5RZUBxAHo7P/z5ouN38/TatCj74ZhfOYHgAVjU04TZKbBRAQ0A5g6BYIq2nyOAiLJs+hIJuSUNo
59or493q+DeZTtanMe2kagfhLK6aeYfeKfev4DiRFWW837viuPPhpgbUjrPoVoLpmctX6Y4jmlc2
8Jl25mEBA5jgb0XRIsDIqwZUwASHR5mV63PUIpxfx1qY0YI154xlSZPdR8/y2++X9Pisd5f/xgJp
sAotPmXNIG0PjzAtyyA84Fj8ZhedJ/V5ScepFFeauaeezavL8KFroNsoIwpKeUdR9YQOVbX186mk
MjBngUDEFSE/RJeoBjQAMRg5C26+dP7/t9Ont0HwSzx81JGmDQJ13ZIG1XIYABUOUXiwkTcXH7SK
HNfuaAEDZdnT25f2pWUUupdEyVrYFRVNYOEia6ViqN2aDDuVB6oKep18EOLOUdNw2MA3N8h1G87X
X+SiUmG3iH509/YTwZdMROrMqHhziy+kBiD6mGde5NIuqi4SH46Tn75rNGovXbXBCFBgw1ro236P
86soriFN7mfsfv2TDoz7eKhEKd33UESIlkC7QqS0No59WHK7/xr8gdhZBahq8eEZpjz/xrh2r86x
GH1WBAeXuLyrgs/P7U8zc4LoJFKAgOsATJlBIwN3Xmadg0mu/wBSfH1e8A9DpGGdU5tBCx5Vq+kW
vFsQS6rjYRXUID3rs8RfmUCbZ35CKMH9q2Cd4FX4GIqnWvYOr/S4L8ONeYWzFvZNfH9WCzgwmpZw
Bf3xsfWMCWzlCJ9b+QDGoms0xlHu3h21d2QmzFoxKLthy4XuMpf2PsfWmNnGNQCt44Hzl6UesH/M
Z1Z6kfOm5AqKtoK+QDklBJs6q/ArNzhyKxAv33ojCqYVcOA3APSITKpPx2GFOuTWPaHgsOM674/o
1Vo4ShOC0iEzmE27Q9RoL7WrxCcKskh2+znc+/4hEosqNRcM3CqLRZIeL4oovOcKMTqcOnKDl761
Yayl04rjA49A8V2nzWr02/DbXsJ+ES0Eqhsc8iaqaQNCqDxptG95UowB2PdpsAZ0L9KjSCNy+axs
S886Bqm0cwDYZjrXA1U38y9z/Wyu7YDlToUWfvompArHs6PZc2h975/bAFL+5gygp7/z1ibvPrYH
LkM9xn8ZXRwVSaU/jBZR1cMenZlpLT/IOoLPo8vbMXXI1hlDaZTr6dBiUZVkn99/P1zBWWRtwdRO
LEtsMAl4JQjSHbZL9jp0ymJRSKzKMt9KgQel6kiSAq0+gSXNv529d8PARWtOy1Tg+3KrjDoTJEqS
oH4V9XQzZ2IaHH2j3N2i22Y8q1rLhW6olrmu6mUBebE0KOkgbMG9XL3sYP8PH4RawzdY9bYsQ3/X
r6Rv+va/jYfU2WZgN/fSux0DcFjRcNetGu2XwD6Y4W2tM9qiRU2rrRRFOVRea1vr2yvBo/K8PppT
N3QBsSrMnyuMShB+qwIpcAN5LEmlOcf4/os5cOq5JsSTMb6UJVo5VAilgNdlV82HaeNrGbhTusBj
FFLPn1zCA0Fa3+bx1Fip6QJaiXKdoBaLyajJ4iBBKdNi2kBWfCxZEDKoLLQY1HbyLgOk1RWhblSV
QqofITF0dk0EdMxwT6C2mpHg7DKQDcySh2U0hYyOZ8HVuTItzywRS6GS2x7a131n/ASWmhi37MFQ
Pnyhagm0dSIBvl7r6bE44cLiI9l0/yMfZ2pc9TU7ysnKumGBwOjN0bx4yg9UweuE5HAQXdyV66At
4OPxElxZmKV2YeV62OyCzLGPZpZ58MQhzKPl+leuz6oy82kifM/De0CzZdhAfjHbPfpUchh+K6Eo
gxK22M/46CKpq27oUeCxEjpHP01UCx0zmhBDWAlPGyID6UVsgoY9zBjL1QPxMfIPBHEgyJRB+wDK
3u5JdjcTpp2fym1ZqHVCZEBZlmHQP8QsK5qNmMLfu3PvO1B/Ha6ORIs8qbSMvEcU9Oyf1e1nEx6M
5qV1oyWGnhTzyUIi9RdUOLEHrqruZeoIqIJUR7JxwQWdjJsZ5Hpt2BGXgDOXswgDTciYgu4Pv8GO
1KF06mh7QPRlef4XjdWWCXczcJoaPpHt+vhq0pPUXUkw6tPXG6w2KvAjklrXTYcaG9SNDe97/G4w
LlU4ul8kw0VnD/K9IdNXN/ndUt9A8+fKTC7XE+ajsNJesWBHfNGaEgdiudqKGXLwoqgdtM3sJZxR
5ZMie/KekQvfcPACcaPm8x7eVjJD8TWjUTN5oqTRQhuWydWiNCoNWKdNkybzbtqUQCszgRm/IsC0
Get2RvGo3zT9VF9oq8NZ9bm1zSE4rLYZUOd5RI4RDlJHNXhRktcgQvKax3RbxJ5XD+UNbaTRWttA
zFTaV9X1aFOvSwPf4jPLRDh9XgryWYXyVOX4vJLRuwZGlTZsetxlmsqHU40evtCOk1nbIJL9J+U4
m3HLST9JIp0sSIDI4ypAhRhfVHpi8CFjS4c7xXMRoufRtqo5sXsvTPj0PCrWBuNe1er+1ZwEieLd
1On6+J+W2EUA47mYax2JRBDri0DZX+T0ov68+ONBizhtssAOSLfvixBI0StAwKXZZpq6TOG4Ukjy
QH4vKCa11xU658R6b/TTzVLnp+JXmqwsxwIij6xEvxMsdMaMr9EX31MmHBlLtq1wC9xIsz1NrOOv
a9NZcOmrmMEU9O+qkECh3rtdbm+ELXJ5LlDG9sXaKCISXRCBHYbN63CO1M5jdkX+m2u3Pz7rChfQ
nGFxNpcd9QbN+8WugBZd21lQwEdQlLmr7QndEwXMBgoo1Z+QQu8QgvtC7DjSnc4SE0QEinVK93Po
bm00dDKpNhcQkm2Q/d3m/dhxhuVrj2lk+TKWnZjbtRJ4fJj/2ytATBZTvh/9yo7N+j5dkXL/CHq7
s1m5MBP9TyYOupsfB4HteS7QEzhRw/aIyCX7//Db/oBM00yuhXVRmmbZPsuBE0ho7POwlHS41gWP
gAbXK2XmJUTOLLdVa0980Jxq9lMPXcNX6IedpcWzIDZWV9SgAvmSsbbSrURYUNvZ2MEEeOXtKB4i
/uUnIH7vxSX7Jjmz2Fg38qjfZ4PyGp4UNxDSHiNj1UXBO7+16T6KRHrmnLwLkhWCAE9AVAn8UgT3
xokmQxtVv+8F26oKldOG7eaBe6StWzQFt5AqitPbzHCz1FoMr8KgDdNGcThvE9LyKJT8xaZni2ON
/0klFxtRZe7A4Q1xsudGKit4eYkJHXFH0NQZU2+ZRnNCSUvtMLk161p2vOxQx0SKaZWSG4MF6l7q
DrEk0wunTbdlNbpQ7dPnUqJVW63w0SUoikO8rjjw9ux3JBvlK/48JqGQmHiZdiZ0lklOltv0VDdq
olpu67N0vi+6WuEX77Sc7U5Q2dFDsuo048BSX30vAoza1xEu/JdzYGx3UypTSZHInUDFZeq3XTYf
r41kd+TUOZhWiQqkn5oERNG0VT+iVluC//bSZWF764ejGysDxmH7kNiyVaFR4p65OSI/UUoekBtw
F/31y2N2FekauMgKIabd+3ss+M9DWUHWERN2aZYeBHfMBpeKaKsDaaKRBQE5UbObsj1JS8cfYlce
bJ/mccr4q2A2PhT1+e2KgO0KJBiWvIpjG7vFLaLiHC9XlZyjkAx+Ew4MX5pNqE43X47WSBSws0D0
nifg2ouomgPkPXPzCTkDw1x7KMEA7Wys9NxLl9/WbLkScCYvnqk0YUNX6wbnk6aTGnLBiqriuIni
SMHNHB1R1a+r2GL2NyY0vAi2GWqBp749mXUBP7KLuTBLQo42HDJIIdXwSZrq+BWSx2hXgFx9hy3B
lPC0EQR7dVyumdtx9M/3Fyf4xONLKNX+PKIKiqnYzGTnMjB6yiUBUFWAAV9sUu03oHK/otJjaWIg
sEk6Pq6pJwl8i7en4ZB67Uq3W+7LhJmlNis7abWlwzG0LSkMZsLG7VTKwt2/rSc1uYu5IVkYGBn3
PVSzJuJ2jCKV8euh6J/CaCS1IjTFlRgXqdHvyfIdoP6sXEZ/Zt2sEko3Cy100MRTRGQ7t+mAW82C
KHNuIWj5LEt7hPjvm4MAbTJZocBACW9YcGqNGf04eL1VIebhlALfCkp2HqV0bREKhVho1/yZc6qU
SY+V8Sd19vUemk0ZDZzZo3CbwHXCk6vKDkACyZFe9QQXtvrIsVZpR5MJ4JaY1wLkTwtC+RfMiyCQ
FGAzHx8+FRcR9rjSOwY5CZkQpyvlp9h4NE4bEFEjbEHMUA+eHpE2UEGAxuk30v1g/xBvGHqa9rv8
IxwigNA6ZSdrOix8bTQIyqDa/pX2Ce51BeoXVy8B6YLZ40rEIvd9/TIu5VVLp+fvv50WGNlEGe+U
CZhZyx/UKFr2nNBKGr+K+E417F5vESF+pmwOvK+z+huHgLXd3tfxNUUn0DLI8nkHAq66SZ5G6Lqm
AsCenAZh2EF6Cbhp4inM0pCJPACC3b+hu4lM3qG4mVfK7EBxP4kCjGGFz/k2tbHGcPGg3ROKq9D6
JlGHCsG899NdCsbhjB7ijxESsR2I1cm4R1bKJ6FrIrPKn9ZgX97DiMKpQztSs48ax10co+FlqzvF
edb4Wz+aXUAVr62duy79s7Rf/xvgokDsWk9Jfn1M1xhGa2VRQdNfTbKx/dyA+EPo7fe4J9EBUUoL
2YrrIfTXlobn9cMwDBGY6TzbBhTyRTcmLQmih1NraLX4DyHf+YkS151m1tQh76ehkt4NOncIpd8Z
pLd9IubuVMJVi3cVe+a/0tiDF1vmMm0YuE6Lnpwt+YvdsJa6TE1k/LFwixpFChtQPm0gEmeh2teg
SPb8HGmHzmLvfPGBHR/UOeQ0FWlsWjHFIBVLUEQ33hSf2cXWACiTH6bbfQVDIohQLkRhow/y7Mwa
mEFYEtAM+zwPYJaBwztzD87zedDz99qtzVc2kd7Zf5mpj+cGN4QSmE3PYZAapZKBIpdI3KigT8/v
NG2EfgVHhgYmUryidcAMS9ceR4ohnbMOsK4qwW84XWKMCyWANIMO/tzWbHzxg2di7al8/7uSRty6
l9RrEjin9aQ2QoIXU2lIKtP1dzI8lgUqKrEiJLh171Rr18QZqTXeJDG9Gctf54/53/0ZDUklwBWB
fPY8qg74T25jZWegTUBUDZG6xsRGokidfhtJv1Wjhpb99ixB5DMz4kciURnHQL6AcbwX+u0L4vjc
bkHIjXhDGSm20exeUq5pQ8oxb3shTXbbqO5Fh9VZxVENJ+5i5hy2UOR9x5FN9RA8qsHqQuhEPFdN
bhImdx+Id+0B9tE3/gpU2dSZhVMjcCEVD8zFaiA+IXrxSUkKZ4v09/wRnsF0qyIO8sTPOG5h+ObB
M0bai5GfNgHptB/1X2IXbCyFuprK/YebRJ0vDo1hSRHzsLFWC4r8H8jHnZ96oLxq852qGiBCpBrX
XavvCHrBkB+3BD6EmW9oFULNZsp5uBvWP4Equf8I47LuBaY+YIMTMsse7H/1g29/h5wkDvcqfxQ4
5AyF4b6Ow3qBHXdTNBYG5BE4Ol5nR401WgBkK59KT5tLC4vtmv3QxtzBj/rmeUFIcgzylqVe9LT9
lhXf1WfO6BdXYzIlebZc96ZTrF6tVGdwwm6s26IByX/RLvPlJx10nQuMkpolAfu+YhFQbF8ut/Bp
8YlHriSkef9W13BAEbLW4k43k3a+TMn3ZKWV2/zVqDRafeie+W6OP4FkhbZJmWAUZiptL6hm4Nx7
GmbL3aLAC92UUIOx1OQLQQsVmmYK82TePTxGYSuaPTZvTZs8KVM6YicD8WcW4e1giA+vP0f1O7a8
16D6FFoaWuc3HLlic8XMA5aYth6eLsqSYMq0wn1060FeMxBYFzatZrxPTlQPHMoSwrwW/dXMVZ6r
95b2HVdM/XCnUdtoPTmZtjXq/AXe7Zgn+2Tgg3QNBSVw68+l3sQIEEqQR6lXaaPd1CNtgG0df/3w
3m6fi1w0zHKN7OvvnWELZC/WyXOALL6mkd0Vd5NmNtf99l94S6GG+rS34eg5ML0JLX3JDvo3rhxL
0DBBRLVArK0rL7j2/UUqhcp8QoYHovQM5DsJTUuSgfLt42Hif6EmxYJKiEk2W4ZBMjBI5ILOQ4qu
Ygv6/7xrHJ8GASGc+Rb71ize7h/A2J9S7ij2xNF38M+q7soCIO7hk0J07+31ztB3TvgNSpU/UE86
+4Bh969iAVvi51iGGHBASHdgVQ4edPCiV8AwYBSBfNI6f9wVZi2KzY9WLiSNZ0D8cehaEoB47nZw
OI/Yon9oG27umahYVt2YOp77V6HqUBCtb5aUfB3ipgX4LKifweaO7pz7XV4P71zgwew9kuufVDK7
3izwMYCE2M0rhkYQHsklMTjlBXrBH0Apf2L0BtVaJPPqPcBEkJ3DOy/QYGlLl9dT9LXirjWq30n6
OcnXSaJ0Eeumw0lQ5utapb1VD3CyBHmJgmR1ynk44RL1j3yeBqmYwM4cYmCHJRDICZ3jjSNXdrq5
VTMumZuRcrOve2Udz9aqFQQ7omJ3HL9+M1JwWEBO+QqGlnats6ZqzBv/aATRi9GgeYWFcYahMyuO
rD8hfQbn8pd7JCmAfVTwzDimNlvE0KQ/KMUfRkLAs6Wd6yhcRYdxoZaxcfoar0xv4ZJlphQpO2Pd
Q2r4PjM7QT59oNeWySSZ7rAp3znYIxJLd6GULxgHue1+rQNGrC3TmrZLV1xQhjMzBZY8xcjoA+ul
+fX4Er8x6MiJ0tOWM/6M+C4aNnLeSKWtA/dp6OazLrl89mZ1ihXWkT4BdlrGGOpiTf3vg8dmGiwp
v7ToVQD/buWUYPjRODleras9D8SGVoUhGcYhDEc7gMRtJ8kkOe5ea30rStSmN3fFyXCiazqUr3ec
+W/jh1kF1F2QV7c9DUHV9Ily1kUfgfsp2I1V8J9F3iomjE2406ZvFXX12ZfPA/ikEMEdf+KvD+Ac
3oRQfAAIve+gokZe2RC3hthV90tJLrJJWGWE4QmcMat6Ko9kqLde5czaAEbTHbqEO750XrDjO0EG
SnRfMWyAQpTAeiYp5I6prGrCKfSoVv7MG8hZwxwWQ0S7VWaRcypZe6R+vm8sIUhccB4DrU8LqS9M
l5LF6McjmEIHWhKLmny9F5s7I2MMsQQWA+FpAZUBZjRiHS5zXfSjKR8C6rQ75TmWKr3XRNRiJrvT
7Ysed38WcevlYrgAWZl4ctfghvbI7jS6nDnC3RKXvxzbLzDCVmGbfsueOk/sPDUkHViF4vxdek+I
7WrN4MuKKoeksY/fEikkzBp/XNeuAPvBFfLIlo0AN7W7w3aNs6AcktS71ofuTNcOKyw7nOnbXyvQ
UeeBXDBDerDfli/EqX6MZvzl5mySsSjTAQNJ/1lq57v7TWbfRkWWmIJQOMXYDHqzXsp1jl2C/4C8
w11p4GDBEvPOPnd96fPpSTykYAPMg0dCcb+qzPCnGQaaCgppZLJrh75TmB5hqQvW5aCShgMTzQny
s5J62jY8B4iwLznmHDwbtBA3kMQriZ5Nsfv32XY6BWEJchcNzgQfMCOL5RkqQ0dmnNt5dupgBVU9
ruYESqCKoo+8MLGbYe8N2ya0P5CAWgSLMUV2v3em1CSLzA1Xy4B5DFjD4l7txIaSObdhYKHHy8An
nISj8HOm5xtk6eLndp4WDaGqnmEd+fPirXIbNwlgpV2lNoS9fnx+8rtM5ZmQFI/kpsHLpHeR6D47
Fky6+aCUuKHTLjXbSW2FtFgJtD9gscrDcY/fwYaYtOQaUWZvQH9OjUXxBdb0ftH1yA0zizcv9giP
WCYOUidWPftDM7tuExniX18q4V8zOuq+uiqs3H6cNoQL5K9Sjg/8qCZWb3p6+jBwBTZ1+tOJ/CEJ
mMJL3yUcxy9hNQJzqGxbjUFOYcuuRgSoPgmQb6r7gYzYNzQ2stg3FV0pT6W7+et/VTAV1Mje/td7
E8cFD/vwZx6LUd1g6sM8XfJUTiz7U+SdewqhyKnIhTFraquwZdnigj/jUaiwb5KGxR0jd80ntFkH
bEd7RN3+P66cLKv2Tc0iA6slYIJlwo1fHxiGXy8hBUQoyXef3UEDG/eE46WYgMUkXBt9u4ZqAkf8
Htd9pdt75HUmM/8yBsKAqh1s2cT5IRRhWb1Op1HRxbhZ/StDBKnYwzjWjhKmDT7ca8pT5b1vazf7
0dKrmXEBjg6cz2pwVQLrnZCLvpZ1ZFntKKVrLxKeLak87lqi5pC1GpTbD8DCqF+JOy149hvL7iEV
dTcNZwbzCCBOQ6MAc1iJve2kdMTG6+GrssxtJm2NDEm3xPW4tK+ZPnS5pQjEfUvK53dQw/DBKV0w
io62t0O8pihja1uCDyKetu1hEqB96eRTySp6bNb79IsRMrw59hIHYT0INT/1x0mEmg85sVwNAqXo
l2aIGLV6hwloyxB/GOh03ODHy9q/Y7QtIrKkxVLzRDDvedv2VywXuiEiCBTGUG2vkZdMP3yoZbGh
1kcz4tqBtjWhiAn/GIMVSPi9KmNTMznp461e+zSbUx0wYhP99jv0EZGCc86PjBzNGW/kJeYVvW3H
ZidUPDJXvZ3txRZFAoc2x1ByoRVdeuRk81PzZjm5sk9kZuiRrBexREyaTWvJkz414Kyr8fdIpqOU
1P+UAeIumIsL2uAlWFsJTvERkAIrGfhnujPznopywxWnbrz0epkwdNKRF1+d9SgpJFyXy4Nl3JUw
Usq0Wlv5NuB1vtdYU89EPm3E1OhSOH1uMrlAGo20cUAzOaqDUa9JQ+eWDoAXAMzZFepWw7jxc5Xi
VzKgqlstuzwleYW5Ud4q6CBl2aSCNrVt9xD30WcA6+U1OPwCaSh69yT/Cj/6t0/Ops8gWa8BwMFZ
uRm9bJ/gdZre+PwYqsl6IHXSefJNPDehws5Ra0v7/CRbSxhAZ3xk5npY1kJjlMKYSKC5iPuF5g+5
MTXmkPUktslcS06dLZSPofI+i1rtiR+oJrEh1cLhk1NBQdHgwt2xY1Zv4OaQ9qQTSzwpgpduI+5o
D0TiQN2bXQ/GSxhPML41SwMj+lWRu8itiTo1fB2HgVX2AtOmQFy/6flBFEqN04eggvRKQH95KM4V
ziJGYCXCaO/U7zkJKbGsJujymNvhCH1ztrEyFfkTO2DJq2c0U00e3ET9zg9CW16wX53naXdTqX1+
77VVjgSt9gFNZKu860Rd8SlwP9Lqs2vaYspthQRstnEPmEYDw8jQ7qPZB8R1tMHp+jreNriXV4gg
rrlXjVa92ibfp3kt+9hr1v9SmGAOGcecvIkgGY9hf0McMWpYrMUspkvxCwLvzbki+jrBocWl+flh
lNTsC4EIJ1Rei27QRJ6LQhKrOPHBVHyVReP13Do3Vl7yrCzxk58mOOm99A8Go+miYbKh0PFiaznQ
HBjWkXO5B324NrmCX2NHP+dUPJmTWRP8TXUPAvoRbJQNrHJTcnaVKtvKC+OmHC0fhH5956lHA1rT
VC6OmPi7jSYlTTCDbJRe9Trnpfis7fkT4iS80gMXvdp3nYMl0tA0Gwww/Gwn9MEea16IRUV8hf9R
bVoYKf2X51EHFmrYYR4xpAVAiUvwCZY4jENoeuQkrayd1x1DggBNWnooS7kZugCgwCKMHMpFD7PW
rD061MXyV6zOL5YT5IWIq9Ohmn87v2LUcp8W3d0X+709tqbUE43y1D5eG5drhXmGxN2opJeHti3T
1boaa9A7RbkR3u178IeQkmMJA8t0pNprc6RL/V1o6TqFNGVB2jW0tSu+e2u3cbW4ITzCRXhDVC+s
SLiHcxZa1rJKAHg1SbBmoPbOgF13xA37PVSLsmOTksEhPp1QjjNYvzLzmniuiXE77gdNdt9RCmh/
PQEnzqBHjJONeDiVVApH6Wyk7OB2dGGpThmAnjLJEIDUT4gqE53EgJkGG/LCRPktyyrXrrrz2JP7
Lhy2dUgUZd5qJWrukbYPskgYYNZToDI24lLfHWYcpY9UC8l7DsTP/aknB7RHxZMWz8c7qW57CWbm
R8Lhub71C26MKl0AGz/lXRWj1s3ziXk/b2QeeSBTErzvlxIQvlr/O8EhblQzbCbAiTf7DNwJ/ukH
26u99leGuTeZSHPYt9PVPu4Rkf1Rsoi9/efYJMN1UY4cBaAxfF0rVVFOdKqsqtA7V77V23eyml/q
wsqyGIw9tJYkvt7FFHEUwFqADrKLnVAXqXH1S5/QsZfNGWkkvjm5TOv++rbMnHjAIYArLHfDGeFF
720xsP3N6008l67qds0J4hUFS8sU048oDPbL9+avsBWaXLlk/QI/bOvEhafHarqJB7LACmhgTs28
G9K6E0QctH8xPMebECOms+VWGM7GBLRHtcNmLAUO6eHE63yUnx3J0eHBTYfTHyZbKhWdZkZF8Fdt
fqZCOF0klbGzhHSITdkPhlMeM8MRWjMPSeV46V7zyQBFiwXBTddQ2AdhofI3ssin9oAucKK4lnrG
JBu61f3r+42EDBYiDE0evyDijm6Lc1fXz1RHPd4nRv56m0l4TpsNgVGiLtiSPT2LyHGPK6cY1aQZ
0uHMYbgMts0sBGRXSFHo0253rVk+6e6dr3f7zUxW6mh1xDoWpSc0uyjTZJgWwoeaNXFHgvd6B3uQ
xxUJDlUR3Nc5hiX+XIwCim8NgsLdN+l9zoLx7jl+u8bB5aJO2qGxY+gBJfmvZ4Rs0msK1Yq7gKEx
E7ePpi/60/ozHYleY1PtqlwbwxQBO/d1iuTh7JNIUjimIBKLJYZGNClGQoMHL3xkf2u5rGvmP3XU
7wX4SJKkuPoxRnGyahbERCVV8MypPtjuawepnS9k57jyi7uj39LjkrI85gLmSSEwCh572bfDBO0Q
4hmNa/J4emJlqtYo3OfB8RinB3pytFUubswNv7DaLv0QB2QKfD2cl3hQ1wDCPoZuHZi0HpQUWQWJ
N+eY112Mf3uuSfhYQ/XOG5Uoj11317a8mA9BvTQTIiyYu4sLHclfir7fu/y5Wrf/iR3LWJXHJJ11
+zgRak+S5NlE4J3BHf6uu5AOksroKHfgWK29wEVuomp+lN4ZXMt/+gCvwYjfHN2Exl5FgxeHg9gv
BOYkLEf7V+rbjWKBA2aJxVGGdo3WJ/D01Ajr2MXpHKfJvh7FhK74l/OrRyGSrrf++GfEKROrFoUi
gcrARAdP25t3V89IT5pKno+vHnie9xeM1iia8PgLB5ThZdMImRZqydoV9diRt71nyXRkGJMT39od
8Jv1eEbzh5cxm6c41cfpXOixFC2uD1QEXEBcAgBvNtIpGqNGCQ2vxqsC3wBfreFAUrYDCWyF66ub
7uxp7O3dVOUXhJJWntu/xn1JjCmKD/jEKe0m+UC2GaSV+Xwb7Lg1PRHv4m2r3Qb5W3ghu3hlxup3
T56quD24Ztmth+SEPJMili+iEI//E4WC0AZUD6TrflcwkElSNyqyfcwOE73nEn9Jz3o46RVD8dG5
QO+fnkv2rDEpeTrEVbDi9dWbXBiayiWpUA6+74B0XMy8+LDZA2OQ1vEcquHoa5qA1w1tN9scxiFT
hZ912oZmYBXq/s19Bp/ZYPXMBTH80i+s8wuSdtuTLIAoVG5l7zAhJcVgbFhSM7z5YzCNWXoCaI3m
nQZrj6bEV1R8ooGOgoZYOUHjZbdXBqNhqXTOZQE3UEIbMiUqIvDATii4rDiMSjL05nTvq8bdUXEU
9p0yIXftUjhPpG7sZiAck6J5YVpSXCWwml7JZKRUznPb5+GV44x9wBJoC1ceu0o6y6wf2MkYyCO2
cLK1uhDj/QsFWGDcawq1vmPuB0N8liuTg2zvNTABab+W5a9R3KGdhFZOk+neOZpYTuSN/qcBokau
uJLuTwjTRREeMcmb2o2REVZFnVbrprCLQWg+W8UZFH9LsOBkab5AFJtWcJ45S7sSEjJi5ISalqcO
F2mfgMYcyo0Z6thCAAuCeRuthuAkqzWLIGaMVvZE22ArFi3lOlWR9fgM9LZO5j+v6i3wC+X87Y1o
Gp5lAJQ/Pi6ncjsla0K6URQta3DpFyntQMy37lSYdGY2vFpEg5VWF7jPPDQ9x+pzCVQ3nJq7zMAa
SHzI0383BrTWlZqTPk9JAjmXc0qIdc76Qop9CyTxw7gPdLjcjt7ull4lU/8t69+awAUaQtBT5Tzd
fGHk6BkrtmqtWHoPlHV0Ai1HwxHQUdbtUDAO/f1FZS9ZgDl2Sp0/ehi840waQhAfFHb/BvY9tlFQ
jOHoXt8f5wO6xAX1p3jaW1dfThuRTRlZwvuNEZlEDEkBWCJnJAJC+zeWNy2lR73rleO36rFZFBFy
NcAyfd6Nkvpts/A3eV38rKx3nXorHCjsAf+GqyUgCMgXVu8K0GYefwK5vzUmwh3GkCvnCd5tXIC+
UZzzd9/OAHCA8mylIrBGg63CXtdKJpVOzyFYjIkJsgWG/tuwlmZka99Xf6RwYU6e4UZaGmBWSJzk
FH9qJZb17Z7OVwwNmfdt5SkvNWXcI/LEruu/WsRqYJbnk077ijZhlCUBokyip2iPJJny0I7shveC
AUeyBC3gDnhkSkajdzZkZSjG8ZjT5Q+NTCpJDbwExSMLvUx9a6UVj9phaxSQ8AFf8i0OhEQtPomj
eRRHdrdZlEXHy3mlJxN0boRk8makLkHHty5xhX7/mJHBbUYavTshM32gl3iz29iW8E+YazOu9CTb
md+QtC5H88PhGtdA/4JmyLScf54OMJG1jwK7HOV9wv8iZXz5EJUOtBrLm1sSRx31oxP/58KZaspw
yuPWnBGexiDAyRoOVHg06XglE4kbOQN15Zm8+4Y5R4B/674kied564Bk3gGiA7DBPFI6jY3O3Byc
G+EeOPDOY+LmBHrU5Q/9st+YSzRhdhWAuz2uvFH8tb51aiyx9IvT1erQJvh3pCFJTLpMtGIM42h9
1G+6A5Itl5ng+OukNZyybjrDZK7R736j3U0uGe47QbwdkgjgvWtqAUlnbwdd8rrSjE4Sq7eTnJ3q
zOlFmUEY2ZQfsJiVO5b+UkVOheaNqFWEcnaSGGdRXWBJK0DIPJZ0r7KFJNIvWRkCOqR4969olka+
0WSUbQQEFL7S3MeOMVmspfrPJ6kuWNCqMCGniUI0nv/9e0LlmfUvJptRFdHgoks4FTFsmc7B5y3R
2yfpUHGQ9DyVFrc52xX3D2OxZQIcHDzqwgAdNpEjQTEvOfjnltVm/oG2yiGUrjbAMLZUmRP2iXjU
8RU5oBaSiiEyVHU51V+vy1sv8foaPhkUbG68+ioKxYZKxh7tvyCwOJHUqc5sSvJYPw4SOG4IGq3t
22rsrAIUULj4zhTNHk52BvDPDShM3sgilLOd31xWspkngti/3kUitFHTbnQYs2QW1C+SrJBXTCfi
7WIjptyrHK/bkbyYY9x7ARGWZnlOUlcH/jbQJafB+10KTIGAmIWIvcYhom2Auq5FXYFUUktIozC6
LWlG3h2HplwNouuGYV7eSKb6tWGU3xbu5ePxiS6+eGnB5MvP7vhK0m+Z6zqqyCksUAq2nm6a+YFt
HUjc5MhCiucADpMSar3DKlPv6fGc3cHWSqrswIdZ5Aa8nvx3eim3WS6/5m2CvMcvWuSytq+FMvWs
gUMVQi026P6x9CNVyPqvpZpuFmKcrTZVBQ6rNFVff4bntPXC//e+DaNT1s9mQl+nxS+5sgDuA1w9
ZLFeeBfNNY8wz8KdtlUdplovRlPqomXbwUY+VXC1QlMmKdCKZFUtIOmQApS1WSp/gZxYgfUdqUbM
Jl3rUmlQc1N9dlasY/bYJfKNLG4xHF7i0pLwvPTL0mfaF8RV2rMM1jgRLaFET17sAPKIJFwu5IhR
yPpgSuoxbS73vWU3W7Mo4zZuBzmWVUMB17WclzDJmsPcgUNa7JgGtB1cOgxDR1CZnxI4+vn5Mr8c
pL4PsFxsmZ1RLZqulNZg6qqs5TvmvZjLMS2MCTiRbx5tV2Y245RLntpF0bikKqU1ej4exy/7rAQr
IC3VvuMNbSgXSZbMgBZQqG6nbT8NffvvI+447pytYwyXXOzEvF74nMOASn4BN+5gO8FuE4BpSDVb
ldxAveNfZYJBWYM+coJEdfTaIJM+knVYtwogK3l6V4Jbad4RdmjOpWcEIbfUOtY+EaE7FWvqdLHW
RRa7ffJsjuf2b6bwve4Q0C40odSyhgRF4i8TSFdHgFARq9yumlkXaFDWy48VYqz9Ckv8sDue5l4g
63zpetsSZ9hFuE8nvvrehkgHgWizi3/vSstTw1P49reUta7HtiU0dEamkJqbrCYkCEoSOdgXJ/nG
FuqL/DPYQ/O9Hb9d76CxLCaRD/RtnErMVrbTK+PehQJ5HZ6VJDudgTd9bGyWpQMlkq5rhFnYX2mE
x897do/fY3zShgkYPF/eBfJXUL7ivTBsLCcRVHZDXtZ2f2jSUBSCJ5lqSqiv+xnqAtC8RgTFyfR5
iZG4XL8/4xe6n71MfhPB/TczIcNereafaYyvXlvLjTWQiWPQ4HXxpwBSO+pTOX5BDfVgneJ3Nduf
/rnlX9ce31GmYSfkxrbMC308Rjj+1ggts6GkePuo8g2DQhynIn3SE9YPFbIy6q/cfEVxEhPGuN6+
8vxuUVUhkGT7C/152aipxQe3j+WRydjiLrKuBxuhCcKDTRHjpDLfT+9BBxbwqdcK68VjdtUJZCOw
kiRo0H/LchLefinU5VlThpyuwbGMvyRbRQ39Lm04UFUnZbssSICSUAVyuUivt5qD7OT6TFpCjtH4
Ldlmdfr5LBAsUIqMGIwJIrygoRCXJXlMHkB4uUAwcxb4Ri1Obq0QCmY8w97l6pvofWuvWV62lC/0
BJf40llHuBax3aJcOmt6L3hvP9pdM8zfpQstYupjpA9uCPuu6MNw8CKM4Q+Ga+zuQjOqkfn65lBx
GrNv+CRMixlZeEizRDF+nvgSr5aWNGCFuX6iy346jb4J6A52pQ2saKkHcMwO4oM5xn7e6fTXtRhk
Ihm8Fww2/FLZ/IBExhrOJzW47vXKPU75N2rK2jWSRCDYCGTjxdzwJHJQMSF1E96QclwgQ2bdPV/Q
McXL6M2+kCLxP8l243LY7dKmA/fht5Wf83MHTzmIXUQI1/rh2PrzNTDCq7Vob4+YQVjR4qQWz7e1
Zkji1WHIFAQPwu61kJHy7BAedVrlQw6xwLI0vZtpn8REjhRkjGPfExxR9naM0Iy7SCK2Xj6Q35WN
xPDl7vyOZq92ItZgQtLe+8CAzIAK0twSnGL4nT+lXpsRZn+SGaFSj+S38ZT/h2ByaY6PKC8Y5PO3
kceBjnsnw16Dvc4knKPjcB5zP+MFUURp0TC1+TocEXgDz9DTvDfcFY5/PIl4LzHRWKZzVjZ2o8r6
kOjmk+bdhm7FV8JIOJhQBE+Q6q7pfWeenbdAWw/mwNxan8CYYJ6vhfUpYty2TdtTVFjeiiEDR0rl
/j6RFhb2uKltedL4vPaj5FgU9qVIK+yFjqLgbzLlCBoD5/rldUl02+ZVpMS/WACDIcBmNJ5Cp8UE
0Rl0laOiWL4N1db+FtfeedCoGjHLM1EaxuynMRDL3dfljDu8DXjm3VTSoWgU3LBO6IXTuDQCUH1c
jVfu+6prwjX8w0baxhXS2rtp6+rqIo0N2Fegc8D7sbXfghCLJpSFbVPQY5av6lsP3n12gMacjmd9
0T6gyrSNemlzzhCPNZJ/n7vtturRA8HdGcNz6L54V1yTkP5kDo4Pa7QZRMqSuAE8tzu48LKnCsDq
u6y1lQ0jS+Q+cFm1UUo19ERSE6KGgW1FfgnGSmcD5VMmuosCyMUEDlKfYbeFtr6FuDpUtORvx1Hz
tB3cQQF6QnwKDgy/xlsuNQAriAXg4Db1DY7LDmudCakNxfBAQTOa7d4zvNvtP+3GP1N+W1QZjswC
POQLvDbJ9hmEMJREWzFHk9duF7QEapUYXJ3HzLJANSYb65Q7EKZibb1RIZmsCS/LQHZhR/gIUx11
/xAMAp2lGG4h8CB3SnDvQAhGlDg9nwJAFkPSmJSZDXcbluU4WayvFv4D1hmnj/PQf+Y1Ymv61msH
aCTY+f8HGrm1xl8JiPzgRcblx8kFkGfCJC+V7SGWv1ZcChcbP1czFkgSv5THSJxQdtMHOKZCaTGo
fw+owZor7Zhf1+BfBXY738/BTw3F73dXunLisPhksG7ECoY8iqwZJS0aLQdQ+GjlgveqsG+i//ZB
7L1cC7dPhdPyScjy667UwKv/64K0/cIx3KXJ5CpfZix9XMtnnO+LtG0s40DonNaaocAo8+AScLKP
ZqzuCXXyo6fZ6iFjDXaXXhzfMqRdHk7vmVSkQrEfbyAjSTBUBjpx2ky/yZtlJpYJyhwhSrLf/hEn
9r285YGSAHGiiHZVgw2ILpzOW8m5404DRumfnqz29qd6AO09FXRo68kr6UE5NxPjw1ap950UeCl1
XOOu4FtaUYtM0vVQqXyLQULwEMn6mCfHhRXmVUzVq51Xlkdh96RPpBF3gx1khW7de94Zsfv1eZEd
EER6ZY3VGdpgPGXm3jKPZ3toFAka9XegKB1wofvvqmZdmvNavuLEJFg/BcW+J/1mn5BMaMnUqJWv
yn+Eyhg6OEno6QWB7VwK5SApB13rZdYgH9U/gF9ZxDfL9AabX0mdwNEWn8kQPDzAuTplj+cmnRpr
IJAezoRy30JECQdXlq/L97EOkvk51PqkxGjR9koOjkB4IfEoHcFm6iPSh6RNUFHan38fRsg7BtZg
m4/pUi6SwZukctZBjNm0wvzsr/AVgc6lltpN26amv9xEoTyfBAXDLrvOJtrC7g3YvpIaDPzedcbV
Q6ugDO69p8+KHfDyNyAOV9BZ/r5DmZspKh/EyWOEa463sIIc3+cTk8SPC6BqAA7ncYwFL0qlFaFQ
KVZSU3nG1tjWxpp3RUHtUZIRb99w0K0BZ77rQzDJqdZvJZcSahM9qcm5rAuWWidLpJ3dpo9gXulk
dZgSLHY7+y15LQHhIZewBVnZ1PVZ66ecanzH1Wa6eqPsQK5ie2EuUTuR+8EX0Cu9DQutUm9Rixpe
pVwFpse5vpaCCnPxcJK1cxNQaCcLT+KH9iaB5svhrJwdVTzuz1mfarkJrvEs7gQh+MZJweiVd87y
O9MxNWfsSY7m1DPSmTnXsLYdR7BBMeuUirrMrVIEb3yc75U/2Ol7H3meBZyyner2gwldm9HBby/0
TATHnTiCvX8s9CXs9xfYc94GTWmZKjqGvLk+I09Pjxwr+EFrVFlzPlZK/gRYZoDDNdQaNXTEDkwG
Uu8gFgXwIFCeiQutf+NLs/GX+wUZfdGT3EA1PUcjprGwIaH065YPVvoKa+R1w2Gb4Lt9t/RYlyMf
nqrEPuvS7LrZgcNplVzUM2OhusALhnFrC+DKx7S9budVJi0UY4TVBYiu/gUosIkgUzwgc0ZTxPVW
fFVELIdJ76XaZJpMKVV8QbO+tOiFveaCFnNLpiV4G7Z3ltnr0Wv5CNz5FCOE2ewVdPrHvAti+1yp
5LEEP5Umsca220grEhJwyNWzb5Dqhy8cVC/EhPxc+GeFKvnAIt9C14HPtDKBIbj+6bwVofc2V1bW
LlkdErePIQ1mJXr3hKFTUFx9ezyQrQPaKxN2hudFQFjvHXXJwYvBnWdDI70Vny8k3nOUxsIqVHI9
TytGbE6F727scbo5HUOWOtEW+ZI5mLJtdeATTgqlb8a2Fgrl1eo+r3T08ABGa4LdS+CkSCtk6WOx
OZi/FGx8b+48z5AOxcd5+f+rVwCLudvdG9QMTLr42b4rM40cid0i6IVi/nLiTQl2G3CaqgVYItO7
mhQKG6sh+FiO7ilC2JG4rgJXEcjRtyzl1sThVEQqE42Mr0/o3YsEKLstnsl0ag7nyMirjKTqQNWV
5wWsZJMbpvX2VDum2tcR9d34TLC3uDbELeq9iQHfluY1wxAsrjqLxWbGw5hWHkRnCdA4SlONxWrx
uGIaZO7DNwTCI/ahSqmCx39AMoF7fFiFczdgjNCJ9aeu56GvHTjQWRiB2bW+e0jiaiZS8xdZWdtp
TrmoueFZb6qn99qPdBIxCZ0u3fgCXMVSK+vYi8oySkw4NwE7PuyepOg4KHCdrkyGiCmy1+3KC4Uc
oUZNXlm8fI8PMFfKKXa+fMegaOXAoYkHcXx+CptnUCHgniM1Ew5sMzrBPSQUTI85HNGJBxXWkJKn
YNQfuO2gOybA3EXllsqlof3svGeKozk5iwMETfExPAZm/ZiAE7CRneNH8K2ZrwmB5tRLcZeq1H/p
RKQKxbKNJsL/slaJymX83PnnaehJo+LBi5GjigHn9/DEg3K/1iLIdp1J7D+Uh9OUFHP9/dHv44uL
54V/qMztS8fIJutdw/M9b0Uz+UeyGxfR1HtSsqmcIcbNdSN/9awoxOdC455YDxyuZ1edjiPuADhD
rkf/QRwimdb6HFvzCcfG3KAqSglQg8j9++W9n1wTJrxXNV+Zpij1aYGtPizhUp8PCN//o2+/PdML
JQSVA/5jsAv/koExP6Kbla+rWgpdcsjZWr/lkvauKVOPXC+O/GuhjYYRDdAJi5/FQtPvzUnZYFKy
fem4Mvi8u2KIVT/xUGE4yCavmaPDpuj2/6atxajE9kztjObmvCqgVgXDsmsEDGW9gUGinRdRzh4Z
VbVgj12LoxHWQrIV4tlXhv8EYKHXr1APx1JkOxYnXEBDRs30kL81QJ/e7uZ3nti+E4YFputQHkDf
UnEw3RWRn58zkEE/KZQ2lG+DhkryJdMtmIAnr/1bGve8rgQJASj7upfWi3ZIMV8k5Mz4xasAeb4A
xnzyexHo4ntlynBuinMwQh7hDrSbyuTQwip6XUmT69xLQPaSPfJLH716p6+iWfyprO135DUw0FqA
m/WUisbunNKPJKzfupLuFdYZJA1ojXiz+mOZYLV2QvYcUNvMp71MG8ziHE+kxoqHegOXNGkSt56n
AjCIMLtZKpKgsePbNj+d3hXbUCqnz3mzcaj826Ig28JBK/XiWN8MzKzjfc1vwrbGJI8rA4DzLmjf
EeIMHYYIIWne+Eb01ArVeFsokh8oKLZmqs5IayCY30VA0TcigQ/qP3IAFrAzeGHmhT/lBEBrZSu9
AhxsrEQDQJR+uvvTCdLkTD5oc+tpySZgBYSsysHaA08cIeZgR+RE2eyUOdU16J1Ln/8kwAQwYZYQ
JvnQUpMBOkbSFtPNHtykk1r5YCNKIerRITEBRgFb6l8mZ1RCBuPeDZZQfJ4CNcYTtHpa8yUdwQUx
g+WvP01GJkrOBiDvwVkWBC9TBW2w5Cy2ZRrl1CwULdEyaQXn6Dao6BewGiRUXfXoKjq9nVLbOdH3
LGsKf2WU9nzkal7EUHdjrN7qqHun2e4DtQWsIOLqbrnrkqu9PNPVur7l/Rs+SeaeDqblWmEXM73q
vckEm76IoxQB8vaJpcg5JSW0+iZEu6KOp7360boEtokz1l9RuUdiUhlaGFVDNHyor3JViIO+P/UH
QMnx9XKK8G5dCxhus6H1ESc0/AMA7c8beBkIy6OJItlPY6yn0FrxjUTL611UtvfoxBhL0g8uwJud
tG5fEfQtr9AF/6I9CmLHfsQhilAiOzhmXtO8xMpsveoDlFPnD2x9p06BUL1p73WX5W4uSWld7J/Y
RSuvREXmUPD4eiG241yb62/JORpZDB48sBqKg2jAaUwME+jiyuoX0BXtk1RAaeoY1q8G/O1SnXhq
kgsfDUgu/QmpT1+EPfytMs45H5xDUdczluzGvNI3+3SX5rEefmZkU/1m+uWL43F7MVJPe38cuIXC
3I9tVd/57y0dHOeP4+66H1kmVL59xlN01Z7+DLpL4BoeCeltCjh8Izwn8mTbMYB/ptaPs8EzgJlX
QJNQo6jgqr+JzYZvS5kjy67ZAybffMAND8gbJh5kKdLbg8TEvjtnw81EsMtebC/8XwMeVkuJnrE9
YJ5HjsS9ZnHgdLmzatn+0B3hrkeEsWEgGgv2hkW5EEC+nVR0gHGJP4dtTkKa6xG1htoLnn2uh2rT
Lc/g1pl0YS28H27OgEZQbKrQPPhqRByuT4KPsJwwwk7uTCOhHBXlCkQYKHDPAjmyFvgJmIpVMcQ2
TJb3Fg9VnsUtZ2A6C7CGFSTo/Aqwo9U2Cec8YdKAIolW97BhjWtiK/SNgt4RCgvDIrzfiIscmhkG
x80HE6dS8XzHdi+Swv0sNJOYGfa/HA2xB3lAFswuV79qU43w3FNySAABxgZNDPBL1mF1lCSR/+dH
TyYhEO+LfhsozEjYrWRo/ZUtvj8RzLmFKgaBQ0FkbJYNafINAB0Qt6ZQR4/VW8IAeG1KAm6QiBhB
c1y9/WqTo2reNHxBPHRxP3hhlRJCNXxjQIub5NOzYJlYmHRMJp+jwXs/U9OdBAdAMnGvjDeWlZxN
08jBpzUHSO+VJtBe3LEvHD39MG6APGNvHGyoZPZ+/iq9HThop3MuNR357ewJ/b/IJb6XzgHHrq65
5fvOKqkA8XZKZGXLTK64z+5RXbjx3oAvsBh1vLuuBVYUYbEMWUR/l8dyfW4LsroNyQfX9rmPpZlV
Wf1uJl6ydO5TnosBZfG/RDX/e3/T/pH14chLc9DuITP40Pj53x0qGcgUsAqwcCnrAwNqyrtasWQr
tKUFuLwwlDwGJ9hWfQ+BJJ0Cs2mf9OTiK7mXgWBtfS0piDQ4MDt/FAzoi+M73Fn474zzL77wfBXp
4ymH3A8+Ea3A5fa3n5TT5wuEoOnht4/GyEr8Q0oaVQr6GzvlLqmz5oRO2/wryMUOxeriRWjgh3Km
QZI+J1jX6jAiPXIYt6IuszybRwPMnz4WzXqm4V2YLaP6tEINcZxTgtF8ZtkJQaplIMrdn61E3j0W
1L3xDGCFKGmEv3dc61YffIh/zviqmhmgeChMh1oaZSjVYqYFeyI21XZFRZ7of1TTQunaupXDoFkL
rKWyqctC5GxS+FYxw7Z6csoayZ98lsUg415y1l+jRzD++nowyY0AxIVxciObHSiROF5qzg4u5543
Vc+L07XGfyIvSKLPrzwJXFbdD3w2gNXtcI9AFhUbWJEqfhn+Z9aISTD0vJ/8bC9lWAG/EkNx1qV0
+L2gjkL1cQ4+CZMek9nf4+GGE78Cc6O/RyQRJXkFSj6/uhb1GLWqR/huWG4JxZxkkypwpvgLdYcn
i9mxjfkh7bpVxyVXvc2r3L7uOK3ScWuL01JPgHKxk8+n4lgZic5Hw/O1ClKqHLiMvbKr9iRD1U/i
b+py35XGYTFXY7JxWxqx/u3ZBq6JLLH2tEj7NiG2ZoMypk2T7136/o6DNyv+fFj8VWJ0SeI3xaOY
rmwUsR/AR7jwImmCHhdWal9/Fi6tF9idiV6asXApRavT6q+7AkbjM1xquRvcFt0vcussxVtCeh3I
lmX/gHzU/tY8nr+0Fnzj1Nc0nhBAMFrhh1TSE3Z8GiLoMVfbpL1bLgmge6+Stm/dIgCYlHRhpQWT
oBvnmOxkR+NHJhf+KgIcCTLnFOZ6W0jHcAbCxrrZPPp1mq0YjkK2TO96scY78VurNHZV3WefDJ0X
MFP3Y2OUEEwEV66qiEr+v7Vm22N7WWNWyWtqghsETYJ8IK8i5lfRBHZGWW9PKr47NqwEjSUDsqs/
9qWr9qvoSJMFxTrehIU/LV7UB/TZ7xOzusQkW22rK+8caUguyftXuQ9JsTspqb3+D9R0ZheHaoXt
GlVXUajZ0A76KXRb/MYokLISr7ze9fQHQcp6VLVU455NHUQVsNVwGmpeInvxZRQAkctn2rfHf1Vp
Vm5kFDVQjWN3aCex/HfqnBfftq6QYxoSB0ykLRSumWmItGP1ZkusuLYPtBmnABmuvkL926W1qHsq
2XbTj1J25PkjJsAz4YLxjC/rP0ryBzvqX/wRt7LOUaQHvnfsehjdhSCVokI+hOD+WLz4GpzmX3GW
/4zdjJTi5w6FJYtoEdQoECg4x4oheN259MuSKTkcztUDqkxCK64FBxnjH+1bIu70GS3YLXSVJGGg
+x9MbwIFYxLyD+A0qgRVkZDSuZiZEspdJvU3GxLuVfp2kE2Me2KgKLz23UlsMFg7rgBaX+/zkhON
YMhbnLwzWNqyl2cqh/fzaDiHLUKTLQswSb6jO0WH1zQ6DW/wbVci1pLBA3Ed1xrB5CnCI3gXpwew
fCuq1SPjTSeVoA/xtOv0nlMC53WhoYVOkIEmPhSisVYEmI5Q+JhT0wbxuMu4iIHJElubLYl7Ntcd
6yphnQw7f9i9XnuDTauDduJ3jXiffvs+e6KM6btaLsIblc2VpjMA8aHKNG1QqJ3Oamt7CyC/hhbY
zuupJSgfRuFOZX6mt0B8UtA3qJLBlsQ91tvErUn9alUaJ9V1q2EVCO2qLRhOr5DezvVimOY3mLRp
cRDCk4BMvfTZ57v/vdP9NH65+pYUETEQAy6i1lWNEq65U3FTBzAorkWlYbtGmDNwuZcOyiVbtie/
URbb5zqDDTw7TZCPuZ342cJbpf8BNGkZfHh+EY1m/WggEwLYA1JsnA12xtALvUv65HviV4ftS5+q
kF+k2NXhUV6jI3hCuoQBGWje/Ko5iMA+dXK7eAH7Frjd3YeBY3jnJVGbiwkfWpnALi+Yj/rDsOSv
w9VKIr1jklC3z8vkcBgIRW1Fh2CxQwpyGZj9JnW/sNdYmvjB7gTyhpgAjrk24PbbIpJx0FMvrCkH
iWrq1EwLs/Qn3mm4VjpJw37JSfzxeqTM1FJhaWmpyrJvZrxPCYKavaAqbb7fDSJi92Mtb8REsCbe
qBsjAqQQmwoMuGuTr4y0onfHi1I0rBSVrRBgJ/JS863qJdo8DG8LsQKZ94++UFwteroHEDGRJ3Md
zsC6ya140x0qoFi4XMARPhVXabNO/JO+lfQGQ7VW+LpDE2AA8zqGtiPbQgxoW/eJdmyLWszohrqJ
F7+0sKh1ugoq8VBdHcqRxszamF/jp6oFqQH4XMcXOw/KVofHRSl+/Z1Lc5WRwp8vWuOvHA4vlH2R
rqYquJL8KOvYfftkYsB9J7DXPUpzSN1xm0oBW8JiG+CL6ogv7lgujAthv87hPbtV6hw2zcfTVCe7
WRLvPEKNmEKKNVnnac+e/Zhr9Vr/WLm4iwMyo2tZDDqx3gI7Qp3mEC2vMeYIUNXNKxwCgtItR4IV
gBxt4N/xSk3I5N/tlZcpCd1ClGPxZg6WnWWFBhDfwTylQkZq8h/4zT77JuUbnA7nNcK3yukhfJQi
rdODQbmu/bWb2xWMHVgFEAjWYWg5ZK8dwgi2Jn60a3sBDBzEQ7U+hS5WuL/7c1zXX6YzKFCrqAiy
PVXgN1wr3uw0pwd0/mEhQBlQ5BtdB1cDUgkozfysMiq8rXCaJmfB2GL6FAj8QzOBJr7PPBEMtwCC
Fi64Wx/b/tVT6IeStH8gn04ihQHl/gEDDGujLejZM9hcrZrFJquWB21/BjMZsW2pPj3OlAU4YQfa
4NbhgGFND0TLHxEKI7sBe4g2unxWpwUeFmzwl1pFIdXpZBAbsnWKrOMF0HE9n5O0IMwnC355N+Uh
mgbVfBEczqobpBraeBWSR/4gxM6/Bi+gsGPxUEQkXGyciTbfUAGzAeXruX8sNQ91r9A+nuZzz+3j
lOtu5JYjXRJFELCK6c2ZJRERPaZp2Nb2BNFlLz8k4MNAWaeQ2ySdTwgajnBNfWHATb05UoB5xsWR
rdu5HTCfXMwrBbP4wa9n9MZzuPO6yqMm6JKVy5Wj3eYH3QBoQORIkMhGX7lYq1uVicnkRqCGprEn
nRlHYQ7j4UxzKLED3OU7agLF1Sl3rVEwj+IeyoY5gDDuRE2Dcty5KyOGoTxxRyiKyKb8tH4BTlRb
xzZzqjFV2TQtTB7aO5nzHWceMht0l8C0ObUsfmvvnsiDH5hsIPyatNQDmjc650nyURAXVNSPVtYH
N2/j9AxUeDAKOtOZxASYERmLyyppgY96uH0P7nCi6YVSNx7/zg6oYqBPATjNXbFhBAyfba1w8Jw6
9LZfnUGxypPp5WtxEAcxisWqjcocKedmSlBtdBO9VifrZEDBOPJo3j7aEYTGM/CyoacpcO+8Upt0
IkczL1cqbOYi1vXQ2zY3D1zTNTLzxk1L4ovQ4mbjiazpRnntEztXRhUalv0bub+pixmHFiI9Dj+v
Dz6MC6i1LE3zA2UkS344ClzEua2ymrM5wnw0xVK4wjgM9E8UcdtvDvBDv12ZlBJpZEMQBt+qy0Cm
+lzZDXdG++fAJ2uy+RxYn2gPYH76iu7WrC/kO9LN7L883ZDygxzofCEuBfpMPpV1SCJP/ULYDRRP
FbpiTQB1uOn1fPXLuP6OkPr0pG8mq1CVJFf1gW1AlmtsV2WQDSErTkeF4Kbx1kQomTlmwXKIcDds
oL1WX9A4tll3VFk02MDVwpynSIm8CILlKTspZc62ZqP9Xgg2FDCIclsy94659aKKayKRrmzJyKK4
Hx+jY3sWB8qwyDcL1MsZPOtRYiUBPfyzAp155LjJwKShlQaBGU4RxCzIpHEmOOWNVcK1Zxxf0dpI
vKWvz0i2v18ijFC/9HXDZ1HlahzLOauJ4nZZ4SV8BDJPOT2FhsEBwFHbrnSE+J13Kjts1rzz/neV
uDcHlu25Ct1nfl2AoWVkWdSxEwCqL5+XiwmYsDC0uS5VCRk0h4D8M/4pmEpEvhQKf9f9/04KlMbQ
tHqHU8HBoU0InzQ2rgS61hnFQiDiJJQP08VOFYdzJZiL3lDbNFpGOZcq993gBmXNBCED3PawiiDj
6hHgq7dqldwAfadMqzXF+u8jTaGz0oh2jns3HBfhDbLBCoDhKLSKKOaLaGWEY3SvyTxw6Gb+MvvD
92ND8qqKEUs34lr6b0ckpC8B3o1ZOu3RTRRT9o70WzLdTTek0T62iYg0kURwdI58HfYk3CLpfcEF
jbGiPgPLOu7U73ZxT7vCHnetItP4sI7rdHq2WgeFxPy/qbW5c4EUuSKNmBmGHMbOGIGjJhToVIdU
dFI+T4Y/CrC2H5aVeabB92FYQseHUrQHxrCVjM5qGgyzYwyoek+/8kwKz9IB7UNBA4uehFG6I7Dd
8bcnukX6Nu6wS0j0/y1AdCeRgbcIAZo5Spke/lDZtx3jhdywMTIgCp4iHW0tNz0SfW4tbJ969f6v
GmeQ9c/gs/Shv6D3Ulg0zZYFfb4ngCghk7SrpMWckBSrWp8BKdpvq6sUVLIIyX/wnBxEoJUYWfK0
tcIz3eBHIFpZ4UQvsJYx9M0V4uWWS4oumLRF+AHEqkKDaHUvx9qwxYDtXRrZ6Kp5fvagbmaOxRwi
0KBAa9/gw4bo/s0f+1WjdilvmULsoy5XakXbFjg/hFISSIGhaPEFyzQY0n28tkHwQGs8G5MBEquc
V2W6OKwAn8QSi4TaRViWtA4Tx4Pdwq7XSno0T2SW4sHKl44MWMm8nnZFnmuU/DPUGFNyCt1mU9S6
GGvKHDprbgXutZMgbRXtJsal1IAIHMZRDAijUZuxybA31wKrc9+yVd0qo9j3honY+PtnE/+rcLPo
EdyfNJ9D2Gn1HRNBYmy10GiH2wmbs6AL9WjZOmPj1q2Jainq5nOnvCQnhnDCRq8fKL+9uieEylJN
/GkPNvW/hBQ5QcbWz/Vfe+ndWiy3AHLrd2ilHPD1jG9XeEzTb7/bPHJi2ELNQs6WN/s2LAFbBScR
mTiXjy2gh2FCKSySjrNwXbu5f/orLiBJ6lWHo3hfZSvcoxu/Cbr1liK8/3Ze+EGWrspXO1tkIAOp
aNUP/60uLudnLQp42yS8wOZrzOasO6Ptbd9p0FJaeI6NYBqNA9hELHpzZuael3TaX6x2oCwTqb+5
kGv1KQzz5mZYnrZoYaZ4yuED+cS7OdCJmpVnJPWuYCrJRtpdOZsvh5CxnF3ompckeBW/GCdGiuap
U/Qx7LJtL8s7bJnAxYnq6uY0ruixSK1i5q8N92kmI7yO89cxwI7ZzttVCUVVzqOeCJgSLpmvFOH5
wwdxGYNSToWkC4kF4x1RccGdzvUndBMWy7aDTEUI+j9Hamw+qIEUJnX84TTV/SQ5Fg+XF00C+dbA
VZPqrufADJHxIyQ2/z7uFlUoJu9FGxaA6bJMan0EkOx2b96wYll/C9bqLnCMWlr+IfHCqlibpCgg
ZJkJaCZo5etTVWJd4JkpssoZHLpvGdPH9hyxSGbWFCYO9p4end1W1DTvdCoX4FJFT7WibEqIcjoh
KDADJ2wfj6a/fSPvuU8AfSwVf8LZpZrTnUAFJ5aJhOJvZ5ZQBy/V74Gsqo2O/lEPHqNNztRir/LD
FBiorKF9gjuF//gqTlTd/1+8AajshWPq3OtHKXaq1hVauYlot5v8a0yJr7D2eP9YsfFklTzilBJt
iPKs8c/ycIMDFPz0Tk5LVARSngo9gYvamNWVeNfwo5IVrui1EDljVAEozeQJ847z6UgWeXvnZ0PA
nu641bFO9WTxj/Xhf2/cC6ty+tf6ZgHSfG6tQxo70a/GABzjQvQbAwjS3UlrlMs+g7WXkCnLK3yP
vhOwQtegWBdsNsl30Q6eaGtF6FJjI9mEsV/IHixPVRqBRCblRdu5cAjIiWI4xm0ejeO59JWbExJq
nkws5Uz6nwVP44sgrka/8dfMAXtEua7s98TJHCIDykkLMwq6HDJj/pjbk+/7OF/IrTBIDdjVgQaF
q5a0+t8pixiu7y+1SChDrYJG6c1e4PFI+N3Tv4GSGBlYW3fBHLrsnGfrqyPCtT5V9m+MYvgM29OG
cVWD6512/PLKBaxj68NJ89fvu+kcuBJrNwFcRw5JzXLO64a6vPQSMhOw3sr9s3kHpNvSlI6i1b7q
5LFSAROnVPq/E8NhOwtNw5OqEZYocFi/k4D1UUUqojQqDWigxp0XISc0ezIX8CkKW0TEYXcueNzM
PfEDVBRhJYmnBWY2rBE9GJ5SpSfLj8rOXSBH98bP4TLdAF+YQ26+AnD5LGt1RrUiv4rzlw191T3e
FG1qUSTyWDI7NSbNT0++QXy5pdj24siwGRsVzr7twW6NfAvGRC+sSOYHjDjmiPzM5kTcdPDS4KYb
Q3D9+7ekw+HdwhONSSayY0es9HyPUDMDkTZIllZ1bU2oRCSwDlt0d8Yo95Ek0k/kWK+vokozOQsf
gHtE+5yKVSOUSR47ReLFKoRMr/z5puSd2RSvS0wxFIRK2u1RJgsNScu0EIe274uMcThiTDkfG5qO
0g5f1X10R/KcwlFkY0yt6q85ue94LCmJr8pc/df2lbRoqjzq1lXLlW5BPqgiyuIvL1oQVddXOJ++
EJve2HkeZ41y9oLp9LW/loI9nvrfezSawNewk80FwJVGOymcAqq5A4neiXmhQASbPW4IisUkWbuP
gqG660HzbBvuxEkwdgj9wncm5tRU4uTP/NHGPGVixYN91FO6GXU+lHEiDN4Jd1TboBmXutPXBO8e
H0NxbzbWnw2ImCeNlVNawBYuwuI+lLJAnl+S67rdC/Ieb2mtRmtV+4gvlq/7kxtwI8Ylr2vl2aCT
bY+8auBUFHQ4OKM7iiQPL7sm+rnTTUgvtEzeuQIU4QXvImXF08fdMLB+fuA0WhwB9qJog90+hK1+
0RH1jopdhIPGgK1b6dSsGIwLHtRAtE74vbOVxYCCMXLSdtJ5OxpRoN7lGZ4YoOX3M4TEU9eT0KVq
IQ8Dcs4El27OvlFIvvhhJWjpDWuzHWdvnRkEXckQ2RIYuFYTXIsg7bxDAxmDVi8KDftxZqTxhun/
5YbMwoXIDnq7qeBmKe5cl+rROg/N9q/S1l2KkFcJg4nFk7sxAexHUTM276ELwyS1JHmQ63NNnXZC
mo0PtbYWS2F7SkP1BJclzSalB0i/8NZbb6b6SZQi2/3BHjxrMm79/DlGaBM6+0NnYBExNq60SL+x
KO042sagV7Z28aBXWCkzzF+D6GI3iCYG6cD1OdBi+6X00dhI5cposwpO74dAfYsIHh2Fc1gWBjPX
+dIY6s17WuN6qZ+4EgAeYKO+5SERtGbg76guYX+xNtv98mztcMoikCrncfJW8FzaQU+Drnk6AUHY
U53PgVazO3TZFqoOCb05V8TYXFPUrmUKG8s6weOdmhBq3OsPHJXhUZL9G89TgH3x/TVLYVJiUdWG
0OAWXIEYCxGSkRNVQrOVu3vUo2RQhj3sZYAGObry/OYyKoOFkYcy41IZ0O0pcAhh3S4LwTedTarc
uYDwYu0g0LfTFx83O5HlcImjuDuB8/JCrLSGds2c3QUbXHOA6XNA2h5oBGvbCePPdOq2VQCWkSS1
5w/UixXgM8ipjW0C1BnS2tJPU9Wu7r8udBnaIMXNI0dXbFpEuzZPLwoFAoHIXQ9kx+saH0HDGNiS
q1q8YHwJNUcGV8QX+04BvOwo53JeXsMPv444L1M8HeceIJSWErC1IL50dgIPeVKdZWIWrtUgLxrl
XjNhrclpGDl4G5t6dz3CRQTyLKbffyBSlHUqIIqbr5ov1gxwoSJ/MGXi4Bw4syT1I2rAZdpNjgF8
9m1OrHZ9cJBbyy9UTrJ2X9qSSep2kuDrISjvAXrqsVx5aih0n0qYvfG8yoNtKuiSRSX+0wBUT/0m
KhywAIAMcqSc0iRYlmN6St8ta2WDOLQ/MdDa3WjM87bMxWoubD3ZMTijxG80nQK6Wy1yIbZORV4Z
87+2/Jrbb7hHhJ3GBc/qSTn8jbSscXt4FAsA8+QPxsYQpMPDGBnB03bhC6OOu74QFfaovI6grIKE
SaOgwiZXzQ/aBvWz4BAYwRVa+LAPQpDC7KoLsu+fYjjXpJKXpc6KaGlyoLO4H3hrm7oJXfVELAeU
g0FyBTIToiVn4U6BIPw1qZYvjNy/AS6a56fhaYLZKgu2bXF/4lEx8Ez9tbvugcEYgoqiFdnJ26Fp
ei/Yz8BNgtj7Mrd4G6+z4d57uCEi88RaaoxB6pYbES6yATB7Hn7rDE0hOpTC/Sxcp9qVfJ4UUADy
6fwWl9a1Wg2eOZQfZJf8t4HJMjYlG+ozYaBc6+FGPHMkvT5/urz03jEmwNo2qOSNRIwOxcOKF4CO
eNJzLaVnIagpIF4VaBl2PHV2MXceqVhPWW8Z4MB5oNHLw7Ik+hxySfzIkTfNOfX+Zw+qOIxJrO6M
tSdpclh4KvURaxi409o5iIxy0ApL3ydr8pH67VXyjpSEFSe6cSGApv7aEVnNwA6y7tzvRluyJhpT
UPyn/6TLM9uUbKDzVQdUwWEG2vIBP+inpnNfkfHc5tmVWZd8u9hiQuuwaA2zH0uSMCkH84OVntA/
mUybMLCBjr3affgKnj89hpo8Hf49lsl7Z04eM9udqTt1W67ktRJVMhdsu6b0w4Dlv9N+n4brQtn9
5yAZ5Dj3KQdYWpFSFCC8mpwtkbkCq6TLvIcKFGs+9tYOC0/pYkS9FgdvVoxWBH5jlNWya1aovafn
C6QE+3S9QEMJo2plRTqchrUmcSDTw+u8OzupQlV8wAnuyBknjdjfiL6SHNHfKLtId6aKNp1WVAHs
nJxx1eWSeFiVA4DHFm0llDOVBItRov3Ufwb8o8StV0JWrOfJrwtPRUzOhynliZn+bHLFVgwXFlkN
ZQu4GuiJxu60uxgrErWr1ymKRBVKrC1mL32gy0gvoa7g1QviOj0iPng7OPoD/UTCVbMtlXU12oYe
HnwjrdM9QWRlEvffNJpHrpvvlOlu+VWRN7YfdTbcUzG83UX31RTMbmjNS5wZXe+59xVHLLJpBbli
TgQlNzouxc88a62urNR9OCRx+s0OZ8aLtbaHBDjQ0XFtO0kMNUzlK4MvyMS0zpsx8r7FQVe7lELj
jFqKwt9rAvFpOOO1AzrYpFJZGsp9Vn5DQrCdWG+X+1kL6S/PvGmY9IyActbnYXChfeusiyagMMFk
Zl0ErhyXnXtc+yhSCQHUrpR1zkODnwLTPHEDdx0vg5NOI6e9NIk7eLn6pOOYYRpcrERPhODi2z2g
qmRpDcPQIgTpKrwp00upP6hkGAO52YJB4F0iszmU1U9Ss7MOtroVrbNU58wzqmFvlD/Qzr3kCxLk
7jEDr4Td+5ed8/MGxT4CaBzOrTvu1/bJh48gBEM63ZMtsELMb7IPNb2hc5BniN0JkwiQqRA1cXIb
O1cpx9bhIbcym7Y4ObZLFFzbBC2JUWTOSnOpNPsVmpulkh4R8l285X1ink3qc1HeVp2Ug5rwcnYx
/d0BuGfsYPZxvS8BEl+dbofe3L8jUceRHk2oppFS40OwnHy+QIwh3yIzB/VM3FEAkG6JMkiftsOI
aZg7OPj/baq9fuOJTWc/w5QiNTYCnboxwn9j5TZqubzj69Bb6e4rbaT2EtEmEGHHXCzhEZJWiv2Q
k4pe3M5rLlM+xPfPkEd2wWzYCxUIeB01KrFLKbn+CJezwXTAsB8udMisbkJhWGnF1zqRsTC7XkzA
H446gaZndThy8/JDCSLv0nG49FPa8Ppt5bfoW0+tSv4GLjQ2Y5CEcx2L8Luls75w46IqA8IK9cMs
cDrUdDhkwqH76ehW2rtLha0+WuirhPk2maz8w3A3vlVsOfDwrQ8NbYAX+s6ZYyE7zBZm8R/snacT
je+FoppakcaW4CofwIUWmVavRfoOd9eC52jrFzgFUhmtBFxWKw9OegMYSdOsaoOng2BkAtFiZ9dC
UBzIZ+MEeG92du1XuJdpayG9pLD+lxuhHAovRrp13Y89+sPxxN3lLemK1Arb7YsH0BxMbwFkfCNP
OT1PYKUi6l/aYh5f/h2+pg7mZMhK8OjweLoSuHFXshjLNS2QQ0XuPp7yrxBNtvNU3X5s4xX+PWQ7
d66bVRZX+AV/od33j7xbpoNoBp8aI7sIDGdri7XwAiU1VlfDh+G9GMuKcX1H927732O4qFU2clOL
x5h6nSUgde0FVXH5uA7y6yE7YZdHesTTKpVlBOusvKnooFsuzmwluW7sZOUzBX9hAV8xnOXJ3loK
yivpn4lRAuwLLeXnfWRgN4K6cgmtMV9wKN5N6DMzIciDTkhpBgqmYPH4a91bWbDR5aEGgmQj50xu
W2FreytOOHtQl/jjG5izeGMhQyhuk9ZtAror5NXwsq99c91eJcOan3FpjgBNnKDn9VuNbrBav/aL
vbBiBaetYxi1/pAOHFRpN4M7/nIeYGIRSlrfTUKdLpOAOd1JT9Z7EroJymREsW+yr1v8h3bLeNay
U0Ka5RmRRciV1Vz5VWqwGoLHDDqUVgsqjiBpsHuWZnjC6WZHGMRdV0b55c9fr6V1pmqHWI8UkZlg
DcbJTVE6AvkHVyB1XzeVou57Pf0h+8uDu/IzGpI0HUxHGveX01LGFVpnSQvQZHLCn18PsIFmD00y
hiZeZ+2HIrzrPvKSBpF6NJ8Pp4MoKf8TFsFsYvl41553SzYsNLkcXBG73dopTod9RoYV6WKZx2HJ
DEsGIOj4tT39OI2HS0gRoXA7iwg1w2VFUNZaI8KGlKecfzngbfpNIIURStapSIRCyJmiOhBF+yfu
MBnXVcUIGsSdY8V8fW7/9FUi6e5Ru79l+59PQQSgxLp2yy1Eith6l+2R4IkRtQbMF8isQsLgHSAF
6pN517PiwtXu51rRm/H8xdlrgQi9MiOwkgv6nBRfzZ+aaBvMgLbONV4ZXEW+Mbuuu/3fSdwMlZxq
HFU4K3tWw48XnwoyFrScO4eVym+O8NIrrDCkKRBNl8eJ5qgtfSNZi5GDx+xKhc2YlfFGlxeUMcSe
cEC2klL2sbGOwHW0PG6rk4+6JutM3HM1Wmivs6I4h7StzIryQl98WvMC9JKE0wiT0McsFcwM2s65
hjjZUFZM80Qjj2jBeaIxnWwmObHIrJFA9IBoH24JSmX6sCdaDNro5iyyr1RsdMIi24ARIjr2Qdzi
4/02ioAFKJuXJ7L0RlvlnjaH5ypleV/rjX/b+G83E7J+PResVOXjhNIxJtHzI6onBUxNTF0ppdr8
RbY+eZ/1LkEutz9p1AUa3gLYjY2hyEq37pWCaSgXSJLGK6j1BEDeaHlHUfSJft/hHNqEogHn8ePM
FyF8cquUL6lHbWVB1z96h0uIS7ZWKp3JL2Lb4ByqbR/E4GXWhcO6t7ijyrWWqJMwIPsJHOVJo9YV
JYDg85PUfDHuZLfW/pQEqaXjWUIXWF5+rNClE/TiVZxhqKOo+QgoMllisJmCVTus7KiOBaA0/+tC
LNBk6hTA5McXnbXdUjeZfcBsUQFW9BIdXGnURZAqWDY480b4FHEH7iJfbvHLaCTzEEMGhqcbO/7x
VkEUqjMWgU+04hcQfkL0ly2jqVq6ZinTnlKmyd0zlR2wBLKpkynNaRrS4CrHsDC04G3Ama6kry1J
22LZfXmKz2w/m8f7c0H0ll1v1LFSTwio/KhQWCjYqLStxOKBqy3QT/9U2D43nQsNyOJxyGDvv8Le
ZmWLZU/ZeBHpbmTnaW2F6LKr9j3zu2/RUn7uk1lGc+2KoisExuLpqacyDKG+MkeefFCbX3bE/0CL
NWfdmvzqZSqwhNoqC4Gdnp4Vt6XEcdX7CNHxtdx6Z0yNT5p1bAF1YeLYxUFvDEDf2i0NqPucBfjG
l0EUF0KA8qHQJ4f39xZaGIcoa3rBXuhYbUm74AjCn7ZHxqjNHZuA4CK2DOW32i+4NwGJLYKVUsI9
GSeO1Nbr6eoe8QzQ27qYkeYpaHrM8xTZYArDaeFq3aMwcovK0HHkNLOZdbRC87R6XYQEXkbI+/mE
kto3AgqRLD6n1BJXNMOwvJi1BW8GGP/yX4OBDkhr4Id9V55kQLQglmGM8wBO7pmBYCd91UKVIMAv
jsFj7eXX6trG4TlwmfCfjXAl/HAYubJox3XGVoFG2bFVwEjrd9Ei4F5RxRR+eMRgzXbinhUTgaEl
Es0RVe4jaUBBeN5aTxIR2XWDcRrGP3kRB57MY5i6BZBgQTWDPeRg3QsvQk/jNfZ8MbdlvSrty+Ea
Zdu6bad8MIwGkuTqdoL3x0RtRvWxFDOAjzNNIeMFd+y5exdRQltaLiKrCWcfKu6jKUKSAI/cxYBM
7zB0Vv9wmtq8XtUQdj9RGXacfk5YEqDFRWD4ZLtrbGke1IumwyMVV49nQuGPccMCoTfm45Gepm3c
hfMJOdehsHDS9a0XitOV3MtEtafAkOhkqThtJJWdzooUO1TG/qB0q4xvnoJxYTnSiCWnw/4vgNiI
IgobkBXjC3aJ0HsKJUpO/M0DpeFifOCGzipw2qnlQJ+Y1tIc/peFRnfCB3J0aBwvQv7IzFMLegtT
04O8KQUtl4pYyI5NzN9BpeKx5iyzWnltEvTWs2y+M4jtUJ/ayeeGOKfbOQ5CKkZpP+eg1O2Ql34B
3Rh6orqiS4gu8FDyDCXZYIYeE+653DnG2LquWIs5+dhpAxyY251nNx5LSGPBNw8KLYFS85e8+Odz
qVMzdfJ+MUPcNBRP8tPcBuaR9+6uIqMWQvfA0GfICABvKEpcJHLSLsA+655rrt8ljCJkDGRQ1aaQ
RND8ULliTZQzBWuQjP5whGQ5Uf0GkVb1Dy2padkGUsoRRMpeoRC5kIYp6g2clVo+GGhxg7xLBBwn
ljqk60r3VY7/8VOoCT0o9yZOa4wf7H+SUEcnswUxmvD4pXqIbj+2ermNn8JOtPT3IJQI2N1atHAR
jBVnIpfQ6549mxF0AUBiP8efM2s6SKCN1eJYt0gp4G9WKzp/fqasrVE5SnfaaWyfTTYAZi1+nsI9
TmhSGjOpHYMLJH5AgU6bW6HdIz6tLqRw3mso9aKU7AXYYVa3lkixDWjR7nu7JNcYB4Qs2TZ1aeJo
dkUngxrFqbjcSrkr6ZLl8+lR25Wf+gb0QiT8Nzu6TOBoAlhZtRQqwYZ/nojbDekmHQMQHx1w2Eqp
+M47drcc+RfGW3cFLuXDLBzRhxMw8VhUiwqUSwjIqYOyUFamfK0smEVO0NTNB+n/H+M4B/rHnEkH
PS3ZGxOw0LfQfDl8RnUGYr3ndPt7jMuIBiAUeDSxEozRljSZM87sYeO6h3KaR/dusZcmtFUMajRJ
TYXjMscY7L8usrIhx/dgEaCVRbJwbQ5w7+heFscD/mDctqJqjNYpmbiKBOxNJh9VJOyDZG6Z1GD9
75pXijWGSEjOGZAo6oVoI2alqVBCQIf/KOm4idx6va1QL12ps8ADYoNW4pdvbDlptPM8GTnVHy2k
E2joh6HyqFCr0X7py7xP05FOJVLkrR4wxrns0/5ptClkqIW0virXyWe/Jfkcvf6MpmSWH6Tu6s3E
LmjhTw/jL8y0LrpGt7f7OAGUL+N2NlSJQiKhQ8g7i+DCRqVx2OhEN+TpKREnAn5asKCyHktarWUS
bDbl8FxKg7HVKHvdw9t9uiXjPLkE8yg9MaXsd7NDPvP59Cd/FiQFa3W0oSMLJBKv/VJVkTl0Y9eG
lQjNi8FWRN5cfFPeC2jHuXOnPLSMpD70ve0UuYd2APW9qnknPwnYinlc0RmdusvKv55feMdS/RnG
eRD2FCUYfxTjtlz1Fo+iDe2Bx1NZIUNZKAzh+ciDqqMZlEoasDqeIQViHPLMYWgT2+uI8iGyGqif
YR0I9ldCzXZtq6vSWzw+uL8FHA9Wg35WZXLRhCqlHmvMdXEgWnVKeX+j8XLLcdZzfbGM7aiG5U29
DULlZKXg2jcW0vS6CmEaNK9Ghd/3YgYYvJdIovQpQhX9rEBrhcQs0dIqEmeakk3Vw+nRYG+pN60/
/Pp+0rZAVN2nzksB7hHjn5AbBmFl6fvWj6fEKAO4Nz56733ynfyUMQ+3xZsms26FsKbR1NpfDxyI
wXkkqryIipYLK3Tyvc08UDXblMaToQ/dCXVKqyrmZCqR7JoYCDjBnx4xqRGjyXMLDdfi0CoNVkn2
yz7tfc8G5PAsZwptVTwHvM+aSE1CdKbjmrbpumvLwBDSMVzHz5vsyWKcRKJGqhaB6uCpReF+htY4
2SqZvwRuO0uzNgTueZrIPxmkFD8fPksLifltynoSD/PRFo1rR1UNl7bW4rUZdFIVM351klK5cmD0
t8OguK9sN8pwD0/KNNvgE3RFFG03gMJVIgjFdkjuPYKQUrENwoSILLck7UQsBAXuXlgc4xTwbtPN
Yaij10G+vzGRdCZhqhncZIrYpEg4wZecYTz60lmU+91hYUvXZHNjkQc9eW+9wamtewGnsTuCmFEB
gKNVZzTy4iYeQVOWXWgUXgT0bWujFAjn2AUkJENEPabL28Oh4qBWMaNV+BzTtXWVLziC4VLbdiY3
P7eakpLysH664wgJ9ADc9NN9G3AG7+frbnyXYqISKDrOOPYzQganKztBNNBnjor8Vnu+rVdBhBRV
i3cfk+hv7g9bA3rKqapxQvlbGzcx9yg4Ww8+/ZyC/LsYW+HkxfAR0UQxSuH7+wX4lOFrpuJkhn7b
wd5rft7VHcZvXpDwABHx/+Fmjf0qDPZAz8JIZ2moAIDnyovQmT5+Rely9qZuhj8ukqgNtpexsbOU
LHx0DBLHl0UTqidPqQse0cbheDZJ68UFR95Ysm7QPRRL1MafRTSYSdgE6mYHsFWklpTKelM01Yms
8H4K9IkyF3FdocK0xLvo3QM5IIG5UTcqS9Zp5p+0A6meMtxCE/pqRj3g+I0eE2lLcwdmJ1cU3c7F
7c3IO7rLyFo7/G2U8U185e2IzevS1kOJQDiuGvQjryTWwIMfG2K0RfP+MOr8IzfDcaNcSOF79wDz
Kikava7hZ0Kfzv6F62zG0geuixKXhfnWIT4RgIe8nQBYphLFlzIqbGWs98emGoFgf8rurrbDkw9h
2lJ1bXvm3YiBu5ce3Ws0Jja52kIoSOycCMNVYpbRCOpRjysVa/NViFfveSIWNIz9otRg1mmG4BO2
aCHGHjDDMNiQ6jWkKG+6aoE5JwG8Cb3FbsoVOMmybZ5Bc3GhrRHWGEAq2scIFxQ6V3eCXWA9JmsZ
lXyrinY/AHkcO2njDeqaKF6YKjiu64166lMPDW8M8gwH/4n3z0c4VGd4GRJsPkYMniujlRWvZ9gJ
mwC3B7p9PVdnW6moSt3jdcscNLhPCtKdAxj2Bk48Wl02OHEZUSzQahvEHzKHxxky6T1IEx2HL1Bp
n+D1co8QsT2wO8Dv+Zvh9JIEY+Ay3MFbS72u4bnotZL5CFSSkOq8B5ZLZ/BSfQWGTHNpLQGILZYz
kVUkqy1DEhJbwUpMoVUK13Mqu9AMP425nBBnRVu3sMAXQQGXNLVHPWHM689I0neBaTW61KuDPMMj
XsKd5UvxbcOSm05Qp/G2VGCpEIS0a1mK2YHiD7lYUXB6iHSP9HcyLmcfE7qRPkedDMUUZSb+l1UC
RplYrcwXSXBfQSt5vC165pOJ8Vc1imOdilGNtJIDJ2ZBK0NsHVio/6fBX7b6OwBvT/mGQVQi879t
gy8eKbaB7b6hlW1J5TFKHT8QL6L5slXFoLI8f4uWVMVyNbQvs+i4Ss//biEObzfOr8B/eS10qwKi
UERdv4BSt8VUkOeBFDbN8sMB3iOo49I3QhMCz98lzC+N4lqWAHhpysL8prLc1T3ca4RFA1bRNjsf
U246l+7OnllaJu+2y7v1AaqF9GELSpqUwxaZCotFTH0NCX1Jr/j/3GUGPdNGfxMnw3Nug6d/39je
fItwfW2WU+jl2DaOdlmBfHwCJCyk1VdoMajF4eBuxh270FwdoboI1/+r/1ykDoZhtYgwQc7ETYRD
RfgNbD9gCF8S6MEiigAeQbGB/n7fi9SeQFGdW1811ake1XSxsTPGNs9Osd52iI9JGE8MBA30ykhm
gx6EPTOMWZvBxazEYzGqXicuAfBD/GyhxTwyjXYawWrgqLETKfkaiI5Sjg6y7uajrWBKxXgpRMae
APgAcpvRhj6dTu4swJXZrBYCgA7rTSSDVGObqM7GwhKBSDEZzQyznddjc89vAHldakcEjbkRdMhw
0pThlWpOTA7garcegLjxMEOCSKX8s7yM3s5oHPdv0QLyIND76Y+nLzPxrf890WAGy6DNfWK0kDQ4
M8bnQ9/nvkUudZye6+wKU/KYWDNAsIK+6IiUUXf6KGFSXsNc3MH2rqUQU8Il0XMKIX7+kwzF1RwA
DLPgSIIxv2TaLBG9AukCVwxCsXWOmYVgd09iGTjmPvfWuTqn/Qeh6bwHQ9WoO3+SHI+C6bFk8g2X
riQySHXFjwk++r7XljDVC9mEhL9LWtjnCV1e+AYhYLGtW/dzuSYfXwND4VjbeMDnwLiql/j2l4Oe
cCNn+51qPLo3WwrlNelQX7+A2cDrbGexHUx2CLZt9FV6lxRD5Rq0RI+szzEZYNQVVpdTjwEMO9by
g4CWDZKDYdmI9S5EHJWv2JbYK7bMflwpWW/1s3h2jWuy3Q25f7uklAjF0KAQW3f/xcLiFb8jfg3K
l44pLXlQ2sBHQ4bs/lhlSx1x+VyuQzBmttkhhV3mZ/EkzMKawncFkh1jdMozc0X2lZKaqMIyyqEh
sEu1ocARZRz91WKbfhJ38usvgmaEErLNcdnn120Hls01RoMbgulkMn1A4keMaXggp5+B2hDSl/o/
M+Ir4ywbmz0Sq5v+jKuM93x18Kou3wJpvIw2CZNW2EkD39qIVRkWsjnAJsfrJnQrHFh4rGeIdyZC
4d8D/CAzjGzqibJKB3PZmkiHLJRNaKu7UFBKcbo0TswgY9HGQpyC86BdZRvxE7eQ+HFrATQFHqlm
KulcMEQGWYKrRd5BeNI0Gjd5usLzKx3oNg1eQlosFPMURDVrlo6PqlbzDA8PR6hoDCSoZQeY351O
bgJp5oAKRZ7jXrLcwXOFJqLNEzm20kKUGD6Kfvh6Nv8I9hw+/MHY1P/j3SH0YSK5MEgLWlzGr3oE
UIty7djf+PTza1dqgM/h3EFML8jZN65IC/a2FWP1EBy4xgG/4abS6BQl8paoF0Vu6dUb1C77WWQT
4Lll6Ct2ZYRHYPuRxrx2wf+wPo2EeLEA3ApikYRKadBfmB2Iq/lRTqIujd+pNfnRM38FoQeIr9rI
B0cR/Lqw0V3ZulArQ9TJf83f2L0R2Flb9DXVFNDmdTLKTgIRL99xt9M/OdgFlzAvuLT4IQgV3YJy
wCFG+qYXw+yY71QDJYJUZJs/yb1IJEQ9698NH37nUAwMKPQRy5ttofHOlZu6bgqiRd2OCkrCGHRW
SzWVnhKQZEyvKzpCwmMKLpTL6Dt5bEGO50hSd/f3yNa0A4PvLOBUPY27e6bgCVjh+RlfPO7M5Wdp
L6Hz/u5y+F4PQp+g0cwz9Ij374sQNSqmF1N9FqyO8Qbgoieo2wekEAVsAW6z5UzRJWDocUNf/NqJ
HqFTGnvOS3FvXidqJwVSE3AXD61FW98VCA1h9EHF0LSvDVav/KtzK9/ZmxvUFSu5Oefte1Dus6wi
QRPdFSfhgcLemZyvxyaX7sQ7dlvVcwDJQTl2RDwQT4O8DG49xbguK+1FC0c9W2C1sAWP8aaJVZaR
rl6cn2HgMv9wghS/M0GoR/kmCdW6zect+0NuxukD3Fi7bCS5WFyp0LFntEi5IBh3t5eS91RIFbOE
BlkTyzDngLnxAX7A8xqQkwcmUUF038bOxkb9tTusbsIbTOMzt5+x+QwV05Lg+dQZGlaPQWeGrX+k
es+ni2eBfA5gUf8TL5C4NftDHuq6UY07mEq0Y8chW1pb8k5ynMYvnGJ4mSKsDbjTuKLehsfV7THy
xsaRVd/pr45869O+P7Zp7/IVFs7WAscU/+TlmShXQcNWWmqn1K+wCU9xeKOPb6OINPgUXNGFbUoA
B/5gJQnCICqD6O5OG7yXhObXOaHMeXx8JyBAjdcJrfufZms67Krd/sWdplPJbdQCAif+7YAex466
sqYXJiPrxfnykVpblPI+SP5N1eM4xWN/oNM0tlxb+WH3JfdSv1dZ7stGeLyi8dY4bm7fZZuGSWKm
gbdfOOdtIZQNoqRiH5o/DVvEIaxzb+D3qAXvz+9leq6d5goJ7QxztNBrz/yG8imHy/BmL50uS6sN
mNVgBp0tqiScIVH0BTu64zV9Q4chcHVwwxbV5GgVl8YesIUfPhtC0VqD45HdZz2vgtQt69H4JELH
oUK3wBMuhn+AEuyrUs8bFsErWKUPVSusHcPFqbmyivFxPxjeNMAfpcfXK0/GFRihqnnGYPTTyIsb
UVvt+XAS+n0yT4PUmsDqmcAYYSFknbuW8xCt9kw+fMoSIWhfD487AQg+obUm9wY7GArd2k2sB6Op
22rngzlvdJ3J/8etbjxnOgtVpEY/uPQ0lKpZAdg7PuW7/UieCXj6f+ahFZwu5t14ATQpgNos5ZHP
fa6bSDImA0CfLpvy5zkFCmwFwYMh3Rl5nPOPxmBnvwKHblg443uhl2hiXuvNjXHZD4O2YWky54Zb
TcGrJP6ZPl64OLMGWNQJVu/cGq7j6SYsifBsj8lrOh8iz/vIJ2br0cdvgWVdpVRJjAAgvgCajwsJ
7l2DHsxfh1v7gF2O8VJrGu+SiVZe5K6GBR33aZ8uOp+M28Au1S4ov9kWsuBAeyh6IkjoJxkg7lC1
eW2+geLDwZS/iOArHph/CfEDTxnduSCNGAroO5SWr/rTJz319pTOQxqGWnZSO7KMMd/sMnEVt6V/
7nIekMvYi45ctYO8nx6tAx0c4ase9xnQVc94GxF31sziJNGjgnO6AXORywxQelujeI9Ls87JUcIF
CE0xOVdFupWBfz8c/s9bsMjiJSavh04+fZqaxPVOct/2tuD8abYV2TNLunO7S9zJ/h9L6lDeywzy
CtGBEBtV1f/qJKP4lkBlFeEBGIXcqZSZyOVIF8ZRpR6AxkeBBSeNcRGrMwdMxnOAScQBcAJMklWv
77BXesBZBN3LV4/NA9WKVtKtwWjpSEAFpBe2f/yQZcJpti2vgY/HOfy0/PnMtMQaM20OMnrNyenI
ryFAwvptaLHssj3A5Y2SByVaqnwtcME8FO24WFtCyj4+GOnY9N6LURQKCQdARlx7SQw9SuN3/Z6n
dj+l3+G0xeU1GuSqOwIXoH+lrdGxZW4KxyRjTnW0PsRwBrVVsXo85XophjjeZNXSxubVWLkx6PIC
8dIdZdStmVjhsZHTeaXlQK1vCJqfmjXgSMe2KYdIsh3vmoPj0YAdc55ZbJ2UxvBD1QiIiGX5Nrzm
gTLB4Q8vsb0UMHisMdJmuuaaeFC82rtLuwOglA5wo2S/ecCMXVD4zZSd3b/CHWbJLtsGz3kMsZu+
K3ZCcz5pcuHJTF9LC71FHDVlHHifimsUzrtw9WEn6IuegeJCKnLhInB0pftnohH3aDjn51i+vEL0
XbrfKq4+wHY8so+OxQNfXxkoi0jw+E7jDC8lJC6gk0SBTbEHm4X7JO69uQpseQ7OO2YH3TMPkjV7
ppkeZGN5DRzX7seRe+Vq83tpsc1WkDti4TIbrCt92EAPJAQ6BIcbjn+0arTDXO0y1GA2GTdcieKD
IajT/CJxMv0dpzQb+FEDcO5N40gGLbd74sbz4BSgaU5xBlma4gl7xi/J9/j+K9l1DVHo+NkKPajZ
xVmoou+mHI6gOlV7QSUbBHTxLRvX502wWyhZ66Gsblyl1Il46U3IqBiDT8bikZbARVolq6jeBypD
uB6ROkUKWfsZz9SKYVNFyIVEmZyn2/6omcseEDagpdkeTpZWTUhVWpAhQ9bvtiB4Mi7sDlgV5Zp/
Q0u/SdnXbaFFsP+rCfQT2ReM2+qRpBraoOdylKCEhzjKPYpBzjMPOZqKVU7eRgV1fT/SA46qyZUU
McNzpUZ2vK79HAEjt0Hbw6Vob9/CNtoHIMKNEiOA6qUOw+vG/R6wdCpTharUG+kKsi/5zr83bgED
H3qbdZ2d8yiyKou89knvXnYoh/CxmjD5axqIgjS0X98+3gs3igITYC5zqGnzsfPvLnZP7iW5Oono
v6Gg+r8jGHaQ/y24uoLHGvj3+FoAilZ3QJ2ov7X/BEsDZgicilgWu1bRAl2Dl95B6mNMEsfIhWYY
1s65739T0Kgb30x26ANGU+ud6aud7J20n+ppR1TEl8jdsbJA3a9QJ55Ta6rf6OvzdNbigj8dZ9so
Pu+mmws71YWI1mgDPUhe/wqNL+NgYGn2G4+xvFx+VWANOTIi/66g6ck+7kTJONQBi0rBbtgM0by2
ZNqbBpVWkFNwI3cxGK7rd3QCNiISAuEUiyOxOVchJP2CksYm/uIvfpSooH0I8U06YKaK/3PD1HQn
KdofGSK2OvzUvhkAlv7t1ZNIXBqy4LfDxTslMR+XrrowG9YUApON6AH8MgTVeVU3v2vbmEQTRfyV
xuge2CoHQsdc00uRdV0MPhn6DbgMMwybVekzn0b03XtiOcbbhBM8CiEsv2U+0R3QkiOjS2hRYE6b
bOnTbYeiy/A1bCcjYtj2BtwNcEWLxLECDf6hil8u98onUYE+tVRs99SbwuYdlm9tBfDnZx0hWvvU
yUzjPOHSPV7cIUy0QpbOt8q/CAObIER/JCMKnvPHtIakDg9/JhVA5t3BR7308tu/X01wgA+UmEyi
+ddI/KRU4Yfy/xQfC3a5huD9jGCgKi0i+Le/E0jd1dn79a0VDc0w5yheQ1b2Rur1YMOeZFO8kUsL
KuvOeVShMon0lJj4Kz7vL3fPX8u3v7Fprh5GtGRcZFMMDZ9OEAZdK49sMBAU4NpvgROYKd6WhUjV
fimmLcI/ROBLTnNRAyU/srceJiMLKfhXPGR1sXt6wLpJYLSEJ6jEwZqMLQRj1jMPBzm92yg3cS+5
YqQ3OGKOcKlE0C+I51Iy7K/HJWosdTNv35KKgE0G1VoGWOwtF2gkh9DC9iBkUdlaRjMexgFH7ndB
MUuc5LpkFzfRoUjAXp8zx/uWp2YOfk2/6Zdu/ErlxvP8VtIkmY8ZsiTbb/0keUhdsBVJC3goTu5/
hlqaKUH/qQDlnIeGlkdekJQ5hdrA5kj3EPnKH6/xGT7YASk4tIAVnqHPv0Aek9K3OAT5+UIz22kZ
HIjNN3ghrKEO+cMM5qbC2qjOXW5CyKdQpqXGYpLE4ZwoQrRny4e4mi5ZVNgD1vHbMpy9ansbdeO0
4I0MSXfZBqrE5p5Xbc2csBitJRjAmY1GwX6dWBrwlr3NREYPXB+DoW6tG9H4wijODxBvMNWvNKD6
RdRotAVgjHMTlAxz3/FUZy22B9hBAeicM7vqoucfBzg1Dy0o68svz7JdmdbOIBqwfJST90ErUCIU
7VeOtK0BkOksMz37Fv2ji9H1nlB96hSfg1O0D62OXrLxm8O541c4HwCIWXcLTcVhioKuBPYMJKV7
IsyZPLR6EYv9OFVP3ZVqkuQysCFt/+ELXsFa9jfY5OAh2Vu0Uhzaaz36OqBh3Hz9TOUbrBuDz8uh
U/c1vBn21bGG8QXFSUN6sVX6iUXZA0dlmWDdhKFtgHcV3FufzDOI1bJjOlTbiuaLQaWMgyRQ2Dny
3xG9Y1yneSQeyuBkPU+Pst4bQS4keXsoFY3Om4384t4SXeFrLkCnSvieNtOHP5kcPeggztgVih+J
XK7mS0xaj0SuntaO8AwrHmhEX+Sh83ynRkY0pttLBLxhwm9X4cpfsVxke4+sasuGSRdKCtS4KvIg
gBIM9DDqxE5jvFydkVOjyuhvK9F7NrUKM2KxRU/p1n93CgjLFxQImLI+Nifz+gOWzl4VKeADEzt/
FYkNk0lW8OxD781jNQO1ftGaVlP8gFzhZp5fa47xasPkV5RPuBJ+FMd2SNXwWGncX0vXU++bZJO6
+mX31vM5VH4sY13uPxX8AShVvr+VJBELxLnHCa8W3hzYley80sXbSZzQSQXY96UFH5fY1k8xMUIA
b4QFqsFOnjzjbxkv+1eIKdZY/UY5CL4Jj+M5ucrHeNR5Df2iZVZ/crOuPX8GYUj1ZveA2XbmfLRj
b83uniw01W63KCjCjjqlil7QBiOBp0s2WFXkZrMsOSwzTvQXCC5i5eZvFn22V7Ksta48BRSIOh/5
RSKrsK76zxR4D5lVZzw7ZGOGo1Ef8hXb2vF2zWGj63Ma7tykmtHtwlgnU3J/OvJXKwuz5o6SrYUJ
bdHJIz7pIpvAkPMLNOAgiGa9EzntE6MP6ACslJ0zMFdyFnCYc5Yv2s4elgypIPlfXAWRVJodaZT9
mjIS0o/c7iF0CSmG//qwA3kPtt9zLJSxwPH0UZvjyozmh2S582gm61QJU4L4+8mi91gHLP33gmVd
RwxCaybW3FUjUeznqmieYgq/GRTBBoAUq2Dhnud46S63AsFyWZMJMY80af+GYimHeIZAJv96Y5z7
m0NoOmcbWXh3XbnjhUGYIXVHSwGsiKjoQwulCkpWG19FFmyXAcbDl/Q1gI60Wa4jtUJtEVMQEEn1
jTDGgddAPBmpeK0zAIrh+liaOtQEH19eD+wYzkhPkrCqi7dABPJXL6w5cMgPMb0tHgW6RHUxES5r
tXghn2DoB1FCTFbNGdKzN3ddaEQxdbQ15GAx++KcR+Qv43sYBXJ1smytJhfzvvsMYhs3u6Bri0J+
XDLORiTyXqGJ7ULXgO9aVIxwsPcxqM6C5WTqSqfNnn7F678Ar66uRqToXGPt5118SJS1qkZz4mF5
1NEHgv40D2il6B2DvcpirHuOJE68WzBcwONL6BF37i8EjH5wb42RYiMZudcegEuBicOPQSbeUYN9
OlCUMC44bC/cLp8qOsvOCvVSro4CmvnqzHHaE9w3DnvjjqAHkLptuWbz4vmjNdLi5X09al6eIMyJ
fGXWHfUbdWlyOAya09V25zYyDWX+3XLnzWtBbAhzBtXNbj/lo9E2C9wK8Lmf1a1cS9Bx44BjrodN
o7fF9I2aR1XchbWDfextnKKTqel39iXa99AaaBwkbHhzQ2IoheSvCAhFMQE4qcMtPYJM38VR+4/l
SeqHHfDzc5lyL30L1VK1D+mR1vEZbHmuT/qDcPTutsTWgz1+AGPxPIPwGDpACM51QQ16HOc2+MrN
nMtOcmFneqDGHdgOlYbzXfkBaAKJ6PTQGBTmVEr1e45QElGrhplhE6f0w3TIsC1KOtE5s8TTou0F
6W9odjtxIYCILi391q1GlKBW7oysgeRjDeXm87pUCjRG7/DgEKKX/GytAYlX17/dL1HKr1PAVl1o
FoYrZ/BTSt3DsacB4jR6w6R+cpHOFMXW7B+9uHfwmiUKbGOj+T6ixSFteoYOinRoPxqgPnR6J6i8
ZywPzJWZSvc0aL9gOr9IlYYTiKIAgJKZg0hhJUNGpfLZRHV08Lq6qob8HoTkryhYWlDm+1fXlBZa
Sx0Uj8w6GS2EsIMv3IJzcdCtX5K9co6mrEmAFciJ76J+ot0mhEfz/wYjO/gfDTJplR6hj0+4y+jc
GNmNZNz6XNdS4h3uHR3TUlv8i3RbtJCpLcsD8Hyf99nS6bTtuo/MovKQ+8jz0bDpk+WHzEBmAw3X
eKdY6JBP60yP+/Kdzm/pP+4n2dlY1kvzLhDCc1XFqHPxxliY8lbLEEH7NeKJiMw3r3ojodCzRW3d
FwBgK771UlXW0wJShHpqJPiKSt5FmXqn14jqTsIzrnMQ8sdCwTa3QosdKXuq/3VZaFz9Ms7vxU3J
43l5Vc3g5z6J1eDsqbmQlHz+NntDa5RSGpRyrZFnoD87BEQBCRRD1vImlmBWLmOLZOj+T1ZFrc36
D7cJwYTPCmrynYZY3dH8jXZmb3C3cbrEa65FESrhCW+sPlND7FySN71R9ISbaHu9cZHKYY5Acof9
eiNqfdFE8yME01uZdguUKy3zShsn3KAlzB+FZ3Ah5rx2/UOc4FxLRc4+niDEK+GE120jMOzW6rLj
1i03tMgGmGbJWM3xSRO36yMnWlzxz3amwdDf+20927twR02AZwRoiNGMVS9fdPQf79K7cq/jkeC9
S90kbydvTfGx03OcCZzrpbrHlZZNc8BQvdk+3V+TfGqMOnYQpTP7J2EWj+4/XfqJpTkcAaBmKr/A
8CWOyLJWYIYspYAeR5yR/SnRDejozTbddehdXQoUOX9UDmCv2i6eQu/p891R4KwYloEr5dePmVdZ
N7MWhVkawFg/hM2uhvCBdmlNkSCTsoQ6O1eOUfeKkqTsgWh6XmNk74/LtgxedcatNsWOibZGEXJy
OoqTRSc4bqnv/SB+O99LRZjPwt+7h/ABVCEJSyXRwIF9O+GRvvd2p5+vX0pnfgFrrLda2pdXePfH
wbR0WfEEqhF+ocvsQdph55mAm8x4W1aRQBs3C5h3YniRPGrg5sX7lloFCYrNcbUimxrvpDohpiF1
13hE1EJoc9n4ErvhOKqSWmBywQgu66I7ya3aILYHY3mUwwumk6cO1hzeT2M4ziExu4gjj2icmTcS
Civ5D1RrYfbNVguigWMkAIhHpz6KtxZN5DZgNj7jVgcF8bJjPxJkZAM2uKF4TFtELZuDKOEa0YoV
VdD66LBhbCwgwXvC7KQt8weCJd/tD4JSiKKHQm7r2woQD1cSWKKMAwCsdOtdFmWJ+xqqBSdM3EP3
7qB5XRaCL4+GvlPwBBB2L3rUm5DaxbLvi4yHeW/N0jA8t9LKwMC22pzvG0xMWdubTtZ+I2fj1dnz
7cssDRHVD9SMnJG1sirczvL2Jet87/tYOin+P080XgLIpgxaQy/CE/DvZr4i1yM6XhA0DL3aNy35
EJwBtY1MvikKXjAnGk7aBXfnazLe/+QXVXwJWQE/i9nl3/fXRTpWsSOHGyFQ9rfq/I7B6mBjVNDH
ftLw4Yl1CXez7YrpdBc9AsJD0hEYCzcxVyxZhjRizjG+L3cTLQJHpUP7KupuaT7v+2K87l4IW9fU
1HFwZbViCiGh49KwL+6juS31h0DNz0O1osF67lck6xfNAJ0PC6bAYZwmZlvAb6aGfvelDAQ6SarG
H/ceRdMA1Fb1jdgcWjZxEMdkWXr8Chwv3iomujQVvHhUbwG6Y+S9lnWbUi6X7ZhnjOgqADuUE22R
wOkEp5whuYhQggfnpxk9IEGpByU4uuZUCF82pUIwUeUYOBXsMQfNdO3arhIm5ma8im4gfcX54/Gk
odn2gn+Fk5N5vm/BcwWJdhkS2AwDycJjmescKr6yHOptnyXuy6fmx6NJId3cfvpEAqjxuUAo7Crh
0YdO2vhxG9Csn4LC2l7mguddr5dOv/ykH+xAJ9tqZLN/84slspayvay4nKl0II0xLH7p5KEKQ+uq
ERfXr8iYW8GZsL6y8jzeq2VP+ydqkyI6SP0Ju1ruSB5OFxwEYZF9riko8Mxh7oM9zxbZpX0r27Yo
U7qDSjxxl04+O3P6FZ0hVHvUMmBMW5GduloKecaSdssb+oVdZqJ9bL+Jwf369FCvfEzMy3ubXN2Z
Qbyc/ioCH117DKjFi4zB4A4lvtXLABsmzAPW9kUc/jgI2xKEkXZ2dMg21mhHRzQucq+pxGhNDs/D
btdhmvYeh2ViSn/mFUZ3Aebb3iZviM1/Ba48sQmAzDHijwnLn23g/nEz9XjASHnVq8fvrTPGA5jF
IA6icBvNoAe9Xq8UhMSughJwRY+5OEt4g7FpbyinZXBWLvmsaPya/fEx1EAbDnfsMi29lvFf6kTS
o6pkoD6DSOq4kUQCENuxSEwx2fX6QZmnlUFzZY8pdr7Awl/aTAKXd6d5VL3mvOe7uGg0qU3ZFyF9
G+yrqxsavcOchEXzVLf8o7O6y5rUlQ70bEMx1h/iYCT4DxjVUiK7LIgq38jT1u/PdFMwzhaC2NS1
Oszf0qvjesRKiC1MUYX3xoJFjTb07cwNTDwQm9mI4maWSIqY/othssy0M/DGwzavVH3kGLSqgq55
Or9OZlE+skZPc4HJlhbbsJMQtwkmHNyAhzcArDiL6HvxiHeJvGDowE7qnE7waqWnEqXZdnFu91Ul
7XjsQSZTAh/+8hKAdyWVF41mYwfkKcw2sGVxPpTH5fxA/q1do4guAKRa/fap2eP/pKSJQBkB1piB
vP99qAMa9TjjKfFEFBFrpdo4nh4MNnvkBRemGPM+NbRtOBbIr4LctSy6paemdtMKqHfJiyWFFeTM
PsclVniw3HzfRJpuGuAq4Jk7UMU1HBHkSL/ExmN6hV1cY0E7aBSxawfTfm1eJShwT2w3iqzlQZwq
ZumvVFrWUHeHd9Xob+fEQO41e6WlvcHG81ErIvFwr0Rb5bj8Npb9ftxQlu1iicdzyRz689qGgrjk
JdQ+CqIoC+rDOj3tHIyQC2fFQS0Z2LtC9jLxJVXtq/W6Tle3uHSmioP1pZ3ZTm6On+M1jbjCt0tP
YfVGFEAZaUQ6M3+INS6CxtAafUWlHvaBvAIvvrhDmQ8etI+Hx/SB4/TLkJbaQwv2S3uyUNGkXwSl
kvveP7M6moJN5i5xq7+aAlseLR5BvrDOssnQ+wGyyWlhc6crZhV62ua5CVp1J8MplQfhb0MWrG5h
XOzhgXkjxwePkDPdGCztzOhbDl0xJgl5t4bYvs2sxC5NclxW4c3KDUU+XXRGFBGWZWYr3tzN1WWt
c9A8ixSPKInAvxZQcWUCGJJq1kPcOxfuNbU/AVD7Sp2Po3t2nYxwp8ubqWizcGHepM1ccStMV/hx
of39Boow+NjF6gUytdPIeCgumjSYGvMQzxi5ZcVmv4KzJLtFaDXYzByuT/E0YYiruEUTH8bRKPNi
0wQ+ccPvR+0lXKqRzTpHUk2tu4xRTliC11kst2tPeTc4jvTOWCruNN4QmwdIAHRn4TevF0riABfj
KVrPHDV5DstUjhDbzupgU01KRqStRfipuJSi8QxnzP8xKYcxyTAX9xuXJj+i3r0aW33tEuH2lSke
U8n3QRXBhaCKNGCa1UoqG1ilyESFbRnib/iYvQs0j9li8pjISVjD/qoL+pV6fS/c9VJyApZk1ViY
sYOY56BDLWtln9sGovfbJMTNYCxem9+zco0EKsgfwEYauuXZBnJTdYJ7JW6/P46GPWXz0P5Ay8pN
k1NK3tYgNNGQjy0qjJ8pPPDzhFsTWkVR/GB3lXcs4I65jakm2XGjIPTiaStIpHViNg20OnQpt1NL
R9Vpc0skNhTong4t3cJucarbm9ETDq05lo9b3xfRN+GhimBrBfpWTqsmybuZ1Tnf3F+0dRvdatBe
+KOom+WSyPZbQOPX4uSVYfT5ipZ70qmTsDcdm4SP8ozg7osuuf57PRPXtlLc2ugrw9xE2ikZNxN9
bCBWXBlw/abuurB/Q9xuPNicnmc32WvQSV9cIwfbWjUvdbGB0nskoNsIYZpX6ivBbXBg0VPmDyk8
4x00ePjqhNSZYlxVeLUZLrsSAv+T6Ray1pMop2aUdFM4w9RcRusjbOzexzSX7PpPVZsRzkj6LPSf
T5PsVykSYxqRQWJNJkK8CyMaOk84PCPLDRW1hESTGd20snrAc23li36DXZzSrvEOCnEQTvlHo1il
DxZQJMdYop2WN5bPKncSCJeGQ56gWUucAvlRC3+jy5La7pcyYzbQ64kuWUPXp3CytE2Kz3qb6j+W
4GTubZillaoe7eWAbHa/a66kVTPekZlwz8hBHgvK6BgtpTOVzT3eijAacPMxFv78ZcSrq0iiC8Vl
zg4qq5MI7DNvWUg7PE86C3tZZ3QqT1cccZynmdgJX3qz56v7lfnFEECbMtBIAx9AX/2rcLO1U9WD
j4/bAjRomNL4JLW5uml5RhIRFvhB4XaRTVtuE74nzPlcjP7RsIxpkIgyqwo6ldyBwXZe+Eq/T+fy
Lxpj7yy45/0VlfCbEq8cfEL9MA0kcwTveOR96lLSj1KsSbcDb0i2IJREAzMyTcHs4D2mGppkjc6a
jfRnb6A4h+o6R9k7uU0bauokxUpfjeR3oo7EYfIeIeXJIjwa3UG9Q+nwQXWb0gJoRrT4QUC8mzau
5kRGLaXq2x6D0LSAcGY5Cm5z2Y8znLAHZV+4uQmMBtz/wcd64OIl1+DM8iwX8/piuC175k587du2
AA3MIKH+V46jVTtBfzqGzBxFKg7AGww44e0aTjynUBIfrFTUsICsUkvf3VWLzlWc6+w1rgsJDVqj
LW5BRkB7/ToysZ00NgYSip+GshtloeH00kFkzZW+tSXZ35s1GoKXrbv6gajcL6y/7Y50WtUgbv52
CXxSdEDnsEQh3ZLWNYvdbj1ZQVrePxu2d2vh2CGy4TdAhwPsr/Fg4P3bSIfb8GYCD45byATomGmN
wraDhgyZqMfYfvNE4UTw1qWF1wLQBn+duGDIAf3tAi1Y9hRx/nETzVX/c7ea4sB9/xucu/QynHY3
1gm9x8dAk3+DlHZHSfBNw2hXHeLZaCJ1m4y13YXWAYMSJQJ9tVUArAmK3N+sJf5d0JFJ+uH3lvK3
agS8inH8xEMS6tLZKKKlrSgktt2DgjtCtvD+PwA9MkzqPzdoDIQhxTFtrleCfZwTkyWXEDWldLvD
hmOzbqSdSU7IQ3eWbZVEHFg5HBGlXkl4FJbSvdRfDK7WoBUP4IDy4pD9OPbOgU7cqCcwkgztjecA
8vV16nXcPx+ebLsdsjQVVTjH64lja6/PtGQD7st0Wxasz021sNCK9i1IMMtpk074XuVqcqwEUL4t
wBx2Md0/uDPsour7+3DiqZoZ7LCzS+mnONubfpBAKoEwu4tZXWaL4Pq3d6GkS+YEcGPIUrsRlY6s
KEJBwQaJfJ3j480pUrbA5/Bc9IW7/a98U93K5ShHUyQx50OxAfftqd08EGdCify49PuiksJmcX3i
w0A1dMbJKz99TfQzaG+NM5MA0CjWppDm41hhre/3Tpa72m6mViSIzVzvIPEOqUVZTWI2LcH+891f
rVo94jKngAzI+EcbrO+xk062cREX+UQIv9PXIBDr36BWYC4UFWeZmNrm52hxQNHlPmvB2FFWMqEi
hwMcxIUOwFCL5+hEmldkReoF7b1S1hlAlp7FDWmMuE4jIzWu0DBe66sM/7ksIYEE5k4kY6tC+NR9
WGHOe2YsYMSKu4yD18bN72bBfYezLKgMGlLSyHlq5D2NVh+oexDWPUIeUsHoe1X+q+SQerUDXsyt
NEpBX8j8BmLhPT76NcQof50B7OxiukDmgcxIjR0YHajkL+dQ5XpVo4CFjkcqRZ4a3x/LjMFqs4Kf
VfgaPrfJ+PH0XPXLkfWLJ5t025tMkyiLyq6wjnF7HWOds9VynuyztkWS80LdM806320kXcKEVE5Y
xHHY3v5CfTXe+Aps22gpcNzgpJoHNiZKq3IxwWVzThS0X3RM21lackrs/oD5Lzi1EuuuJvv1RLD9
4UeyMTRnkKXBOnlpWJqChOF41ykl9Y2iBiF9Jic93FEjJR6LcUo2Fdpji0XUu/tlGxSO4MVzVoLc
oDxUDnya4/cGA1YKh05cXp8RTEBBFLFlyMJQjhPF7uCE7HBTINVzzen/ZUQjoPrAZgHKKRcvjwYm
LJxdLCnyhAkGwj3Ey69V98zPMTbUxwIodMWW7Ja5pYX5bk7AVO4hr+XwD5yrMuoyjnglPCxckijA
mt45u3gHsBKdjZeMZtgiT+X62f8pbrjwZ+iB1ogV8Z14AJPD/jB+2VattcDqImftl5E6Rj+MAtYT
FwZISkbg9J3LiNEmXfswBFJGEGRDZOGTR8dtd6ykrPygtjAwrIWzfHlGZFzA5xC+kNyUdtc3RHaR
Ma6BdCet419mImXTLLt0as7ByhlGNB3TyPlbSTjZ+XGtRgjkt/aotWTfDGqNGoLpMGRgTUdYuigM
c/I+hlfoOHi7jbBx9L6JgHrNDRlljeYHW57n5YxXfEqyWDQDuA5d0i3q3JHWbRzDaZQZZAq9GvWV
OjN7VrB2+Iy9y8+pLgjBpK9hU8HKtNIfwJtFNxSOiF3pV4v37IHJYeQPzxSVsQcVBf5crH5NbIJz
s6hMMcXM0H0Ak0FBQ7H++me0vsxtiYViu/LOX3oNnIoDAAmWCJtIJ7vuX9AnvmSECEyFHFHob3fC
OsZUQSTPT3W76rw0dvRd+IqGY1kJs6QWCgAK1Sg4PWGuJAkd5R82zu5iu2iemA8xf3kH35Kzdk0w
OquN98RjbG9qmH/sjMUKY9tdrgRGLD6GDEbCriP82QfW/DA0c/wX/qsu7dixSZCUOp//PxzEkl5J
xiK2ZOP8UWxQJ8c/K55/RZYI1zW5eOunPwZwN+QPj3/6g2nV03NsO1b1BQRpHj4eMgUqt9fBnHM+
tOjpE+EfJ5LtkeJ7h7V5zZg3HJm80IfB/iwadL8qKWbE7Wy8ksnEOKgk2dslDFiXRsTHRNJyRwSb
w+SnzMeoaAhcv5HlI44L0GlxKZDguk5c5YpRYTKmVCbzQDUPHLkXyiet+HCv0ZL1gH5u0m9X7CSU
UVMbaXgdsLAmMCCv+19lB0KY9f/s9LmVVOlfvCLnZpm11gfBpaxvZZZ0VIAwyJfXKrOfbXHrjyum
/hMaRjRB4IbCMsZBDrmbpv9bx14VWxPiOO2hai3loxle3KE1hHUuGO/TinMMc8KnJ9yoXTzBIPun
QDbXPJx6La4Yl9vmp4GGMsTk4qmtaI9cWUOPlrgz4cW4FJaIv3avqUfqY4Y514EPrgymsji00pGH
tN8iXXwR0Wd+gdLsXCTj4JCUMeBrNjVemEU9jw8M9rVcriM3kQUuxIUfJRpts4v8AanwQGVvUJ6o
6bXTOVI598k123/DprCWCajxQpaFOMEumSRbiejpsfZxk5gfBiP5ZlzAeyEndoDSoKSmhbOBeefO
C/z/6yjfDzx32DPx/HWIQ4MTL4FGVPkqQix6eFkKk4CEwWNSEqvOVp6dMLZDUa3N4//bEZvHPNfy
28eRiwrkorkhsuPquU5J+Fnjd0K0hqZR08i1ti6+SzOA9sx+3XwQ721r7lexnP20nDHCj+LQsiJi
IJJFlPc+cYjWEibdkdEKclKp0SqAsJD0zDu7UwMjxqatp1A0yj+bP3D01o1sHY3WZbkYY6qRGSr1
yiP4svgQMxSPM5o2hbs2ZagdVWYwTw6qT9d4dlmiZzZEgr2bZuJt3jBxFCP1d1CvLVb9giBoXf6H
taGpTvEynWAjTMhwQHzfyDOQZNN3aVeIubzlMVmtcpZA+86fwe41a5jCO8JHa0B/vT7GUUeiUS82
NR5+uc+KsAaAXV8wBoDiT8Jyuun7wnQ6gVPRv3w0swZe3oaoWpNi9fbpTZ7GHxEcqnDVz36lN9ch
nlW1/2GVWSmLv+t6VS8BmaxyVik74GxCevFDFTekn+bwIp4uHVGnmC9YRgdbxo1S8Qo0qAPFBNU3
8wsxnX3UGMKw7Y7rwkymr7fxbyWyJrBhsGYIo+NVug8wunh5vE2/t78oi96VAiNQUh2A/leuYnU4
0lFtwpObkIoWGiLwpsC956B2LaAflNPmDi6WPwlnNyB95siKC0b6g3/oTLU3m0NfSbZ7wuT9TiAO
WbvcvNhUaizmPsTtBmVf5Ur217XsWgiakpeQv9xa7+aPDeDEv+9Jw1IMzL24dIASopbSsZsZ9ouE
rkjiLp8OLdh28eWtT7KKcyb9lOdIw3cZPIdfbZXmexmkDqbG9f1xjYAigfipEDfqCw6KLQKVY9/n
apmjExnr/NaCZH3uw/iYEtnDs6omaPqvR0SQ4pnX08DN8VeJd1fkUmbO70qPTzX5fYiQjqw5DPHk
bB9wInSxvDmi1CyTLdYslfLW1pPxIPPQ39HVxBuL4ZYElpLJe65RSSMGcEoydY0DIKwmrnGqDGHy
ABVnaFBfSYW1w0VN+D2Xg9K84LHs9yqou1ECM68HN67fEgnX2f8ubuvYT/nPZkCbrUFul5Q5tU/H
iun34MxtS2edZ6OCqnOka4O/hGQvZim7z6soHkRD8Ko7PkyAFQb7BLFC0/p7wLwl7/6OuXnq/Wpu
qekXI1ayLplHDFwzhrahXl64tAqghlDeNy5UNdrEF7fQjucc+YZGyx5umi0TXpUqG8jL60tuPWnq
7uorD/KfnAxF0Jon3dn6tgXwJ40yqelqltvb7KVsNzfstattozYXaCa9UHJPO/2d+cRzVgIDloyF
Qdf5HkQAB1pABkgfMpTemDorfoaF2ffc/X+hfgW5jKoNCQNEMd+W52LHrO937tEUpCbMvZ3TtTzN
XT5v2qMc19mOZ58h15bj2yqa936uOT9TZk/L7/0sW+Gm7kJ1BaqyJ7V+k7JRwQMkCBmZeCtD8lpl
cKo30ug7C2LJCgCNKNBp1SBzx6n4dzA/M2NcGWPismzlMDM8+y44pvDG5Prkl4EvTC5g5ZVbu9xj
KLgOY8u5I0zA1ukfjKaew0DOui366SetrSkwAjePX4nZsYCq+VTArYLGM6/ZNFJpKRK2uva1e2Ga
KM7EcwGOBvy08Xx7siYVq6gkJz6temMfKMtRSPK6SHkzQ2rSGE5lRY6kjfvZrJW3V08XqkL9wMYY
gv/l4fuPmyrgz2wODOcZr3wRizsrYY68gsrBz1sFRWu9+499j2k+S/G/lih0x5nlri6h0FhVc1Hb
5jEEQDnbyrniK51xXQWa33mwPaf8XrHIpfvUMxZytAH8neY5Xsazi17aYOZQj5j+is5qU2esjDKm
YIAWxow724h8ujE8LpZK2Y896SpxI+6pHSF3+U/fmk7ZITqkIlPWXUqKgWdQ4/+9JnLIh+THE+jB
5yIlR71CjZnPevfSpQbJrMK1Riph97cQLasZPBMs9MTR+USImfH4e/VaRlpAeqi+g1C8WdjS2AAJ
tnzxszGAmOcm3M5LSIsy5Qcxb0S8UdXZQVVTvWWRrKV+LLb0Tii9J7es1jbfAE0aQq1oj8qO0WIx
ZGz6HqJLCHvnp/H/0RUGoKFNRp9nDrW62mgxyJbtuyZDvNThmbgxwVH+N85m2nu+Y7rBKCdN4gj8
pqzR2Tcu/tqdlQ/yuWwlVg05Adqbg0Pks4cMOwn35AGiFWWbbC88tqF0iRUsXHCLZkKd/HbTttTE
z+ctOreAwXOalaOd02eaOEeVwhKOrCo2NCR0nTI1jUqtGlmPkFF7UbgtAyj39VujtpR45KJYnKJA
Wt1Ed+6LuVDKxhBdgtD0tl8fpXXJzIrZakBYgEko7qL4G/9K6FMHFsaRmrcM/yBzkah5ry0oyTyR
8XpJIEImv6lfZqt5YxcBano9Ns0PpvEsKWQjaKgogWT6Pq7vN0GGvbQni++v5Tnv1cdwXXOH1nkS
RNuqkQ9HKU+x3mlVRxfWrPSG8OOs6/lZpRPPFYfq6S4rgBaaBSl9+lE034fgQ7NDTRnjRChYn3to
SVBTAkdOfXLvgitrr/exYii+zutpEjQYgWOdeageDH5dAJ3672ALqpZqhk6cC1ypFhC1ahzQQ3H8
R8oJSQIYbB6GhhNzckh6jvGasJ37UtF5ctEOAwftQ1TC31977cQkaVfgCFvcbSFCJ96TGqt2nZFZ
829EM9JG9/NmsPvCRKfZAr1nQEKn90cYuCTYvD20aMLyTM90D+U5gil/JzT1rCYm4XOA/EQaQjnG
sLSJJE0mfS6bdww9vDwgav/odgjnXhM/Vuf9DDt9XaATwA4Kgk4us7aKOq7vLrUGjf6EpPfbM5Li
inbm0wO0keOR55Oqq0ygdtJ7X6XB7MLvlQeVIYbEByZN+hQGgMxgw0Nzg845OrJJb9RbeYMy1P/8
tdEDlWiBFxxalf3aGi4NIyCKp8eWWocBmYeOnc4jWxNPBynPERt+XNgeJ/CDVX0IK2C9k+cC0byR
5uCMK3JIxBIzOgAHqLFdWxMR6kAC3YxMmVdHvnWBtpExnDN5f0dgV7eazXkjIqOETlM5E/HFF5m7
Ijegl+VAk2Q+WJNuB4OVWQiWV5Z+Vo9F3mUrvpMPQuwUTC2fTT0u7tx/D8dG1sO7PczbR4wV4zkY
nRUfsMmiXF/58QATnfmt8LK0Hsbif1Pp4Ltp/Rf64Pn+nsqmVGH8Gojlna8SXVGHINDjJlxQiLN1
npyH4PxAKSDvHa6JzSeU6GaUWMxfkkVOCBzmW2iET44zQtA/iGPNrlxv7zSr0CvIRglTcvcHFtd4
4pluQGbREo7XK8o3OUooiXbjlc1bTwo23Tj3NtzyBbY5z09KR7S04r56GcG8/qhFJFAJo/e6yMQt
ULUtC2EadSKUlnee0CkHejv4o90Zi+WoHKQWknoRcm1P74EoGw1Hb/KKo0LO+3yoFI09QugAuyv1
TRb2UfxoRZxHegxTQHNn8kh90TeRDVoQVBFbZ0u7Qxz7yVS7eZ8iQ/mTCA4+GITXEVH85FvlxE69
8ru1PebRlyHtWPUYKxYkUtfAly8HtGLTt5XF6FWk1Mvg7+ZhDjQtrNnDeBxGoCsq/V1XYHGK+8VJ
iQCO7tUUEi6Ia53PM1Y8NYpyRoLvKg6W8peQxUiAkSjQUtgikbyK7XkTxQZxeQW3QcC7pNjA7cd9
YJIGv+JfIFz3wSE8nFnS7MLUk4xrkpOsm0IzZniW2hlXWaVnD24j2eZRo+CxBMcy41Sy9eLNe1+5
xbawYurWl1JrDgnTwn84x/nlnsdQfZ6xGp+MDiC2bpcixynQK9Mz3exylZlQdA50srllxJPeFalI
DtoDvmC97GMMYr1g8iM9kAZGc4j7MpxOV0wobNZWrOcJymP7uC+5nIoZyRT32ia2cu8/x2bjJcSh
zMrkMig6HJ70EI0xUxqHXht7FRGkt02Hf6j9fglgDD/qjEiHFdvoUTT2S4DxIfkdhDyMlWHMDElB
E+zvo8TgxlEOBWmlCR6pPBrN1Dm5UJv3ESFFCn3a3+AC/PjkJhh0jlSKSGq/aGZEltRRQudQ5ClP
rVU6bArt3M5I8jEIqIN4NCn1L9oAmosCqgjNKkvgyY6iab9rswYFJBcu6DbtJ/dyDwKnvft8oRP3
ridgZhvLa45nMU+KVJSdES3CoI6iM8c3vIfFMfAfRMkf1cAYXO0Tclc6pwz9JSVMB57zH0aO2eII
4fxUMlWrmy43CJqVcC9F8L/TUKXVZNDHjOBk7IkKdAzX8IccgPoV4UCHrAiFkQlyrH9uvkpgRIrx
oIgs31AgkfVwCp9y8o4eGf0PhMR98x62D2ERKGDcJHkuDFWzgU1GUFnF2YhSQzxa9JaiCOk3tIq1
KSyQxnTq1t6+W0mq2FWT+ItBNvjJCY2G2+MYCzUQQCzH9BzujmigAwn88nlpE2JR/p67aoMnlQlZ
sNeXbgUmfhw6OYoj+aVplf9yrQ9yec00khjlsMJf1msceAr+waKNXVV4cEgXKWKmlvzpIG+F0D6b
E2X2Xff1hCN6eznZc0NzUbeUnkeZFuG4wXL7Xk7LZssAXPjfdESBqpnRkFitEcl0ZXZJ8j4QOYOx
ddlE2Ony8YYRIh4EoqN9deM9vjVihV7vZqx15bR1tJqwV+O6MMfncydvKqTcAdMd0OqjGUopGyc0
mOVzrr/+uWdMNkO9MwcUf6BU9pdPX53OfdXRCt7ouVe8YPiJgdkTrCpSIbynQtk7m9kBalxYkhZO
Junez2GE1tpZd5HKHxby25RcEtp1rr8KT+cA+e00FpGgrlJICTRdOJZL7yWtzX/GYqWuHxveBxvE
wNhMAoIOYxd3Aktc3F7/qPYUuZY8aZRcUu9knwdw/FMlr6iCqbkpuO1Mz5B35F3YOGwGKrqprjUB
CkvSoPgnshNh8OIzI8MGY0u905MvqmuAq/DzqKKS8XLr8e0VrKC2M45E+fsKZJOlK9xGDD+Ybdh+
O8e4aUtwSuHbGR5NS9WNzbWIbN5yZ8crNMsUbTXxqtRNm3JGmkS099s5/oOZ4fFKNv+zPR7cp6YT
tawtJUmbt5TcUrvE701oGNrG4Ec2hF+E2zhQpn8WNPu+dZ45J558frOSsuW41k8ECiClMCErjjuJ
OEsLLirpwqLNUVeARfn8sRiW5I3+3myPtJGLZC3KsQ8r/utDrI0jIQLPHwg8/qliE49q6foVkd5K
ZMWMgh6eiNtrnQGQ6Hxcc7WJrLpVmJFWFVDcsY2T9UVOuqfAZ7oQ/u6yQpI7oyvODXpO/6ONhD9l
pDKBs9eWDZbgvqpTRAls3NhuA67dUQeNtZxZId3S7J5hK4BUtWuBbDe8CrKGDgMD+YxQY/CuzyoJ
5vDUAUo73eDhuJdPZIWhJwyT/bKVPExTgfNoKfpkWV7IS41VPSYqpcwcIobL8JImBe3L2T3Bre4e
NO7ksI7xLBS4IPJt7/FbJi/Usq6wQm50gtG0wCTcRS54fhh9Fz6pEw5CkAGGZbGNILqPRS9TR4bb
0N7f1k52ng0p+6BgkWgzid+ftefpQwHjoiUvk8lURYYHgwNw4+Q0EY2qnehAhqaMolk6xbql2Ium
4SaKmvty+bcxlDCNmeN25KynDST1rUI2+eA8gndDwwzS8h7B2iVASOSAvF2bGxs3/49YRU2X3g/E
lbn0+gy6/mrKAeVHdTrf36ScI4xelAjDgGABsZon4YNdi0v8jxSy4qpzJlibZUpZaLEqpgEMswN4
AL8HsyUPnXBqUk3DuSDEqG+VHcCN4CayVVnAl7bOLDx17oGt8LdoEKOY0JWMVmndTkZ81uiunh7Q
SzXd0CPCiVgtE+MnurDAUPv6HrOsPFWJf6UCNGg91DSvvrTvV0IcUupVlPH+nCKYhEjU35p4fiX+
ndaKyOEgvqbOWUVPl4ezQIhSSY+Y/EVqdtjtwo/5tO/XYW9Mw8AcYZfQjqI4lb0JnirV4H2e3QdC
9h9ZNQlTI8hQde8VcfuSGXzX4ZQHgqE1Rzi03DkPwkbCJYteVXPnU1JsgSx0Vk/pkKC9/JnwEvk+
cc2XshkWZlivSXRxJtOHrGwZtC4og/rT975Y29n6Pqt/jtT2dFHAviDE7jBAXZ/y+pQA+k41Bxlu
Qp/qCoSbGTH9xmvMjdypkzfvroxnGgHvSr+kidudumRh/VbVbS4KVbPyqmviV8k4+tjK+55A5IoU
pmSleKdcqE0/wW08vBZ8GCw4SiCVtcXnx6tNF331sOsLGcACrxy91Fqgi162CzxalcmHyt8Xh9yG
44ia+EfiHhOMe/8Cl53XFxRHpkiKlSyKvEegL14iF/nPIAV2T+tNIyv2xEzasGOm/jjJKYw6oZjk
U0qqzyAgDDPgi22jJMX4qAZJRUoTSD0mRhXTML3IBr8Sidv6XyDp32YGMKOt8L1KAFHaGQaeolOH
UeE1ttb75FFTytWG5n6kvrVriovFcnpWjR36jcx/Z+/JfqO22w1ZKMdWeHCuCdOJNQoBRY20JqlR
XClb8D08SzWdLrbZHoxyRqMgYhfN+OpBi7NJmgTLqXl7BXnwh7kIDERod0oK7V4b/3bmPbsMbDl3
eYumQowa+WNbPFtUfxTc5tu3n72UA+99JAIav191Nvj6okZzsVyiA4XTBLuvEtf/80G37Fg1fR6r
UpH5mU1ZxoFlAZG9RJUlUtHIa2BgcwEMI02EguS+mrDw28BqmK61MnMAptG5pLDcLm3Jlppw+GCt
Xz89JNInsLJS72mdfcAdni8xegaxtWqp6xgUF7ns5LD+SawubgreqOCEi0imnX3rqmxUA7lKfF05
/VoamXhiWob8YSSK6YCZFG8U1wykfjAac/x2Lx8fXtleh072pnqkRn8my1F+jMQRje7so6zGUe1i
51ysL17mA7PLRJVBWqsUpnyPQSpanlyNyTXhFmtzR5YUYMvPJ6upxoGiqwtP4hWR4N82o1RasK8G
Qj/vRXDd3KMkoOhIAQVNb8R9nBwGCuERfah8Gf3bjSpeYxAcWLAUkn0pfURRQHlJDr6OUJJqQvzz
qcNJAX+V9hv0JhBVSlaHgFiTKL6GJGCQuF1ZOmfqPvqljJy3tqlCvlSaxLeyzKcT2CZhHtFpd8RA
szMiYv8YoP2/FU/NL237twSzyXAGHad7ytdzjRXjmRZpBwuBmS3nurDuuSxYMfjQYO5c7UZn6fY2
b1S66V4kf9H+GRyRX6TOM41SuVjYjbqpoqqzvQh4NXgIVN4nI1G6Doe1CQd7CsJiTOrllrhqVpqk
hGDfGMHuuMZUKu7LjqQ6fpWtpgMsTVpgr4FhJTyKI+T1QOvYyStnhMotw9HfI+MnouDf1vbNjjGd
AzpRJzubzFf6ubI2+bj1HJE0Olsv8oO2bOnffKoB/zV7sXbgnHBopDbZXi6esdUG4lQ5eE5LEGP6
LtVubyB/K1vgjP/FrVEJGgOvfvBuBUb6q8ukC+5M1i05BQviq+0+WEy0s3x9RQhr2lp6HJd/hRvv
8HPbMVjAcXUmYXuYPaFuKHzwh+W5lbsuPpxUWF9oFBTfCCsRvVXbncU2H4aa5sIDwXs172JzI+o6
7A2/XW3H5p+L+qENzBPKKKxliGrHirF3HLNG5tjbVXIracdx9B7VBzcMdyr0kHB5eGI7r7jc/SAw
NQi4AmU0Y1GBBqzqlTEXRnYQk2Dk+0ruEJOH18vRBNX7tEg+KOHTaZlyn5XODzsALI4jSr6v9t5s
nj5/9UYkikdDyUZRucWsRzIp+yVsGmjUvmix/Mu9yS0kHpm18sq6cCkfl3hHyeXIyZApeoE1Qyml
94flk0AQGJ6MRkaW0itaaPw3bhxbrhu765UqbmrZJkOQlensGmlpEkvkC1AGMz2Hjv9MfyqD3Qdr
+1S1ro1sQjzEXwOsyBkZGTA2iyRZSwWOW5k1fvD5Pzd60mJyLiOmDcdu98mugBEl4FGE7v/5+E/X
YXpwwOc8OKdu0fgbXlKYiL1Hxs+T9GzC6ZnQ3EXW9mNasGFlFV0b9jKb+OGEtrRiIJtBdj9lpDCy
oTeuJaw7O3CBUZwwZfn26bvJnl2E5dhGtvDGT7wUUtYuRtGOAMZzuE8QUfr6xkrkGINgum7l+S+B
wIZCCdLxw78qXimfEudszLIsu5tfFkguS0Hh5b+P8fUHkcd98i9SsjfJAEiozyIMbqUaDL1BeRDd
rIORyTBmJPaIDh4nX1uFVhvgIlWjTBdfxi9fX23xrrpz6XCrHvkItV53HPTFPamuMnO4SWcPLUbV
9Kf8Isgwaz01iQpxgQAKtVZhevMK59Gr8lBOF4WgbUgzG2EeMMp8oQI5EeQePeZw9btSTKDVXnqa
ZUH6Nb/rIg7aIWYrsIom6Y24Xh3mkUt62mr5CAdDrscOh9NC0pXFP6HJTkU/w1Xtdt0JFB6lonVS
Jyafq0qov5xkwiUvXlf6yYQvzOFmvk5ohJiA1XqwaChblPWzonTrwmVzcfWdUWrRntW+tuklU4R1
unSl3biVohFthYOMcERC06aj3vRMFmzHM5C+L5fyiiOeFZFRALqL4MUbSfRsHgtHuTZkgPtCvIYQ
4TQ+vHh/0aelcrLzWw8dgzbJt0VOVz1vcpC5XYZRTLdDce7Fl9837N5s9mQ9T9puGYRXY6ANOkzi
nv0HrW+vLU5R0Dl3Dl+65lTNY+ANg2NPniTTVKmgDvCNlgXd5kbfRLYue37lXiBQakUc8FuD8GN4
kh75PynuX/9j7EredFFtpz9jn7fdkkBBj3cBM7qaDi6BEhiDgjjugUo1abooFeMhJ65Ypps9yZ7n
6gwOHsfSLEvJZgCnzNninGMRkQQwQ8Pdi1D5uAxFtzirgcJPY4r964btMCq7s4lVvKvoYSkUV4+U
qsGMFzw7mb3nlxZRXsb7z+sYPbruLGyYZLPx1SJWXtoAIjZCVAsxsB3Ft4t9mP65WCez2r2ztUQI
pE1RG62BoccqSRmy/LqCOZPs+Io+dUxjix/roODmqA5MoyCsvKszVuyMTrbZINmPpM79+WBk3SEv
nnvbzqswyja3GCxIcWhzlSHHtPXgTsmOVcQ6nviJF+0pmO3iQFXqP9pCcAj684tawQVDGxk59nQE
GMohVZk5Zf4fJJlIP0q7/xY7IgUvsPNaLTRWiQZivmcJ3px2sd+yVXi6RIoOONllEw2LP6dadMLv
UdsHoOJ3C8/hrl+qzNgRiC3/DriQ9BZjO0Qg2kcytfNK1DkD/hlYeMHMaVdKARBAdXUVeYM0cT8h
BeTNiiy0zri/H7PosAaHNFEutqxYnhh8Via1L2iiJQAdUbF5+93rC8W5P2JneoBqIJji4FK3xesf
Jrwq4CoexOcebTtb0Hq1qopYxmdnuXeBX7hSFnAe2kwoSobTCw62YfM/eRDBHLOGNXN4PprUto1B
FcL+dpdRaUgdCRQYONWVOsfrG784Zpsx0706IzOj7rYr4FqBVHrtJse+OykqhR4eetYbdufLskgx
XmKdBFv89u71/2miev9K9y49fPXUFg23Tec91zjSy8zSsHq2auV9YjjCMhIxOd8JjQF9q1MqQ/ye
KKUKa0nc88+Rb3viJfdbtbfbHI1n+0auPEHrCkjQ1nBI9n6muM/u/+y+w3ij6CbyW1+euchf3Du8
YPt+nTTZAMFFI53noWOb2pALeIQoc23lw6YqapMQXWLUiD4Tg3aFBmkDlysFxlXDPVAvIyXsedXx
zpmEBSDLFmtslIvGVbhFjvTic6jjU+yWBwba+zEjZGvaNDbeZeTOl+z3obIKNmc8THcVgEu1g5L9
dDSCkGbYlsAy8dR5hUhgxbrTdJkV7JNCD+OtJhg77mbrMkosigDGmGSnuoeuokn0lZttxnzof/Il
UMjSxmh9HdPHi9ENyQ3kqMllNzXDDJIWPsCow9wLxWazivQGxpVouQmrKkvcp1IthaJMQAlxQM8x
jNDQhtWmUVUBSBcVRPMN0Muknx6NkXfxLpeCDzIeY4UWkTIMUdPP/azMkX84/2YRb0PJkDljmRc1
j2R+x7xugTCgGVyUO1QzUO7QIamgUK9fuy4McYLdldPhFPrarBQu3MO1eyYqyPvaqmQXCSvFVQVf
50ZpBfUtq8qGKHPh5SDo51fou9fElbU6ENZ2YShbNG9gKWEXQUWNhilFQnqlluQ2eIpfYVFWWlt3
C9At9S5iQsB71C5PllZWVyNcpU7iqdmT6RDX3JUO1MRyXK0xBaCq9ihUrEbBTw1odIR32VQI6e8S
sikPPa2nSPlbwfPDgSXyXjGHXCsazBliC9a4THA5Bk4ONR3QwDG101uJm/Og8yjZRwc4TVOepaFd
w+c5JS/S96EYzimMm8URRNmtI8bTZkm1nlGqDBnNkd3PSeP6/7EJCe5fzFpHvSoePqLIZI0rdU7T
6QMGlpte4V4npCB70tYLT2hlCFgd35Q5GfTYSzvheorG6uxRlybWKQBhv9hP3YjIg942ktMFJ6YF
Cy7xgciLzzycZPEbq4V2HWZEONfAGESxdmvNHGGEZ0TCIlQfFz0uLhdO/ujw1RD4yLXrnNEm67UC
tUxKHN2PWFL2GkElz1O3YOKcagVhn/Xqie/6JjZcP3zZ/T91dmvKuITGoSUI+Ll0NBwRQTf8DS5Z
dpjGb5snJDgWmwUnN9hN5r10vWB9ajfg+SbZshA3mrKDRFgj1NyPDZz+6nkgoyrE6ONg5Q0WP7ZV
9onXbOsaRyvPw1xZG2kPAEpDuGoSjQ0HXbfSW46CNYjKbhCPiRkyzV6VqU/4BToFELj+/GZgOj4G
0LpjXASN2KK96tkXnVszcBSI6UluHIsbVrbN4CCRHy4gJ5gDKrhs8NTOPRziysc8DVBTd0QpAww4
K5KFtGy1trYKKG8AF0JWF82cFoFKm9JdYqHYcJfK8kA/pNsSt3j8UdW2tF1Ty3FNvwMkOiCtiw/3
8tczuNUHi6aC1vUYDUv9b/6RnbEmUNvrI/3MXz4tOCoWwlNSlai7njiP1Fe8I/twxZ2Ng9IlbFTU
+w0FziZ/PsnEVPzpvEFp6KdUfS6rWyVC89mMMaBz0dCI2vLt7F9scAVDs/QgJLhzsnqHGLmOtnmY
2kIYfAbH5EnDX2jfVvMgkMyoC8wNZDdjHcjeiSQM12+eePtKiqldlq3DN3qehxZxrLN2FWPcFETh
MF641dciAZbcOFevSXK4VMLQEAyIVERSKcgtS6F+GIx++5tyejAbH/43kldqsMkg6tLGrRizlSlP
XU4DtJHcj4uRYobjbxlYCpcAh5YgywJXq2+huwXONRK28MPZmagmhMfBsb9s/e+R3Idy3SrzRQVv
Y3ieVdBVE7U/pnVQ2bGHTpCb6hYDqXJjNFz5LWZ/fUAbeks4OhAGcT1ji98Bedtpb8XaLJzL076S
oCBLyAOoAy9ExfDPYsiuO76mgvPPOKZ5DfchEni8jfM/JOWZDG+K+fuYnvpIkg1yrF+gzFUZONdX
414x5IlPQ3YSmDLVRxhfdq/6fyYU51EKYFPvAEe1241Fi7vzIcSoJfv+EWCA+H6i55yA5Zu22KGW
o8gS1KWyhtG8P/0onaWNks3YLvVgZ3szspCi6ZKP0RzGeFUItuj2+3DMs0VtCplJpDlSdL788SRb
csPnsGNGqljIMbtqC5G/mErA71HpJEZRY6C70mE71FBcZ0fjEywAxlUbCKTsv8pqsQYs5O/ISQ3Z
3622CE2MvlnVUBLNQ3cLGTnu+OW7S5g7yzswSHcLLwnVqaB6/SrEwwcoejOYQlCXwlsqSgS6Vnr7
pkLMtRyGY40+WA0v6528viuPt+kZ1Hhyk+JsPF923pK8hj8bsQV7Zfm3m/YZlFTSGXhgDB5oeb/P
6QH3WAAB4ExWavcuuQCvTK1Zde5H3PrVOJHfGx8+1Z6yrdjNiT6B5RBKkhNUcLc28VHOa4PPGz2J
0dH/2c42MNtKpSnN6TwP3KQLGYWiYOz7seaIUBcwXSrHXzAgsEz7KI4KIHrGm3Q79GnebSXgekR5
esgmawgrxu5opyNRbkkDi1kLmBaoDCOPJJhAISCHkL2fNy1b3gC7BFho6GYVUjcwWmj2OD/CrU1x
jsKfQblbefIzcj76mmjGRNQEL1/SfLau+AI4Q+T2AxuRso7jFMIsCX4Ty1idSlAXJjQFj3wNoJic
78rQLYrGkZGmaJqRlRJBzkrrQpsBfBVn5f/V6sD2MF50RwvibJTaurmw0GZlZJjiahnk0MzvFaJv
BeY6uN6Y6e4XvbgSiN1Se8todLA7e0f3SOROnFtqEMmgaDCWX9BzDp7Psq9GE1dKtVYdoIpJ3hcf
bTYY+gGlqmTDqGea9aIDY+Q2M0wyPyH8l4ioQgHZMXoeEVic7ZJBGJaC4Jva0v4je3QiIBnvpdyk
or2HNVOGEm4j72fv4Zrai3ZLo4hSparyRA8ZHvUl5uuDJUwxJyu6CXBuFNaUs41JES9D1wqK2N5H
ZWdpFxFDpJwrqUpcwNao8OwvQpzjdoZT7ZgFONE5pYHvO+lU/Cky0l6HW/T7DNxxx4L47aa1lQee
kZR6rLehwxq53Ii/FRTIkMvDxCUH+Sgb5dDSFNRBEiOmeDTe2NhW5gtgBWkkKwW80VLaqJ2AWUjY
UCpDeXbIh0jPstx81ghyx5tVy5pwD7JjVlLVUwNOqtqEzGC2GNx8LqvN09HiYvW8zZAxUAtgdNsz
5u8OgQRQNDUMtPyBZG4Z+8hIMZtupEHaRYdzDaBGBH8xUvtVq7mbBHPIkMu107tuywBSfmS6KLBy
mslGPr4ShHbxfEJ7WROKDfFXZ3fX+tmRvgelR2OZu+w/36a1yvIp8GMXIiyUP1ozUYdLswKkjHMZ
UPx+SB17fUNPIyM5P8iJ3KzdGOdticot6QfH2q6DKkuc+iRgLus9fObi3xStSzfT/QJgP7LkRtE4
nYoxJSEFLIMu7G2lm44zclkU6atk/C9PT2IsaQNZItS7MTQcLGNzgLTWKezlVQ60NVsaDbT+EoM3
tOknB4r8OP6RwVFHpLiI9m5pmtp2X9qtfrA/Et+hcs12ElawPbXH9fT3iqYictGGH2qPimEfzbnx
Vl0e7uySvXDlWddESXk84CJdbM3lv//4fnBkXyX2JeYH1ne1hAwjNxjIrC4qmAyG49qBItr+hlyt
G71unEZDicZ6RosvFd+roLFVAHezCx4vur8GYu1/Q+3JI7Ps5cx3tuvXe5kf4GSwmSA4PtI5S6ZU
KAU94TvWuWTDsDh/dtnhpXPKQmhGZD5gMUKIkSosO4rtphvmar9VnqPXUXa7XVPJbxBWPo5KoHng
23cNizhgL2aZ6BDn2PD6PBtGay6fN9pHHM5+DDqDWM/K5apVDYxQ7phCpvuDm5pFamkhV1fTRY4i
9cjvy/w1GBz1IW7ixiQgApbcnvp9j6xWZ57gK+OBxKosacFJ98RzvLuZ3r8SrEYWr3vzDTq2hSDB
F967dsC+aRauT6LgghI00wOQHfGTfm/aaY7jBgZvJBoQ+MfyBNkHN4hcYM5To22rrTHy9hopP4+Y
lVa+qoNnxrgCCYcDeECV+vnGZO3MXciBhQO+YHWFGBYDFP5h5IYuuWq40qTbu5C5/fov+o55KzHq
oU+7NFhImxoVlyfIu2JCSGS+3O5Dh4D9LgkJ4+lRcvWBWbLM5Y/TZqw0gWbhrUxXCfozAlhEUPz8
1Tn+fPcfOWXjPYsd8idv0pBEZpQD+1kJTUJkmV2TkqJq5oQe4t9X/GwiCDYNaZZiggro2XeeqiIg
zdPhnc22b5HQGKJCVeR/ST4WgbuNNXO3CMmCRv1PnoO1wHiT4OEb00cnJFTxSv+mM9cJvJIDaEMQ
48KUEOYcnk6pANR9EE/mQX3tjWcy7XCcXMVT5CmcnirrhvhWlgBIklW6zCD76uo8Jvdd71Zin2DL
DUpqY05TOK5YfeUG68axBEE/sSobpRakuxro7dtiBQ9lw7FfEsiCAoUQOuAnE8DwuB9pOMF/dgG/
Ev/9MXHsVusNTK9pw6fP6MGWaRBdzmd4UfgAUSeXppvfekqQhHhLxaZD9ElFz+WQ/T5QSeqVPMog
gXrDSUTDp41FVjzhIRc9+lsbG7HE+ajttcFbp/lUTr18XQ5qiduj4J5AdfwMLnFWsGxMr6VLRT7S
zPWaU1ORRQ0iJW7LszhHARXejnNZFwRz/VjBKu/mYAVLhHdwy+JLfwAFOIXwcSr7K5QmgUfLmxNN
iZesAx+sJP5tdI2BFO5uan6hHLZMyYYisf79y9EDCsdh/j/NcOYhpKO1r8tVxNXENY/0ERqO1764
PB6Hk2mU/76cJNjvGmtu8W2wGm8mBg1eBsqeuUoZP8BaU+tuypySSB+xhA3/V7a8p6QnDUKfmovi
WBdlMCNdN5TAqq4GC1M2jU+dlNBK3Wi4jG/LXgxOkdCA1uNPEMNd0Aw0MN3Aamy8TCGyuf11pY16
an2TfsceZS1lrBcT1UUzErdhb+vzl16XF6aYuNbfinwr3HUHAqSUTtZkRznY5pfRqOlMYv12Hv1U
KazzpOEWLG7Hs9B7ykBzuxbzIqHKVe3hCgwgUBoYpGRPyIVOqsLIFhCOyjAEmNx1dCSxqDET9M1J
J6qORQViMPXPzlh9Jm1kXls2HrtCfGzICFsoDmiQDeP3RzbZZ6L9fMWPST56aomikEo7mM7bY0OT
0LmcQi/VANjp03G1LS7OsPShfKQLdyxg8mQPtXIJP4A9OrrWv+4V+8/ciog0MAXCIlXX+jsWxzOs
q9WNjYgyidkb6/INQG/ABMKHmHdVyn6SuusuuB0H525UMKPTswFgxmfZesNihh4IJMQIeM1mMWCq
q9vPUBe00Y0dasf0X/CRlp50eVyY7zCznlua5lBMVr/hIG4UMbm+WsKhjASWRnXkRJqeCJtZuQuK
u07YXkIk21i4JN5LB8VNTbSlC/fGAs3UrKzQXO2Pcav9lbclI1jhWlJl1NYzkUd8XZkuzM5XbLLb
P5GmXCOAD6CzRh8PHLRE7RwE06NBA7wsl3C0Vw5pVX6WIOdb5wreQ9SQU1Wq7oaJnMEsPYzuPtH+
pzyS8+9durQJH4zDnyGrNY5V17wfL8hgTY9FL8ntNVaAlj+D396ditL8EBAXWRU9fLrL/ncfM8yb
rpvoplqYbIMPTRYB0PMZboNTDEnqSXr22A5alv52D/IKduz7qWZvrJ1v8puUA2vWj4I76CqRChAt
Fqfl4z8j+A4U4H1SAMeLGrUgXSDBQQhHzcFEOZv5F4NQGhewgoLpeCqBCvyZ2Mv8pz9g9k2LDIeY
mcGRFfz2l7i5FHgM5w+zitrCQzbERSCcyr0+hRv4btQ3WaZE6GvYrdnwKenseQXTolu6d7wzZZ2i
hqw6j6DynvWJ7yzW8UF0A1rQhf5w5QfWoLix41gQltrl7WOUgnQCBVq4au3SOEmTyUucDgKUy2n/
rNLDTCq6WyGa8qLtaDRHe88QZpgT1yHdjeeTZawmpGNlZwZD8RshNBrldu/cqU/pPfVwdqzY/zLg
/1PSwQbd+XbG2jRxkwK3UchxUxjQGWFtq2UmbgyiRp0+KjIqogqGlPOEhyyIv92TRpjhvptTE8Ct
mvNDWfc9Ukw41bgFP/oEEQGJLWBL0bEi6ouFh+rJml+HtQWm7nKmmzZHq231xpsObS6MYkYoRNsY
fVwgmQ3n2pw5qCsoeAHMLaBnVm6hfqLFI3LP7MT88gcRVJrAHdbtYfcm8Q++uooxGbRmWEkIxJDM
emPfVmBtTIQnofi7O9+77wU+Q19Ty69Yx9LTD1OEDtShCT9gc53+7XXHS0fMI7obLiBBccjWzLmC
5lP4WbT7zhkMYdHWrT4URAxcP75l8OZZdrn3an2nteHRcCspH5RA7CUTMMR0/JhSZA/Jpl53mGbA
FrJPELMxbXbvDogKEEgdv1DC62CJbJEakhuFBs+eppj8oE8qnJTM1jwIrLvKE1Erko7Q/bTa9u2e
GTmCSbzRBT8dkE6Q+1MQyYPaeRk6IdGEIEr/8HTRaAmy1N+HrbDE/FbSOwUvKXQIc73ONOdwO9jK
/FmyWVBVP6O3S6H/z3m7KW488hWd/hfzPpuiuHm6B05VUppvFI5Gw70oWGrWzre4SibhvrkcKMaE
JKukG8LlRwcSso6wTGPvDevqcmCwjt3uEhSvlWK0s74eqi2khkOXHJApKz8EIKIlp/ivhWutAQs1
Whu0CUFF89Ho3YoNla5V8GAnPJiRqN20EyEIvr6py/QCqIRQ3W6GuxlrPy66kV2rMCInwLtAxsvC
n1yhtr/m7r99KaIcFEIbhWOv++fs30xl4ZOuuZBIkDJI6ROqg+HFKG4AxMcrWvLzNvVZnzlN/YyZ
Nu9KZ5GhFtzvm8Fh7VkWZULwspspB8nstC6l5pZ7TcyAf6soE1P4IdLclk+RBLr6Dvopt7EKvEcp
cmM23GhEqrPyvmETFprT6aQO3AufJILR31syQ2tYn4XLgFonYFldgDPHfIJvTsd8/aJwPL7X45R1
EGsWKbpHJ0UcJUo1Z7x9cmzjgNITf+24gC12SNg0C6VRxnoVaMdBGb8qX9WhjoESyBrBH5FAZqTg
4YTnF/404XdI0Ro5c+Df2PBHGhfAueBE5PVhfIW97UozXdS11ShVaaWwI2XnuenpXcqlTnRx5mXw
A64MOA7ZBy+qdpFH7jpumd2bxaY7CgBCIUnroih1nbhRVb9QFJHSQhANmZ2nQjCsK4GvHdWk4gV4
UEdoF8P8Oz6QGiriobmHfDNkS5qo6KvvUQ5/DuFAsgZUv2du6e1B6iSohCiFmHCMnUEDCOubbfvl
C4tKFhFW507tGBZekPVTLtI8d83JMQi+OMggg34IexEE10z30r0Aw+RMVq5ywQbhIeb9bStxGE0n
z4MlBpwkyWMJSWoEhoOy2H5sYUnBBbxIHUjAxwgjlK5nlR+QxoOWSXOEKvHNhe6SPEGtoVKlMWf0
DY8E8GntHHA6ZY/g9Y4tOrCHezS3BJlhc+Avo3kXM+OiX4oQySBn/xdNJOVN6aAUqypcy+sWS34s
h7c2xCYLfUuRw+Vk94pj5BC/UN7cfWd8XPbMEV6WL2rZfhRnKQaNr4KzEhw8thJV2L4DQBG+p1yG
KpfxfIdGhIC7H2u8BkkcJRK64Puqxb2lIt439kDVNMJsBX8LmgqnlnYNkr38/Z5jIi1d1Fs4UWJ+
0vzASYdrIf4gxuW9RqHznAYlRKOP+OTVhrfsZ6LHTaUXrGd8HRifYzmC+26NgbgNqdaYXVEU2RGF
PvYxj7WmsgCaQRyTK5ISDnRE8oEGcYu9rt+xisSRdKRsG4kHj7gomj32FmU2e9zS52NeF8+sgqkV
YTGQK+cHnQRIJl5BIpcv+zONvAx4u0+Q+WsDIHtlo7mEhcBDssVc0Z2tT2lx3N35bfTkq8ZA9GKX
2/evjxIlMqNmFJLMMT4WdhUXGGboFuJn88CeautoEV5hnjhcUb0z3rPGUkvB/LR+dL4fcu1SkwIG
0KFSNVdL07QawhXs8Erm0HUNbHgZ+ym70at/jhGnmCS4MJBlNHvuKPsBUUrKEPVXmmuHPmi4h8J7
3RRDLh2BtXTepcZmWb8CgHmlMPD3R1NjJT7fv8fUGklv/pQHArKrkhW7hYgkycHAtFAUQDGSi9Gt
ZsQZh+gEbPr2ZTe47m8Jko0H5fBQja5arEg/WFb/nNjl7JLfkh/+RQ90ngKlC9f9ZaO39aJVb6he
g5PAOwzVuk4TYtDi5lcM8Pn7/5LMqZaeUCBZSIg4jiZ5UH0k4LTdl842TJ82iaBYQ0Y/2GrmHPbv
Nanx+LS1ntVSQnmw7N/lSAd3yWOfu0oyiVe7yuAkySsdYpSreifJC0M99Ns7ijhz5nqMzgFz5kmW
Fng57PEAMNS/GpTqEERk2+Z+CrNzGx8YGYa/3rp1s9jKhF1ima3bcUsTFvCxK1suWfrzQjkT/GKU
vC0yoEsMYziFsLhImkCyLxuNLxRfAmRMuZcPFG0TwnGAQLOmjezl5zfbHx91wPUo9K5yY3gMwJ4F
FMoZ3IV+dN1BkFIqhI+paVJEWTu9id0R7XbOQBNAF6KICira1s22QENGBtObK7ibguiCgl0sfBf+
0bCmZXT6dZHgcYiF4OeF4rtvHm4gspWLdbTb73ZcfMQP/ln16XsusCzTeK68g3635yrnAawaB78l
QtE4LGWHwpTUIB+jhrBno9o2tzZYzoQe29wcN5MrDPh1MAwUY6nmjBSU0+16BeMNcn+VWHYF28TN
G4sSwJ5FY38rqOo9K9jCX47EARI4+F6TA4AvcR6AvFOvzDXG5xx/M1NJ4E9ZHlTa1v6CSVxOZW0f
/xphRzXhoJFiZafTHnt6mEg95B9XKDnX9Gtdo1l4nAoiWalmCT7+rod9Q/f+cQa/h4OzYmrvsv6m
NI5QWT6yiKMElhXtqh3RZecnFYGIbS2jYW5bEeB76dZPo7KYpNbBjdRh+TQJtYAK7cSlNkW95EN7
930xDwnd0fGf/8xTEHAe2URkuaFskMSDgyQC4zsOBCPi0iv2/Qwhd9Qw/X0OGD0j40aWNqOL7Aal
t6DqNI2KJdT9SjAaLw68iXyI/sBsqJo7nmpnsuDe0IRya/NE0s8p2T6gq65DkYPC5tHmoy6kE51A
gC38eLVs5NMs145cqPAxXmFa1BSrB29pqVq27RRJOQbmjm1472K0Azz6jGhvhaWAFWj1XmWqJeCa
p4sMro8gzI4y7MuePBVDSqijsPaDZG3cuJAxoljS3z4UEbrCg3AjPXXECvMj9XIBSka4IEphBjnE
jFglqE+tOGpYFa0IJ/XTpTyNGMm2TFwmBl+8FK2clxRSx+Sib3ZgYVE2vsxkxXNYY1pQmqSzfvxz
G9VObPsEdobiyX4/ZPixRj5CrvqSEBsD8B8+NRULzjpS0zxVE+1LYRruTtOMD6vOX6i9gHWm9SaJ
UOnGMVrBCk6OqfQEj2Z5DJevW5qQCsGyi/E9ogcFB9r6YjvysGpAHQLYVDdaABcDCQC47oWSXAtz
p0Cn5lzZlnkIntokav2qtBztPTQJSpOv0IhlZ/OfHkR7eHSvM097Xh80u1u+a0jSdmFPyX58dWsV
of0FKnWVa9Lemu9xcroVtMoAcSNRY9s1zunTgvsDAnpZH3M1Pi5JKX0D7O+wJ6LUn5Ka365kroEr
wN69fNN+ca31VClkaDmPlGvu9YSsTBZzDToY8iXZ/ZNxGBgs2UV7swrkDQKLmGA52WJELMcIryRR
zDKB7GrdQuHeP3U5uPXPT2lGzmwXapN2maA2pkkSRXW1vEozPPQ21TS7FouU3fhMMrUl19HIUjdI
G0SekEGe4NTi0JWSNFxLHwZZwf9+tbdUI+IIZRJE2PfBzvEGlq+aAGbsdPrb+8c5IakVMHYiua/1
wAkcqEJPtca1qgWHYo7/fKFyqSjvtGJ+DFEuXGZYPwzUYSoQrlTFP9G4hH73JYwlBrnBoje61Y7e
dNy2WyqfQyzxj69UmdAbk2ev3YxyQP6Ca3xBNfaXwchmasFRlBJEtseKKhXtTS0geIetL4DGZI1S
5Ut36Jt4hb8YyHyKvI2emICZAX2OYlaJGef5SLTIGPWJYoUyHNtGftySG/5B6WmVcDhDVC1k40bA
KHh3HOOlc/sSuMxPXgc+zCaTKKhkYGKMisb5Uv5PgJUCc4ChoaBekdQPdfBtBP13yh0BwG9hKOgH
0tqPQZ8dTSeGyr413fWhc+E5ke/9MS3XLku+2LNqd/MtxLC2ZCLmHWoQzflr7NNL4rjQiyMZZfha
9x2WFRieSJ/Tgk4oKlI8eEg9wA/CuxTN50SQEuEEOb4b5NiNHpxGQ1wB7AMk7VBiTrUv2l/OvOoN
3tZBpmH+Q6tqgS3286PceTJovMRNYmJ1aHfuGi9TeuM1MxgQa+nEscZfNtF3ogRw1X22gYxrM5Ly
j/oCTGN/jBuS5+7DV9YjerMXfTpMGVLzZGlzPaFYquH/8ZKlN/zcae0cNQnRCND3tKzrf2zLi7O/
pnvuKUrOq1QopNLXvsyVp3tZ0VvukIiQmgXbMx4WIiO0u2ygPo8dx+Vlqj8s38hKsi4a8rapSrWO
1qrIIVH7ZlFMd4iqLmBesQmsum2G3y2IJTX3XaiwZuSokYYB0NMxDx49NRXaVrA1VlLy7QCQSdRM
V0hUBEBQkI6iimqDlJ+iTCfSDd0t1Xvtecf9GIHdy8mT8/b6EjdRV4QWdGSSiASvMNXWfhUWal8W
tCfmdrLtnxsqRWyj8NOFxqV8X4ZGlzR8ILWPk077Em4eK+Ff2ORdTOo82m6btLVIswZZRtrZ6Z1W
1sFtQ6B5qySF04aNgbO1Pk7P1FHOBuIJ2/styh7rfInXEIPQ6sGRttFpJdKuNSiEkHhMc6iZzoQx
VAEpkRShpo/yl+fydJxhRTJwdzN4G5hFfQgFdXyMfSXqBA7j6gkGkvtxBEsmA+EPRoStl8CZEDc9
/Vy5GT2eTsH84WwbzStiYacoM26F9aild4hqW76CWdcpFOaO4yB4QB2CJKtaCUaa0mezIq0fWLKG
BuYfFuDxe1Mlj1S45U1M6AZTlz/oaHs+uKlk+5fEP0Ovb1MAFTWd5kBiYYu7iN73ikH2EU7aN+er
xt2Cz9qktDvSCEdMfLBskuRJKX/9/GBeA0r0PMdX34tSH+NklNgDN6XDskx53Gbnw/Z5CooIZCtY
kKjSz+YgOI8c5gHovHMnJQ2AXb6MXAaGvId9xmLrxbsbF5jy7URgcfJYM6dJClFEiLsY+AOpbmMX
fJREbwW3bAuC/AgZ5sIWxZ0EQaOqRdmQxUXzaLjvbLsTYS0SjJfy+dxnGwZ+Xxboh1aaozjKw/6Z
dzMx0LY5ds1CPIGuAcMvSZlOZrbCPlmXw47fZru0cNPhpbTLBgIktIwWbFgYs2hWdTHpqJDpLka/
+ACiKtj9WIcvIHOYQGH7dpj4Uh2p5vMMgTnx2fQxNxbmt7Vn/BQuvAPfldTNjsZLEzvX2r3RhiMV
k0xsgTeZGpcX3akWm15//h7WdjRmrg51FzgUMYCFmm7Jcs8zTmWG+6eZl3sBEgEaOZJFHK+lvkpN
WzItyksGBlr6royDXgBY437E3HseNHf5+8LKUfKmRQN4WbGBxqKuJji9JCIAzlxv3zM95OHtOp6m
sjLBA27idyfX7qAG0DJIb8xSgmG+zxqfX17fjhtrM5Nlu58NiPKV1Idffj3/hgOdvL39mnUP6hLs
f82VBywwoISi+zRlF/B3NrZajsNiRDglKb1K0iQ8pTDvsWQy06H4xxMyPLQktvsJ/tbrkZt5wQJA
tioK+Ynrct5qEgHDXWkrMTVyFN3khM1TiUI5zRnXwmyse2GsXisVbVdrdyS/tdb9oR49+3Q8wzzt
g23DXxPgMxmiathdhlqu7qEqgH+YMqAnPq4wV4n7pELeNUYgZaEyXZc/Mt2u9YZWYIGYw5np3VH9
5wY5Q1bUVi2ZEH8qlddDfPoF2mPuGCUJIQ0TzZWFi2A4cmJJ1lDiOboMr1zx+zBlK4w+jilWyH3b
LQZbUfbJBFqSJocaOx3i1wSHvJkd4EeixgnrAjef3gRfD5HzpoyWh8nXk7pfowYyLcaltmnLNUZ/
2fvjiovWucp+Q5pTW3rM3kB4PkcztAU7i8vDxF3wTXqciAbkjyWxiIe1egGjFj2HmkrKjn22T4gU
AO2iINEDRBqoE+zgTRECYBDfEaY5H0j0aBuMUkumOrYt5yiVxa664LCJCiqV1gZ9POJ0KcumqyT4
3ZwrbQ/8Wqmcx5q7rr7hk3W8I1IaVFaLnvMFTWsUPuuwky4GbhnDfdAgU8ZVeM2fc1XEvg+OpPW8
JvkSGyswNpk1Z/WJb2CrYL69gQmclBkrAZGY/COcOsrGszx5fMQCl0YX0efiIaeP7+6t9vJeqC/v
rgvDHffU/etuIHyINpNkcNrn5dU4Ez1CqlMBfTbSdlzBNnvuqS6l54zIR93ymdSylamQzXuA3U6q
EXLziNfFqGafOynBdfN1sTLeNGIM7OwpICZuV9hh+S5T8Lrfe/K+iWCHz2hYh0XSTajfZP9pRN/1
PQDviwX/vljEkIPNdkfRA6zldgItL2Kiy9iQ2PF2JV72q2oBPy+WxbIidSYSzO+Z3pUbLWPhNK3i
IHMuAiSLpoJkUKX/9rBa55ybTpIIg9AaDQfcARwVRPdIuQpICDwunWhuZbc4spSCU+9LbqYD/oaj
8gUBQG689DgnhHo25QHp6fqTyo0XClIr3jgUvxdMRJ+oLYm06JZkGxvGu6GonOpEQbFDlNpyZAYq
G7fay5LMZrNyS+5Na+iMJf/JchdEZkIxTcBLM3jsTve4lbxbAMlKY5zg51a12MuZSiNLyU4K5c18
VUSVe1RwxrAGaDNZ+vDaFyH5qLUrFxwT+7jrO5I2bzwHswLMcDqtYfmOd6Nz4EnTmPnhqlTXpQjH
KPUUhWAmuO6tn9JW4SSAu3dx7f0PUoP/v7L0+7ZbttJwPDH0BlQD+LBgJ61uTb371gOH09YoDIAk
AEGGngcqpIvVwjCrnz6S7a2wewWwWtSq/VyFTzD3dsPoC0VigU/dVGWiKY5SSmESy/MD3D4o8rH+
Zg15dleuz+AK2matLad4Nx55HYcOlMipqKecCO5yuhWIdrR61aRybbLw3o6Wr2P6ltpNCkDgoTAO
KgtiU4WjnCVGMqGIFuOXoOn9p/L5IAuZlbSQd5Wddo6qUaeUrzLa/8VDJxvBSHysnMlDkSzvxbwc
vQP61oinTFSV6d4jns+jDGYqx7rgMVaFfQNmFne7pxBe1QR9cm3znpkm4a0v2HQmh/XWq5xxK5Jd
kFNvafyvAMmsvprjDQ3+0qXyJ5X+B30snrYquurFdNiQyFoGvvU9aSZoP2WDmnO3E4guc6jy3pyK
qq0GfbswN7DRvOiaJXEMuLjYyBaNTWCKWwP5Q9BQumlkMFJbbLwjZLQewKf4EOFNcBMHKqnyZpHI
hXJHUw23yT/RxmbrdPJOG5ypAVDH04SmJxCDkWjPWWq31N7qVU6HHagKrWQ68xfRKIz/1qrCXJ65
0cVyEIGXG8m3eo/nLPFOSd/iCnljqVm7Q0szdL3ojSlt3OjA+nWOzl+B2MtioD/q/BNzlWkj1iyt
U7p1HRVcaNfOA5Dx5fNqd+sb6dnB/f5FFI43cE9h6UtGgu9/9M0/pgu1Sqb++cNArqztMpYNAGdu
FUY4+gyfNMNGsB5dqRCAbmHufxLLQLHwtS3RFU4HewjhyOIcQzKKL44u9jRt4VcKE9KYQ6E2I7ZG
glu21g/ZRmIDGNdKD+o/MYz/DjgZ7gy370NwDQmVG+3Ew6gNg5jqkXmW7UQfv1gY9JAOryerwjZY
9co5PRh8FQckilVJpwtq/2QNEs5QbGhu/hZv+BJ+kUnyrlKivthq+J+TNeILuYfhmTyDQCTM47jt
NHSyavuqsaaO4A8K8pbJp0cdK5U4EsiiviTLolKMdgAOBt73FfMUookiVrIsQliYV6nhm95eV9iB
YUNogN5L5LqkqoDz+/hh46OsF3o9SrP4QqrA2QWLyCJPDZ/SmhKI1prEIA4s9w58Q0vfCcPqsULq
J4CoBA/x17CaBFKmVjTnjj8ZtWFrEAEFgjVSdbaSCETxEMPBkxC3LmgrO4kK7dnS/+0k3JzKC8Yw
s/kPdFX4OiLV74pl/91UbTTTSYE6T5UpQhD4MbmwO0fJyzm2p8PkMpqyDYix5OrkNCHEmVomcY2i
wjwcHvqlnHM+xYKhYYilVrQkr8z8An6iC2UWBkAvgy2k7D7DaVb1bt12VWnEGgaGBYoOA8FUbxEL
Dtzpo430Wa8yiPNEUbepk7i77xKIkKI4QfQThbyTwpqDA1tmPdtA5iKj0pfWSC/+PJELcjX0U1ae
3Kyhv73mLiomzN013ICORQX63LDu7P1Jypi8ToLoiQuOGtsAs3MKXvpkSTd3cQiSEf9j2H1ZrY5r
phuZkniSTUKcbPbqiVHy64kvNmBUFhEVDFaR/35eytidPKU5NBcAjRoBUgKKVSLoGNrniyzwsCl/
v/yKfkGUNOEADX63FcZuHki7mEz7uubmuH8WNIayVJEKK70p6JZHU+4JO1U9WnbFpe1KqTgB1/gZ
ANrYHfmi1geP1lv20ndh0IFJz3JnUzqNk4iHIyLsHcFmqdfmKwPYD2g6gfSQMTpCl33WQly811U9
D69SS2egcgi2LFmZ4E6zyytbCOuLdFOzNpXa2rZFRru1ZOi6K0zjX3GvcNUIds+xplX9HV4ZhfTM
spoExMEWvd6eWZ2286TNa/O4ii0EduH8B3VI+XvmzZDaH+JlvtbHeyESskgFpM9RO/83KLVa4P+0
2yfxC81uz2+X/M+GUQpOD0I7KElGzmglKgBjC1sHet1mOGIya6RlTm4hbYa3vGC6rkcmNQDxMZsg
WGvKTtGK6kqemFEJy8MYBbtKwIrk+e08RXpZgFxE7i6+I4TEJigvv6CH8rLQohuU+MkTVKCv7+bx
51M0QBBRsxOPPn+zX3b/XDqgQPE6n8c3+yyInUZCSjiEEftSuNwXfsUanJDSrWDBxCuOTz+INWO5
4tBeLeOXl+LvWcQP1ngurtq/ISGVEOYLME+Fue69OKlgtVFeeyN6tOi3XN0q6JVwnYlgyN9pd5MO
bGiY0Q+OYvYjGnJ5MlBAbyXF2UoNFuHFhQpg5lyqKMdVvQwG8UNTRvifxePxj+u1k1HdFZQudkT3
FbPrb+0eC/kQvY+yc1lvL9KxQKb0Z8wVt70ebJSVqC2kVpVEyv4Q0RdqEZB30DYsRre8B+Iwaj75
DeB7mVMD4CL9OLVNeT7XHDTkwH0EkHeCsgFmJtXP9sOTR91m9IMiQOdCjLzaBUz6LjJ7uf4twBSA
BSaXuooS7GgxW2eIxcEj6yztWwkONOIGpZ51f8aZh+6dXCu/VdO1/mN7/EVYRVRhyxjH5WmczeWZ
dKjqmZaE84S/8XYkrj4PtHG9ONt5dbhoXQeeACPA6aSX/2l72vDzdWjjTz9iYuMVeSbaNxEiPnIf
GIAdbBDuhPTTOCsaI0yFGCEi9AM8SrDkjBfD9MrlGM2v0gQmQ7mQ1OjsJNvWa5Bey+NpQlSe5uVH
GWzc31ybNBtMiuN2v2iLGEQST6TJxYgtFCsGyEi7PNSNYvXk7TOUnspFt2noz2B9EJsX736yRukS
RRqpBetbkoOyZtSx4XQuY0eEAJRaAwj7vuCNKoSxKzLlSP4zmCci6cVdZJiPDQQq9HdBrJBsvKAf
gR0ULPtuVk7WCROOspjSWUJ8pDLKqKQHGpqakeaJgn/4+hT5lx0wLn8dZ2A2tlJlxJNz0CLq7kD6
ljc+2M6WBMCB+Mz+y2i9IoVpE2cW8lNsQ1QPM1zwWB3ogga1ExmU2DAB9Nl9yV4nGgS2SPmacWKX
efkZns+3GNSavt5fTopLME9kts4WEymd8JriT/+j/Be497QU/lVZHUIzwLKeWbOB+ILBLMaKAmA4
CYwPfTqdKogipYdiH+HRtTKeAu3hgN3muKWzfoVtFLIMomHJiyYGYnbAuTRseogDY0YbxTUAofIU
OnHlW3U8EpgmuGMCobMCxqqMsuLhRXASGlwoIz9ZJGhgecQ6BxD4KNU9HcJ7779/5x72zgpdGxMO
P1vjAQtFNyrpq35z7ACPr90Hb94s81nRSG92GHdQWni17RnA8X3MnmWrLl6akDUMTB1ANVufjcg8
kgQL02G0+oGlJK9aifP1zP4dGGLd9k/12G3vxVsbEA1MQr90hagPeS6SCT50njN2ZmL9rNcXQKmF
2x0jCiIx0AcL9V6vcsTQVkjz1U5vC4lEAjc2jWqA1uRNm9TuqKtZcIq5NCpgKhZcibJrbs+zbjB3
aUfDbLkOlxjwyy0ppBbyZtPdgys14sR6q/ffpgULBFNc8erOucgfv/jrPT7rdNzrclmTQvcTnlMH
430xLBiC/9l/87sZYiHjadYMriTym0U/SBzgEP+R3LiQNdP8ZorEa0s8B1nWmyRAFUuTD5p3Crzu
TO/1k0WEJsOPkeZL2i5PIrI/oxYT5Qw/CA35bHSPtlKZpeECBNEi95ILpPhPLJYe1MT92XfDQi/w
00iGfP7ustq8PC2wtqrRet/p3oyIxGgy4foEMdBk+B0ctbnMhDVpDl8h0ZguOUWMhPSg1YgmB8lD
hw2ETuZm6p+LNR0cW260mp4hngaUEAg0ltWO1IrYTV42EEmRjJ/4lYOh50HKFqbJSTCgBu2RHBzI
qYmUB0IHtjspj3Pr6GMKcoRBuYvZcYiFmmT3wZu70HlTeKGxmiKDe9g8zcaq1Fn2+fywjrsihdvk
I2/RQOYq5tRzb0rLG4hbpDPd1K0FhgJvRIAAWEQWSwnpy4u79KiGVyDS9hMLXCEkRIYgmG9p1n00
tac1ebdR5VTIxPdiBIe70cz5hLw4TSuvHncl5FJSwlfCx0JRFVDwMhSEkuQUeM0qylaq3QrE+KP4
fWMPceCqlO/Zsn9aSiqyZlA5Z6jAQB5FE4aUq+u77H/zCDk0bRdl5cIaQCZ03j0M/tePHCQQFpxV
v+9jpYBIJOxALkNEcheHkomkXYKcQw6npvKBazPa9c1URTol7jceoS3AC5wucySdGticeKdgpzNq
zsgcS676CeWSly5lMpOpPC783JX5o9p8y20T3+L0BwxoJTlybeWjykS4nSDCpnTisRK++uMRCiD8
aC8LlUT41CaAxgWU2RcpKfEiOwwAdXUxCfPzjlThLejGq6ajP8UJOqMdmBWCrWVSiYzcWBL2El3M
EOeb8uMiOW9GShAnwQDzygfv7Rl5oVzVD2WlMvJCE5JbCvKwe0bRIUIi4mOnZsMcd5omiezIG3gs
tqetZJ29OeiiSZggiHjIAlt3xPimEoYs5DCDokjrOTwQEn2IdEkYFHoFYA/92fxCrXEBIyhz9V74
TkttfHmQdKYA4p6uAIFMFKkDfKTFC+Rr5D3z5DEQRsGfr9wKOD1YN7jbpEIberLm1HLjjUwDqarS
HxojLKIb0Nuos4NSajAdLYrtMtBpTvU4A/qTvD7DQ57f6zkltcOQzonSMe9vhDfleWFL9j0gPZ4G
PGTvLLS5dH58YPZ5VbhOMcLMwckY/lT9CKAoiIiP77yxckeMDQ/by5KzTzIjyC+30FSWLZQmvIJG
tdbEig/J3uUTMbRSI15AP5m/1elB2to0H0pDUCLXAM26QHBG/vV889bmFGIIKd5K8uFa7uhz8/co
tQ9KOFw1ySZRlTVE2ta8pNpGo+k+mOHzNMhqBDjenILGfG5WnKQ1x/qxFe17M+801FpE8201LaH+
uqcODk/tkyXon8Ib41h78mB+mGiWtwnFFAekUQMI5qRuL+hJHSPn56rmdupFJIrJHAobyLWyLJ/D
OyGUlisQlfHpjDOOocYhGWpFxZOCvrTRDtEAbrLIVNTQv8GALes630LactNy5/p32UVXdgKe7ZQo
XaPDjoDeTs0TnOnQYRHmFM9EGK94qtp6JO7AwMerhkF8MaQ0Jpi1lLB+JS+kaUL9+Ojp3qYCOvWK
RAnfxK4sd3TqYPK+dSohSfZPfIQKj0pzKvFJ8TluStxqSA6T29MSceYa5Io0AqCRkJmqhXYLoVo4
ANwjTyIYzyWuG4FeZf7B90QItbHipnkpNpryqCTnczxqtB5CM4gtxR+u2QTXtustZ6Gvbs7qIDi0
CqwANGPU+HTmM6pLWhHUuPBei8jKi7q/OF4OXDyu3SOX3E90R6cddvzk4mz+GmPFKow4avmxFRYd
DMp/TPS3yzEa/pf+sgLAlMH+iEFlD/cLEbkaydY25QrXFLSpGfdk9wp+y4g/GCBR8IPIRBBAif5P
13w3niMr+0G6pQPU/i/AkWz6F5ZsToa5hE56ISOwCfMvjX87JblOZTZv/1AJnFYx5f6u/Ui2gURn
GPjw1k0e2ip/Bs7SBZo7cvZzMbvRoKxi9l7B+3jbetWlgzKFPjoUKVhIHQWq33E+qQGCcThj0QOM
Dm3Up1vRbHiBprGFLRuDw3/i5LPB1dVRK/tBFnIms5Dn+NEd0VUUm4cvMY51nL2yqRMze159q3E7
iu0W22DOgtausxj9RmEJ1pPrhicaV87gZs9tkoVqisb78U/eqEtfetpqjAM0eBWXFfad65zli5Z9
oIS6hbWGuk/7ynP0RhU7z5WVScwIASGguWDA601FcSywHNg+uRk1m25JiGtyHvk0t77xd8eLMq2Z
vd2GPk93bvkm7EuAnaKaOp5kYvnHEqjibL1C0sfGSAEj9cTnQndsZj01haXFaU3FCUAWa2VqJCh8
HtgYvbqMZCigYNu3YjuBYrYj5iWq1IPX7ZyPRt+1hQM1Iuz0NXBhRRek5PdgxyXn42e/6Pq05cUY
bcWw6JZyEtWvtvigRhNqnR16XYfB393GzNM/+VLTBnMHtyoaizGPL9bXGS/5nAH2NWEP9nTxAZiI
NNAIYfs//8zEmr7MPIXO1rbKJJdFLFPGr7RBfyzE1KavRVFFfpDfAM4Zbsci4Mo2LthJpImkTWvD
2ghDYFwv84edm23tC/snS0OC7jBqC4Nf089BzshRCWKuq1+cGaMupok6sPoKA1Bp3h1FkMziLbO/
XY9ffhJJYmb+I4hjxTVOLSTgvq3zjQ04zoGIv7ei8n17IvDqpYflfGg1TqQzq2Yvx36VBEsBqzKa
ESwq4qj1I5VjDi/RJiPmSLUYM904L+nkbK2qN2a4O46LrHXNgj25WhoLOLxq7DonDPDy73XxMG6W
95l18m/INBU9E7MHkuZ9QPQvSqKVbnCSMPEyWj7jnnxb72TfEuGTVrcWEvWSlqI0+s07spFCuGrG
4ncmiokD1SFPzPvVv4eKlrKOL1LJQAppaJvD55kFPvR5jZ7x1vPYWLEcnq8vP41I9lekwDjgbwfW
uO69fDvNWpEKi5oU4mh5nABm3B9OmgZUW7wSLnI1D1TytrNWHhgfE8X9gvMvqetXY6W9+DMpelw+
9lWYQ/Kmfl7cS3o26yCQ0biWim/0tGuS9fNVs6OqOr8rO/yqwuARDR30dKNjVFz3/1VqnVy2PPw4
ji5rWYeINdIC2C+9uFV0rcIoV4BM/suui0UoDlPVtP0G5OpU3NB3AEsLAjSey15X8alb982h0ySA
ZbkVNnO4tDa+PiztAWnu4ZbnCSYyy+oowOA3+FwIPz/15DM8PHQ7cqAte2DnI3izrKhpToGSeD79
ASE7M7Zz3kJ06doI7ayqi0WPuKzEbvzqMaIeH/YFABWEt2luAjfEJkLhg7ny0ume9FQrRINr7Z6J
RitW9a8rOF3bNa0gAdnQj137sTCsh6+4Xya67atJVTCUo9IBroGbo5xUy+XXOggEwMqgmxtzjkNd
bQk0u6XtFZtglnRBM3IZzBGOEh+thfOv34Dq/lRdqNYesmajityvxMI9BmuMYkb15oOp1uRTBboI
3URZNSET2i7Wqi78bQyFQxyIeu9u1D07k0QF6NZ7Py1aTAhSC4FkUjzOdmpEZev979a3BNimS9o0
vuhKhB0v3qspbBU4ObwF/ABLlh0b1OKNR3AHfePeA7w6gW6prUWlxi/V5c3LiCxPGa80OZBg6Kld
YLYi6Obl1BX8xGxvhptbhwTsNELeEj0T/FCQuWRKsK3S9lxzvL9NqwuFeI3fvhih5Z4KgnaDLuD/
K8XfErKDok79T6G7GLtQvHTVAo67q1kX+YTsZVoen4S1iixqz74eu3Ou6D7djwYbYUdvXwXQJIHB
esprzPasVR1AcYX/QltQN2rIJPK9Uq2UOFrP8OfQ+NFxCzjh/g819ARx6DkPqAs0Jp21rZk7aUc+
u2B4dALaqh/AKbYYvTjNNykHPdoS4DoTtONvt9V+AHNrZA90xVUu76+nYCDo/AmaSeCUYRhAwI5v
VT7A0YChAnpgaItACHz6lbi19dr4wWwk4U177ErOW5Wo9usW8VymfTztRIL7TTCvi3YfYeJtXo9T
EEEKZFE9w9pVShJA63bpbU1UzL3VZYChBH6E4lLWtkJ7l5fAGoi8/ZQntxVyHgfbuPSfH8BbU+is
kHsU0ftbJWzgFb8wmWdLPxnWk9jxlTsptzpgR/Grf5cQqksDej+X+DyR2m+jfhysjAfJkYDUcFeY
Jb5mCxK/rVexc7xDBviIIeY+PZfF9GyCCsUEcOpy5tmQJJlt1OHYA4yfkYSx1/4c5yzSEcNWDvvo
e8o+KMhJuFLh9vG2970ZaZR8/ISwzZLen2NejnZYk90qsa2xgg/6vadCnvyikkoJa4RsNR6BNNLf
/heCkCYrKtihVVhxDHl3P56lnCHM1vB2pL1M4sf+bJrCwZQAlaye7DHzEcpXO4rXHdSHeHlo6hUs
QeDfIanfYXw8HLtrSaenhgX2ea+k6rLe75H43kNri7KnQ0aucr9Dsm+TFYu5wWDXb1I+ox+YezbV
tZz7aeOYd6z2IgjoDCb7wlnCJ1mVBsGWpmL3VKaQA5OhlyKMBY3X/sarzoR+yyHsLb19gqKTLYXg
IO0nkf3QPD/8BR6eVX4DnuDDsVUcGBD9VxWez8WDojBvNNJnc+uRuu1KvpUdVriD4Ny8wXZc85Yi
VMwjJiZ8Gkg8fVv5BHgpdtzmiLOfK2BuJ2ws+XvrGJlIZGM1xsssO29V1n3HNH7k73l+MJr9wdsE
83UnW31uY12xCdkyOtpLeoiONUi2iFGKCjUeEPJuwudjOjYu5OgzizVNjxtZq4G/ezefe8TKXlFw
d6ZiUTWXTJ2gaZUjALRVsUENmsJf/f2K4rvjrJ6ea+z1rVab+auuqzNADU0m4yKW+pDU3s1hoQzg
fkmcnk3G61HPT13P41XWLns1PFRU/C5fD7TweO4Da4iEdpFPhkOLG7RGt5i7N4PrlBU//2Sq22AD
Be/BFmCXtNiIFCC+bOlmgrLbNAW8v4a99Kvq+ro9stVFFbapYFgPBtCIGb6l/mSVr0KWsJU74mjr
8kDhsI34HtkpjarwVVOry+xUraYyQIPtEY7gkQjpBLpgzslQ9FFfPnZrQ48VZ5xW09CQLcdKhwFA
4U1jeEUUKsbHVObF5zqX+7mIiAurwZq+h5dhZHoKV2bX+IkbSTsmSgpOgYY+sZUIu4dIwmFfgI/S
B4smxDIjUfwuAqCv7Yre5KSGRbJ/dUYBBfJa2MURgUaik0mNZVlGt/TBGspaN3Yeu3pYd1+DgbRr
ZbCTN1LYk1ataHN/lfHUbMzxD62Uq0muCjoy5XZt4aUkkK4Xk5pLlgDZaz7wtB8/BuwmXOH7FBOI
pWjK+bHHPIktz2o+T+VVY4g7Y0RULBtAh1Q7IKQbD9FK9dLoSfiWyAfsbvzuQYlhqecyQ17GxT0+
tWtcnyErnuSeCOCR1Tnf/N5/qfwZvv7urupv6n4dST3zEfD+uW4l4jZEeETRNV2OyfeEcxRhsAee
q/arefDHUwubwhnGa4qwlsxv68b7msMYnDjKwGLDKhWoxFA2kTWCOVwIEB7dChSWt5/beZiQEp4Y
pEX6yt2GD06DW54/7vnjVlJOFeROzkxsnP3JqtCiig6ZCzvrMscR8W+vLyYEuWCv62O0PrWOmwaB
w6TkIRK2ZjubFZKGmRzoeKiXyGXxmnlQv592NUnoK5oT7yZ9SXBwoW2UT6H8jMmSI4Wv9Yx4bq05
l7gJ93rwFEzTPcGO2Gxn5jjuoasVO/e4O40ySR/1U9GkunVV0vmzliK5bclPafErUL0mcAGWC6N5
651kPLF3meuko8OR5JFKoBFV8WYSTwdua784ypHep5E+rVbDBEy+azEsdmpjrZRT91/0semUphEA
mXNC5qf+jVJ7sDSv4lG84J3KCFV9UqpERnquwYKGzUhJcrQq0DyojbSqgRyDvNDzLs00DSYfZiUd
0VuzTwiMpBjIz2d8odUV2cCw4VIS/oA4WIXUn9teJNRsPYkDbkL+FABM+WvnC4Qj5AT25tIDU0PN
YeAscIu3pjgpfyf8JPRAPvcm4mWFnvekbKkMLFCC0jWLuoA/QXLNbOrlLDlxMcy0zHv51zFhZ5JC
qTKKdoaPeyRhK+ZHm09dVFOt+Z+Rpb6AXpsGsbWty6/FbE9M+VmaERfqJ+O8/Z8N9IjzzdJfPcj4
Nb2WRVZzPGByal7bnGSj/YiukBA7SXsl1PUfsDeZ8vUWBQ/gZb7VefgK6QnGkTr39f10AObrGa0P
w9aBRFYB6joi0xjyJKa2aAouGyrRaw9y7tZUkZS/0k38McWHVLiFUY75fpju8Sf5xoElb5FAWos5
TSotkEObFRrQN6vtmf/YVQIHPz7IXd4KAryalq1onTlgaVGAFsXyGQdqIIRNUJloYazIHJMoNR5X
CP0U4KzAtr3YoAaQKqN1zEidE3bbYbASuYwbAtyvwTRJpIqCAaE13L72L5DQ2Age118kZV+7A4ds
IAYjPgNBcnI4YFRd5QuJ6n49PJSVre3kB1JXUi2HnJ6rrhF6krLLw9YTq/ojmziHlUFjNCNiUFLP
lNUWOxguqmZC9VOMBVGngHHWa30pQLw9UlqqTPrnrWBnKgOFCtWYeJHn1dNl2+MIogclHokGwZ1V
owppaaDEpvjJ7LV2CNt/DG1B9eQe5xwBC78FPWuS27aeuSpXvMe1WRF4W2xELLnsNqHp3PM0BsV2
XfYFvhrDKrL1XSn2PBew0Vei8qPJMQJ/ICvsB7qsm7skpD4+csqjkZgLmoqtU3TnvrqNrayYpqOE
AdVnMDN94kv6gERYb0lQ90ogs/nlwycExs1MIOhrmQIAMTwbSkH7dBUibns55e3HQSpmAnmgZoqF
ahpXMiEYDz0f8yXbBiWIptlYFICmQeoqAfnJ2Ieo/jY3C5Qn3TDe4/Z/3XvrUDousfhp9Usm80e3
I6UkxmSpPYL+mAoFqEzWIBVBaZBAR5n9Dhnys7tzM4lXRzt8RqqqEXaJ10UnzFVgM6IAUK15Zjo4
wXvcciuMoXfSqomdPU9bS0D9g01Ui/4uZLZKW8dTl2WSbKRapeli2FOqDHyBPf9826ll54hR8dG7
oAraNsrnbQXeZmMTm7sdE3R5ivEzptxRzAUDal5mwYxRbQzJrn9FY/VQtKGWTQmrFoFylamf10oy
uoEtyjGNBpKs79NQgbSrbfU5KFqrwJWSB6foJqpl3dPFJbPGcw2Zrl/wH5JxQHFdd50rNYDurHi5
lVkDqVhhHVwxXsOa2hrkkkw9K8t7dwcE36BBocY42gfHhOGPXfNqsoYnDx7iK6a8p4arCh1cVCF6
z+MubzL8WeipZ+8gUIjDAymmzA6VebfUrGHV9zGvAc05Zo53mzpG1qDUjTYNZlQKDACqYIFCaNZd
LQ9xWQIeL7YGj1poVB3/S7TrMjMNvlU3+EtUlbGhAnM6/QrZ2f4DQ0/0CdJfHwmuh0nkDrfbzebR
RXRUDeSX0Cc7j+R38yHiQHOmT0k53aie9wirGa3o10ojaP6Q1ion+r0EVszYPMvwjYLuOgPSRZTP
2qwsDCpl8Lr2AXHVDikjshnLbFVhK1ziIX+yNrXbjcM0oIY+EYDbalVIhqQ6NSdCdJPLHb0tV63k
K27P6ssg4NjmYtWQR4gRllMdJqKgVnC3bZjb1ELNuU/M6E0n58NRUD6o1K1Sj/VO65UlzLsEuBbn
xIni1UEbW/xvni/OoC25a001SJC9EkkAClbixBmFZ89iplChGcmiOGylnGWZfjr3wciNARssUq6U
VUC0K7gJopQkDI+B+dVFQHoKpw9c5S1+VtJw9UT9mlnpg1zInfXy4QAMVBtUlwcTeMMdrXbTMjlv
ro3G9Ftme2PTqRMVKIDR5AMCZmKNfh17h1zJDKJt+iZgD6C1SI7SDRXCFOLrmR6gf6CA3guwzv3T
2j12QAj+WRXBD+vdMfhQbJOY/GLrzfk02QAZEvOdoNiqysSAIBYeHDsu2zwWqxfvIt85pc5dOG6D
h9X+GhhmtaxHkRZfZyDd0Rv6WVHi6XFs94k9K/vhjfkJsVY1cKAKxTlx8ZEUmV1a0elDxno4F3nM
M0dqUYadLc+YR4pLYTWaCun3usCVNc+OI/D9vLBQLtSdZe0e0TZPjAbvQ/3EC1FRj4kZ8pqIOISq
VJgLFmcS+7AQcO01Ro1/gSzcIEK4yBu5FgAcKTjGZjhMvzJE8GbvYiHPZT+92L2UQPg8Lay9Y7nA
o8JR067/bWbhYFJus2XhIBQYDr7pjRlISBV+cN7taFv5kLD+ZmGFcllSINihD3DSwYFnxVxSq2j8
Cx1BT7laPcO8FqWtbRCZiShGu6vqAgvD8Lubr5XTEFnT3k9nJj8SGvdILKYQLvjCPhE4VbBlbbeu
/Lvpb91fY9aIzXif8inXbHIG3L00R+h+U5sQrGgCnrPF2SzOtAg1dIkHRC5SHI1Wb6X1ZacXLoju
SDC5W+7Zrl5dy+eVdbKDF6hAiBMIC3ExeF/N06vt4C0jfYa2Fn4I49fBnZvqcbNJtYH0G3xsHvRT
YeHbzvt3uweiV+sgqq+4qVr3Vlm2F4yTxBVsmMMbrGqT0yOviI5NaDjmr+kLQrAmcjmmpMnSCdxc
FTmrpqUKQm/HjYSR8M90w8nK2vzI88zrsxYoStdzeh/frH0YqX+Qc7tzA7IgwEXawtD4gM+osdN6
GiopRNb5Igq8hJ8WChGkzPgbjsp1VyCcZH9o2OJtHy1vH3jqwWzC0sCcTXDy92KhatmNQD83YYW5
P8n6q7wfbGlla6m0OIVDuW+ifx6Cd9843yOHdjKNWseSyvqr9CVBMuPWqLc/fQvj8X8GB/RusKWN
j0fscLrpZceOA2nVoyHy2Xh2H0hvPSMZteHEgDwtpS2Ro48c1gGVRx4rZx9fy9/3sx5NgIFvlvsv
0328kEXDKbHjO4hnfJogK5eU37z0CTzbuMgbmJav/BysgKP0mVH+m4LkNfBVqLkfs3VhSMPy4T//
WcSy+DaT2Uhph1z4ya8VWgObmfYnfsLV+Hc0UrKMrO9iPWXzOgjQy7yCoWyx67oNSZoriSGH7N1w
bW/hMo5CWN51ZR7cC1RLdquWU4f0cIZDcFft5cN6C2Pd1jKEAsGInwZuiRaScnqJojx5twd/5mfm
RF/UORClWD60BZ80m5x90VZI2BuzA1XRoYSdt8jTwIUt6FJhcXc+MJnTDkDQhZxJYTNWEQtdBGS+
v4y2s9/kkMIs55QxE1uynBpg0C+N5b781IYQhhmfea6cjU4F9tUi3R1SxkRO+4lm40Y68zXWiI2t
SRvS4NspXwDETnkgPgDtsp2jM/S888jkbXH+tEWx73hnhgegDjRSzrVzdXgewNItEPZg32z8ho6I
F72+MhYF2DEMtejto8IKf9a7kSAE2ZuVK85ZOMNADJYZOyqbL73W8v75VrYK1rslO9zJwtuMfP/W
PY/NwNggtvfXPRMTwFjPlpykxo2B1bvvWQwHpmO+jR8Mjr3gAhRPbJ+y4M/1pfd1cspD32lILjxa
mEi5Vl8X6KBi+odszNalPgivYlv0XBX2E3aXqysLNdHuHgqBOHbemz9t9GvNZc8rL91Tpp8mtJ9N
I1FiVJiXJSJgn4OKNVCWZ873HXl7XoF+9Soi6hcwuspvHBxJPC6vzYpxXi2KMOlQ4MwOSJ6ykKkq
i0g8kefsezTWEwHn0tx13RAQFO4SdXMEgmibMLHq0ZEZGX2xpE4QRS0cDbnCsDLJHUwwFiIW3/OL
UDnDF6r3mj237Mucf0Oxfp6q75BNfUs88LFGnkFvGkHZLAuK/vee1bETgoyybIhqY2btkmXll36z
fV1C+FUio1VoSBGCCGXcDKAyu4cOYrnJ0O2+LN8WMX1Ff+TgMJPjdnRNZGncXBJFTSl4cXooL5dq
kJQ/Co3gUidpxqEu+yu1u31xCXWjxNuKgBv3LhdrsTKalzQMHWCTaeCowveVhZGJVlEEMIxxiijd
MphPobsqPYz1fHrqLGSJd7eQowTW+/QkEyTM5tRUDqUScuEqAa/bZQS6S5vb6xAk0EIV1pjja/+V
wFJcV05KgPf+ERHj+pwbCQ4NWVJJnN1xL9MuPpiLfZQ8CIfchHtGTLjhSoEY8GegnkUsQTAmYDvK
aZl69k0L6t6nAsIdBPAnIp/SLzanLec/V2DL08pQFrLB94cQiKno0Nya0OOJcmHAz8DLHwV0oz6Y
WvokOIQqH2xE2t8CROFoxPvw4zNJJFxJK15PTKPetgro+tmM9yxT2xTP1AaIHoEPRbjyH8/dgR03
ZWjrKfAThjqEmwAp++o1ljdu4kQEb5sKZXrzpsszHFmGbKNxUiK4Bft7GyugHnxHYXa5W23sSU5d
lEddB712soKFBuf3NYluBklyVP0F+Qrn93koOFEHaH2II91w16dXzgBnB9x6YEIN7tD302fs+6Pp
Yms6Hnmerw6Wtcs9WxdbqOVuIatiHC82HFLDKT3zBdEIap8hP2F2tHDrYbHRaVLElIgZ15PIWkI4
zwkucRs6NzmETiIfoou7hUiqzV9ateeKtVMnA1PiKkGChviojU7G7gB9s+lhAexUcGhCQYmexu0y
D+xEhJGK1kGZ+eGet+5GSc+E9i+JSlHtNtH96MOfGaUbyl7N9xVcKRqG5f+mMq2+/pReX0GKAWUC
0vo4vf9Usgo+gUa6yhUhoNH2D1jqAMDL8yxEeu6x8Yneqq0ZEruQmkKdxmGAeWCUvprh6axAmSzV
DilIUBtbKa2+D0hwQ+5da/XfbsQkMWYcSfweiTbPwCWYTnxGwUBVSdLikc0OYWq7u6Qh6w3tdS0i
+M0W9VADn4C7ZjVCEuNbZGbK3UW5QJoA5UfqVqd2gOCkQalgZrqYPokBf3evlK8D5uvkSqiR/cN4
pG/t0TWIY5Uu1BsTiyKaAIZAuII2DQUehY02HluikqlS5ECuX0dZLi+mtQ+OhGkMPrGoZ1lxU5f2
nkP3/enB5yU8VcuFA/cGM93WS+n9xIPad9U8kOVFJpVOhOX80ZspvzlzUIVX8pJlrX4niB5MB/UF
gbtJDxCFu7+QJ16ukduwTV4BKh4g4KadGC0+HQRyBTtypyjfpFijpgwcp1ydWu0zFNkctFpgAa3F
EYApl8cMO+5HrZYMJ0B8eWrSCSoUpMHL59DPhss+EIsxA1BtglsRJnOyzEpZBuSrrX2SIl+u/YDa
HWb0zqCSKxnAEkraCRocqp6KFxUWDnTHIJJO5hEGQtNfL/TIEkE5tnfVsXTvtRVv6ADvKEJ4j6JA
rNTijegRVaCx/0AuOD0h3dBimH6df3kblFZiqNxuVRQBSIy0HMwF0VYx4i0vMB9AhbANnfyDKzXo
nBvFRTPeBFI2Y4dqV1ZmVatC7P1MpxZk9E19SK8HoEkabKzgSHgXPj6Ef3lsjrg+zxBUWW8UNNXE
2bD620xBJB6jBrlcpZBQsOwLvbZA0EiK+i7rZn2dh4H0xj1V5SCm5nAfT2KmINYR07VNU/2ydvsl
QvYJ1Ba+iHeTln0IOn0OpXuzjI2LotXhex68BO4s4Bv+SIDbFC9DQ5Bgo7wJZkkpA3X2Jwz91kHt
F43n8GjjBE+5xB5rXWy3hbYJ/iK/OQ/SeI4o5+Lqaq6FkaLt2sOrXfsz65e6NcK74NDb2dS3G+88
DNUTKrLEYhmiRNxYEvYAobGC0V9gSk3izEzycFRPO5yjZF6l666IUH637/l+v5Q/I8cJqRf9T41d
FVuem535g2TYTZKrZWhFDRtZpvI0e1unXC39B14vj9Rfh3sLHLsBQ5seadil3if+x4ak4HyEB7A5
wpYJTYPBGpyb4OLCH/i0/HWdOYsbjJMOhWRqYmJTb40KLz4GPvT56TCeyty1QPgURr+hrSCMapEn
AZhwzH4y7TvC1MO9CojQN95IBWOY206aKJHtnhmBMMNko60y/KMnBBEInZuXF3/zSUXy5SX2cUwD
FbY7a4ZhV+3nIVPja94OTvTzHTHF1G2BmfaQLA0q28q5jr+IGoYjHf5f1ZhkO3ISHdoUfA/3OIZu
2hRCxIKKaOE9utlmkiEDxhe+WY7WIylDtiOaavGkw2/vTJjimFtGTEg6r4patNdV53a7oSwUIF8R
RV5JLHFgZv2EeUlErg20NMI8OXEOe1z2T+8muBni9GgaAzYWfpZtBG2GQQ6AurVEi5ZnINcE+uLI
gxmYzDfrBng+Th6HDirzNvLnu25q68MU/TOW4zfAcMV7WYuVWiJ4Mtm9XuzSxq520iFCkor3TEw6
KQ3stWWJUZb8hfFJgzbOHbgrAzhsF2zS77Cz9zQQrZt+6fIz2ELfDHWau5E5sePG42Fnsgtsc9mR
tZ2GIqfOFLj1E6YvJI8OdqAixDEUOCUGfEgS/51Olhb5lS0hOdVdWPDBIfaBrWqraQsa52yLlKrm
sgMQ2bYJsIlEiAk2kvTmI+HHshRHhygO0CyiLC0q+eDcdM45qbAHSTIdyHa+CnyeoHEp4zfqaVj8
nGfhyXGG+vArPDhHgHuS2Zwk4b3bBV3x8OiqCZMhNNb7qdQGhOi4TfVSwMjWlnlrErb3M3H+keZj
e788Za0dvgx2zNScKb31+0IQrnf6pvXkpYfHi+qinQ2DFjmTzxYUoVyoRz4IpM5AUsSHEDJriq2f
5/BWoXS+2wwORP/yk3214TtGRJ3AVdUbdoXghArsUg56Nblbb1PJ5Fcy/xoUXNq2uaAo/TmgZnbZ
AFWqbmxtTf56rIvbJknLDK2GkU8ZVelKykMgrg5DnKQajZDtEgKEbR6UoYZa/KLbR2jZBsuI9Vm6
eXRNhUbXJvjmjKMUWlDdqekCwEEb1kWsFA2UHCxQmhzC56r7v4/dNbi10qvxiGctc2rm1HgrTyBx
r3X+hYDL2zLsiwF6pT8kWYgrcRMUXaCaaJNlOQmKH2xb8Kf0dmOGqJX2hONZuzulq/iITUARJYCU
HIjABzGI6BfVRGhIpx2DwixNI+V87bywFgS/WLPMHFXY9nxe0V0DztcnUa6xwNAfR9eZ7eTba5QT
GSCamVMgSCsUmwBlZmQVo+Um7skBwB0kramlKeCYv1i4CsipuJH4UzvJessqxwoEgyhqNlzRKy1c
gG9du8zZpTtBIza3r41CQBM5rEyzAFR+YyplDOBml72f5oLz7yXKtZrL8xLRk6Ypeh66b56vE8vX
9WZGIrhXJvH5AvErKVvfAuW7u9zv7LzjOThOxdnr81GmZJ2puES2vMUKKb+2nXWaSqoBH0qLjY6o
rA==
`protect end_protected
