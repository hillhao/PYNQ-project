`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aE0tvinbUqvf5G8iOWas6gNREbQuFk502egCNjwMc3+6gJd1I/BMUUOX5qQW09U6Dz5QTjdYJeMu
BdednffRbA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TxHuajnnriiCieyaOeo9vEVhhF6E0SlcfsloChiDnNzjEUcYBpuq90q934s0YN7gjbNB0y1YXP38
pO4aJVjVDHtgQc9hcVKRWCY+SLmm5NBnnvyrRkfa1PktkKJTQZj/2gDjcjMMkYju1+vwg3fkU5nY
tsiE/5oiQtekBd9qRb8=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TRVYph4LWhyYSztF+Z3kg9/DCgkRHkIxQd6pSTadaFLNK1pvjGVtz0coatC+8yBwXBpX8qH8pzgQ
eNtjZnHnmvvppsUnB3oT6GtHc8ZbOa5d2Pj5SYg8kq4qu1uvfBeQT5muEZocwJvcgDBZu0eyl4w2
D4nfAZ8n7VvlQGJ2pBU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TjdfrWruver+LNuSAogn8BUyDQhgT3unSr7d0ijUBW1pudWt7H8m43PM8C8F7GMGzoWSF/RwCRYt
K6EugueA6QJd9LwzrdeAH4J/7I45u9gLMWiuuoM2cxfkeA47taOn3YjbGhh7rRhDVMMDMGl8lAts
/WC578wsx7/Kx4rPZCFeJs7vBgb3/Z7cWixNXgXGe3fG8S/EqIPmho59+DIMrDvuoe6+2+duNsqq
FJnSqNcVlUB9kG8hH5hBVdjojRaG+WQRK1rxYjrP64CPOq1e2YeEjjObyQtUJlHZY4+5XnuuWNcD
IxrY1SFnW9N8gMm4+A9f5tk91IVoOBOR5bjHAQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dCaVnjYyDp8nNCbNOvnWD0ph47Hfz6TwHBWBIT1D3Y8I512RR5NwO8EaHtEllb0XbPk4RlKQUeJL
d4O56C3Xshtj0ztIeOCB6w2BGZ0ZEUUwLdxV4+uuCxg61xJTJbC5+98CI9c/dtj9t2jMXzOU5h03
9MP5Wd3x9jbAVoP7BVdxxYS21+bHd4j1yGKAyHwF3+Tq5hhF2BCYYLhowUHMA4a3WtlRvpMZybEZ
sr5a78W4wf+yigfsrYc8n4VIXH1K4KG4ybyQm60HF6fAQ23jiveqAWn317Lt2qi8mYhDGgrGYBXE
1fQjLr5As56kCk+4ZclnC+wS/LbCXoKf3u77Ow==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DjxadBnRj2ZC5Ujr1SHVkZRc/Ios5hhXUgItDDGYCBZgSlKScWNPNwHjrjJo0NYfOqYSgc8VYsZu
JDynCsDDqHNm56VKSTQwfXo1O2TPWokWbrgHHPsQYSZ+nxg2VdkUbeg8Y2eEXLHF67iGA1nOj7kG
R9cr6uM5e1CRoCPRESTqyzPE6q2lSlRI2BPq7cLUOotIKiaxo5KoUkqQyzmfC2q9AfbyU482iOG0
UJ6N0/Zwdh76iQhF4kEqeuNAA32bMVkg8FlXyKyKTGdVOtMJaHYbMZSIHPc60uQmH23NdbO73ebD
cToEBhdGO3wMx3ZvsZDMGkINdTsfEDB78KoFYA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 114672)
`protect data_block
Nc8QsCX7toNDZag8DW98RZEWogv4xfDtEiKxiDynQgkUIxEQwWFhhlXMQ5Y+B5yO4kvsRpcyI5E7
gDmjvzcad9V9qb1EYVW9VTF6vGm/ngNPtBKoOEBH/Gcxyx5DjHp9T/DMn8yxSv6jAlxg/2kwQeyP
sjFaeVmFfePLcxQH/cBrRoSXH5smdZPLzlU0w3Du3Rhc2s24RVUqz+gUKf07eUtsa3BBAGPQ5EWq
Q9AsKKfjwza9qVBpvm4zkTTsH/75dnka/skc89kG92cGKx6+AHBYzv1QUX6ViDUCVUY/KBQb2Oxx
FkMAzKD+Ta4xh2yN2NF+FG8iVj7gJlol7v4uykNai1IIQCWNIL795zRMvZR7yYoT2pGN0Nua+OsD
boc9D09i7cY8EUGaVKh1l4qk2yqNgP5kUzJCEnXO+GmDio61NlAJkp6FOk87HvGMhsXniGZ2bKPv
ci7OczdmbBWm8joiqYJSlWib3VnSLMMFDlD9DtcuAWIfTVUnKuUa/Xe2K+s2CswUCH96t3qjRW8t
L8FAfY74z+U9DkK0k1Lvq3ac3ojb0sN80b3BzHfKIglhV4NxkEqs1mK9nx1lgBygB1dKbGj0P+LW
34Ctkw3to0pANntqUsPG/489PBIgm/xUpLCKHRwKTruc32buvxLMFzjTLf8sh/v2+oaFtWAm4hMA
FE0q7Cj1m9CNpPtB7j7hKjYImOhn4kBeVOVPlGTLfc3eA7dAkAopM5AnKx5l5J7j4OuEf8X/tLHO
v7r3V5Nv5IlsMJ4hSjcs8R9EWoCHELOYQyNhoit1v8x3N7/ArSMRDRsr02g2zTScdvyjgEXJ2Zx/
jRCk63b4Z+BHRtHrd86ez5/eIvY8Zt8b1KfVDNKO7VcqraO7grN1KIDyOW0d9PeCokTirZ5Px4du
Wys8d4qWaw+F/MC6fSSRjdEiY6jUt5eLIX/L7u9Jjhqc39eY9D/vBHkBxApRrb7VzrIN+PqytBIt
tzprtpSzF4JFgHvTOiSrMqfpecU0vY8LuApzyVqv/KyYLUejXSlOCOxwD192sMJ/sUSsaCsRe9Sl
eabrr9Abt0TIuXDbc/bLgOfc2b8mvv+ezE+aJ8pfV4d0xlqsbi00aHvYNarN8qsHI5bfj1ZQCR43
nWQZq2/1oG4L85QiNRheXVP0x0vlFAx4DbFq0gXhDIGCicbFbB0Flbh6LCHrvABJlIVeQkOoX5Iv
PwOEri3wzQy1zxzK0YgqIqVTSRf5bUQjP6b+Y3/+2YfRDoNVq/laUT8QKqXV+aLctEKMJGOs5t2i
v6s48d2RevqciSXpLvWF3BvtVI8jYkwqGNCZmxNcgQFYVOo6Y2UbaoPdrX4jmKNsY19G7wgvWsV6
7rXB2Tan1qEejC9NlpWbfQ3YgVwB+QKPLxzCpwMEO+4aCIgb518b01z34hYneVonhnNRkC/+Xcq7
YYfUICdb1joDJRTO6LkzJD5fVR1fiEssSYQV+6Y+2iu+6D1EtKWLdNbN4FmPj4QtSIYk5o2idJOI
jm5NrF9fSXXJxmP0iZqC4Q8THffAiZSewLTFabSjkfr11wLG59J6PYkS4CQ+vjnIIh20ioSCSGBp
qk+ffmpXe0dl3xxdgDH5AWo7ZmMa6u3yYdTEkHYesgGhj/inLJNNEuMFQkFRSbAYywaoMW1tktak
T6c6HFLvFnx8dM2XxajnBPD3Cc5atRiRc/7UqlM448qSD68dtC2rUuCRkXkYAWU8iso/ToOclTEm
7u1VZZGBe4TiPCMezZOhd2fv3ZK3By32+qPRjz8KUbK8R0kbjSoyHzaNk5PFG+tLA7mb72z/GkCs
S+5bd5xOjRDHX2KznJ4rxTtDpo6VCzlV4A/vJ3UA0+DL/pbFH6ZIpFAExQQDvLs22LQh0SzVwOyT
50la0BRquaDr1JAXdEvsHsa0o1SDmV+u+8nia7AZz8xVNY8SSQGbt9+2X6dw9h56KwSwArBnUzyV
F57LgiqTRhBw/7yse+u7bW1y6NnbKBrAa98gsK1H32jhae11IPppPrcDTPYuymj3QEsRsDjoHImv
NuS/tYFpO3aJIN9DeVR9QrGCFTg9yNhW6jkvYq8f7Et/aPAEWzfgO8Yvggpa4ot6PN83Jqh/wFQZ
GzRutxXUVfu0sopR/x3HaE3smNgtLUWwCytEnAq9HN0FgKC78SUKCCKV99SScNet6UtK9OhUZF9v
H9yb105oIsdf3cd633XP7jVbIVshMlBJsPpaTOtBPIABobqIatVSOLR3nQZVsx4Ruh3utoyGNJ+H
6uE/NDayP7b/ApEF0r8WrK4iOnm8k/eM3orCDQm/zeYc7MbZatnWqHEhoRtjKElU6uWrI1XyZMvi
9/lFAaWn3QLn86iLdBx2cOq6u9GG8UsaP4u9IWmpSydlMi3sNtzFvhFq49jUNkvhf25y2XH01MxR
4UhJQJ+HhuyYG8HM4IngfOuN1MFcm5kB+1yxVvNqB2DU13q89qgj4KAa5zzuIwGZjIhLjgS5MxfT
TfK0Iv/q+Z2lINW671wQd/HJeYGEc8tvNu1JJoSlhoEKynP53YlG1wWQLO0A22ixaTD1P6HAF5Lg
g8TnaIZr7nfewTW9QBpMR0pA0C/My/fxrySt2QXByD452IS+yXODcyeqbkAuutgB8hrnV8aRM/VA
e0naIhlQ2TMOohWhn/xvH1V22H6QKRV98Hu1vEXjccpXUfEZUw3nBwhOu80iY6zmu7argxEq4Nqs
P9qW75St3h/syZJK4nbIbPDX/SvP1x2YU7gn3Ua/E+VPqJOScIC41tTpgxZQPkS6RhGrtnnsYcMv
khzvP+tGUfZWcxBMdZ8z6Qq0cvISoktBvomksqiTYcrz+6hiAADH/6K8curtPw7l2J1zXGooZma3
TJoieCwr19YmTwPlgXyRO2guxlqwLZ501Uw6mlYj0P3rT3qs39eHmL94ANjl0oj2FcbXHaH+od0h
Nml46iKmifNJd5hvHndLm0bOWUUAeYDJ4+a61moCNhSJ/LaDFcy/GpA2/oHaqDQOh2jaFKGBWn9b
ULhxHwxxpd0wpDxjrZ0aG/aCgMKnUjGSFQJC/znZySjIVW2Qg+pPjSIO6A+0uVqn4JXCKcv44/Yo
CuAG/91oymsk+hgHA5fWhd9RcKf6pdlmo212tEo8yTm/xCW0SlegqWTshA1DNyBr/zh68VJbC2oJ
/0T+dqg8OVq7SkU4mzXJvFSOjcYrFGf2ufgg0S/56M5/8WQEP5sZwtSemh4s4YAjB+6K8VwW5LMh
k2styD75Iss8246XrqjR4hhGcqpRKWWs3oQh5jOwiiT/P8oere/3oII1K91vY7ky0t24cdMo5fT0
LguY5zqojEIbWfBQV4dg44OAdzxRoVvxSuDX777Z0Dy2+7SVelbktekVDCCBLio9+CUG7gHdYK/Q
NEhSivMZWeq2y5pgfZ+3iiNZZyZFZEyOI6mj6aBkasVkfAAR54rPMvJoHZQ4a60zCsYgwI1ZNKEq
TknY1CUSJpxQf2mdgjbXPCoZUIzuS/NPAg70dMyFOVPGYhrUmNXLKjRjKOf03rlBV95BkofkecVW
HXTZOeCJUaM9ICFaYIUfWgD2IT8vZPQNbJrhOgutARqU1D7RXCsx6FP65tL73YckGZJwS5J5TQqo
WOg7QGMBRJdyGY2bd3lH/GqGr9BzFlkrCBlvzPoOuFm6JdTuZYOlwigNKIZu1qCK/dTDqNBlteUA
bITTC1fFcrPokMvrD07/noc2IgMYUf4peG+RPLJDgZD6rlSloFh3VItOVp589L27+pf4AmJQG0t4
SUjnjO1lqNOUCzEETmGBF6qY0WyKToM5MTX2xCERMMw03Cn07HHH6lW0yUF+vWQPNwlx3g5NVZCJ
b7WhrrWdX7mOC6tsn30VpKj8OeGpwUNEX85N6b5hF17uiGbkX855UFaRNah9oGUkWKQtq8IZtqB5
UYehyhXl8i65Jf7sJgPOLNOUMre8J8/QYDJlqRZKv71xkPFWRAPtlExwHnEpgwmnVsLm1GnufSIu
sQAiz0UZ9aOWGYY5XlWRzsWlpep2h6zEHp4eXc6q8Y80vIyd07EtpA21APnBAkbXpiDBIYsVPkUz
NAVOzjeNJGVdHdapejHu9hOOFtfwSVCLlNVSWOpDj6GFbvgYEf9uc/oppYgCnyHlj7/xBs2HqvOc
lI3dAEufW43/Gex/fMyxMB7VJA468ELeEq62sHmkFV9Zb3VlokdDj9PV7vXIeEB4ILNwXligJX+R
ybZdrzPOGTIXdfpLyX+Ibg8zWXysY3GLCooiKNpenE9cZhoYrHiqlr5vnystz5jyosBQe2FUqXvz
kZoUZwDA1zvw8PIfHbvTMYD6VSroJFonUCwYbyLFq5mqa2UsZOrs8lYGRYIkYx3E+NOq5T0u73T1
1iZBD6JJurL5l3DZlJ5SwjSYA0qYTN1qeSsuKoDhMRtDza5QIqMbbqP5JbAZW+Ym46qYz8U35tG5
j1yW4DZqwCKt1AHMAN2U402/EGpAl+i2a9sioYyHFhK7janD/dfJJgvjSF6y+VVDqvVBtnwdCNFL
A/cyFQnErWIZ2ya+XSVWIZW3dpx6tCVqnpPCg9360ewWW3wbR97QAcpFzl6ohYOc+e92kYinp1lf
x0+Mph0qKp7k9xvV/nx+AMm9OxGYyP5/thOfVPuGgSE+tDgIIjbU5TrfTwA2CoDa95exTM/goMyU
UzG5iHWDXBwpCnHxScTufTD1zklETAP86vbj1Yg2dJy9PRjcgDphEHra/dDc2lV5Ts733ExUA5Bp
rXa1GQTLBJwaClZrFLJGe180L97C28AtlwSyV+0ynkQ1bMBKismaDA3gvKxyo62IuTcJ2aX0/l5I
wdtaRW97c1lqIuUGyCUTGeQ4LvYHZzR25JzyHfpxNO0xmvkg4fWosaTV32dscWFhs87O4qqqgnna
XMdCoYQh7dQr3OzzKhq4vODpX/RYIepHr1gV68Lg3u1FI6jkrY+C1dQBtHlx0XcWaRSq2A5EbEjQ
4yGED7nLx04QDHHx4l5gXgYlCZLIbeAct70m05LvJGF3yEdb7+vkBHPYOqiAhT8BKoD28vhonJxG
Ao372HvJh7RFqmatDLrGEvVuqBIWBDxFiJYJiCfbf5Io6hYESl/Xdvj2RUu+iKZBJvjz46hymfrR
X+wpb9hrrVmWdN+VK+/a1Th2pXts5HCMmuVkVCbEItK8jxeEkkCg2KCe0cHy7Px/DhCF9DC8NdGB
iLePMAqgnm0V3Mam/PWZBRc31g7wzJZna0QJOJWIal+Fwr/xxOzz8IKq/ezkAGhNvOd97kN88dKA
uNgrJ/01FzafZPo7tVgsQCf0rKYh3sXDyX7iDSNJm/Jw/01jljgLCQHZue8QONZasdQCDVKfFWI6
wZM6ZHlbMRAM9dW95J/hKTG7yEgTdokwd2LtvVM/dXHZox8CONC3U/JEwQdB/qW+E1ghp2Jwod/4
ONvTMvOnUbx44IB3GTB0VtkYsTuOObZz+65OLqGY5IGu/G7aEZCBrLjhwKly4NIwjeSnNQr/3BHm
VKfE0RYNFLB/ScRtTXmp5dygTAIUWpdvPYEPvvYP+LOJTE43BpoFNenC0OarYNpUj/HSqK5KKd5R
6BLNqcYb2/JBTKkzo3FuSM2T580sL4nVu8utQuJVSeWdec1BX1DQvBlQ5WLsnpqi2N9GsD3JhXwO
ysCyrKNeJR0r3VZHoaF7pbszkXgue6SwCczejSJgTdJiUNPlBMhQkS3lpkbZPpFTQfyBfbOY8pmi
QKIoXz+ElmF+bt0qg3WwX7ygQQSS3knYv4ulVC7lvSIA/grxLtmy85ccEn76XCtGu2Vv7WbzeuEn
nEF6ybMOr1G6ZPeCNB83cFQwQ2OF3n/5IWVneVA/Mt5xlI/PA4JOVmtAFnyIur5oWYHMR7vP46jT
mJeRzML+UnK1DkGdo5rCOzw0QYxhHNw0dGTI2DkSdlgH2r3jkTOglauAOSoTgtPZg2Xn2GyNVHtk
OYs+9iUyO0XX2FUC0DLgX6Lff/XaiVbpBLiDKrxU+RA8BITCH4QvtHqDm1OnfrT+oDii32kx4ET2
4CjX3gbAKHsiA+6LPq8GbkKoHA4lW/rlHzU5mFDVUKx8g8/f+kZpdYPky115Vs9lLtXbl8pbBLDR
UWyn1KQIYj+8aCpJCK+3gOhHNIPfeLUYkCFBs2pNFTonncDNV/RcAU2XY1FBdIGDZmk2Dmkq/5ph
aMcHD66CS9BmMWOSr+apYuXPZN7fH0Vf1YvduuYV8+JDl/mTVR1OoA7M26uvlC2d7B6r//SmN5MS
7Rsywr4YI4TOh0FfHteHgFsVnwkT2FEQu856n8IMguE7w3Kd1Ebk0IiaBevRdFBOEoRMxbq4PnFI
j/Y6bDaEPpk46vx+ye/g9cC3loRGRmAn1WXuB3lN6CeDqQ0kZOJZS6alUcAm80zrMyhZ/F8ch1S+
r09m8+8YLsSK78I5t7cK2gK6ycHXeQ/xC/oi5gsdq23MzWUN7Gr+jaYOIhgP33DlXL87wKVwrs9l
AUthNkqV8oW9BNKfDv5rQwZYxKiv3B68EGA8OIIEm0Juea2tqT6Zax40H+kgBln40U/kU6q6a4Js
WjNW/an+8329N7nxUE2Kt2jB2Hkkpqbh233aF/1FesG7C0a7PSg09ZHQQ77txtTCx0ZzF7Zmwsal
mRlH5smDjIwCq7nJyHvCJWEsHgjoV10LPykKpSzuIYNijooIeNHm3BSQ/42Z2zmro7cGo0j+cDqq
p0+TRN7MjlBGFMGvo7++klupyDHmY3+6c2pR62Bpdx7wDLl1bJlU+08FOGdbkJqKj29aZaX8fUFX
crGEtPgypqUsojvmgXhB49M8tdZAEoFIvtWxlGNo63Ma53lRr+AbQq83j5C87xpV4Q5GiDaMjvRu
nrhryWbQcYCKVe1WA+4iKDfd2hxMHxqRCacuAX7aWTS+lVJzS2CI71SvFWP4zY9L/d+eudNtRkDT
//nFLIdnnJftDo8j4UrlYy3fUlpelDhrD24OxK7v5IoNt7aPUriDqhid4oawO8S+sXDK2NGRSEQ2
19sgwUsLErqnpWaXIdkQ8OCUg56VnTCnEj339M7Exlacb32p8m+71hLu7JOKtiek/YG/f3GfZ27q
u/+HDSXCg8RjxrY5m+TH92vmBllRNMpTsya5Lx1tXgIB86LgnngW9XVocir2/e4oYD0YuAel4NK6
IqyqHlf2JiMTsJ2bI9J8eySCZ1k6fVE1P+BjYSRVj2btHSF0m0bNa+T9ib5bNWk8E3ps+29+l9dY
S/exm5B6lInWieIhlvyrlgrSsBlWfVWwUjlSast/vBwYLaX3FLNttj6tvQZ5tdgJ9c6xJbrLJa4+
WcFOtXPfTlAnhvgLUHF3YvRFDxledEtIH23swDf6maqq1YYTN4JyMyaT+Pb6zMPJpB179Axwq/Lu
SaBrVI2ZGKVMHATNy7E/ARo9BdsR/f5UjRtzHBePC2TqBBINo3QL5lBNhALXxHj7SVVYAYZoah/9
/lJNx1EzxHhht55978KIEOCWAVu6wcDL3Ad6CHX0x6nD90BrwDDhfkZVjxG7FPcI3yCr6A3/3PDr
3NU6xCFdoXcA66f7m4CcWeF//ifhh29snHEtnDARkqjdvwbwGvwC9cbYhQ4/o+cAsBG/1cZBRDHP
bEXGRIThsOUIAMykS9sUD40jqOcf7ShFbCKTVXGuGGAo2OxO01gw/XBc6BsS6htMepLfiNvCSUey
6t2WJ9pv9OQ5Dc8MzbIiP0VuMpIfV6LHIRsZ2b/EByp4DHHMlY37HKS4YxaBPpzYZLz0kdPbexyA
++AhQQweL5P3mZvVB+Xe8hnoomim04aH3dIiYl6fIzE7EG7JIGLjgeYfu4ORMEbs3KZSAnpKeF39
pqJKWRM/eagJqFhwzAHcxnrvmONWwOJqrFQQcz8WLsB6EHIHvHUZDq3dVvf551/R9VdHt9WMnZ5W
fqUAe45OkMXEUWYNU3D5SC6v159e5DX5kEupegJDYSbkkW68wGDKa2941DYHreYMHYcMVNUu24te
x/53oM1O1kQ//NNN5f172PtFmQRWclg0LlJNXzPr8gS8XDg/wxasT/MZwdEeqZBZ057RoCks8UFn
lFwU6r1pgzOF+64DY7fsJlk/AGL+gihiXiCSgtQ2iSAvhvZKF2tqiyyFPFmDH2oWvEqixF/6EleN
nrKyFkUJxGOLZ9zNBtCvS8xz8DLGOS9x4cYn4ZWEOzhb1ZbHsTH1h30Pbf317rUTWpQKueLOvFOU
hLu0ADyBHxh7Hu8ZpPSFWge+cMvX/OwUWrP00smiCKRngPhbKjwjRkEpeaRRwddnqLZMcb1IOuKA
WQOyi+Zq7JSUUs5xDrHf12yFcu2vE7sa4MWFvxnZpHe7ucr0ZE9G0JJjjg/GVB/E+rpm1sqk2Ek8
U8mk/uRCmCcQsasTGBs5r5EiQjPwj+qBn2jiIcGZlT95oHI5FCSC6714Wan5TSmyN9UV2j7QRAR6
tjj1UMC1tZiBk0+o1f/Z1Oj8BZSs2lwFgedpyS5Pz/l6EqUTv6XzBklM2gyY5b88tcaPuiZU1UWy
8qMH/+McLWbU81BohXvPYnLwAT6PvuSvZEGkiKp7PZl3uQXXCp3yqi4/HbDBTT1rNX0KO8y9FnGd
GBprU+9O+5CRXoBxZRdxv9uJIJHFDU3Ty3MCz7hR70+ytchViYi4XzD7xG08355lYdVmGF0N+e75
Crb6vjzTYUXnSRX9IlXunjH27IFXw7uk4Nc+xWshtfKWS4+9X+0CnU5JhrpV6x3vI/I1aSONLieZ
XeZkNJj1D0NkaRdBe98O67SJ4sbWesn2jGMlnP6QB5g5pSHhRscYpCrdz0mEOokxncUOIKDGiYF4
YcaRZXiUSLdLkgh5E2uHEVPCiz3r+XXjUwX66l8m1qHdP3PGGMdnDf60+aaAQ+JLj/XsLr1+fIhW
31e4MvyiSHuI6p4Lcu+hgke5vsUw1cIGUG29KwYqLCDbghSFMeH9uivR6HlicYKVatGIx0MZeQkF
JiKgQm/gEqkFesunhht97XK2lBofS0CBiJ9rLR0QvmbBOUf9Q5j+nsqdDovZX6UtYIiZKlxz7sPh
mTG5p7DqKwDghYEIB1cNK+P2ZfHFXcYj9mfHIZoVUz20a6kCVbK5R05s/xw/b0Ve9M3yDSWZHlq3
KLnVXSI8UVF0tvONGLQ/zfjwPS3oUYTL7ZrFD0cj2KG2h9dBBVqzkfk2YlwjEJ4NkW9tZJMa6gau
2s3Hy/QBGFjtI7UiEGDuSz0f70cXGrXBiLkdl5Up1LsfAvxNzRH+DzY5wGR6loZ0sxILH2jX00T/
hlxlKQdq39jZY11RBNN5By05Qb2ZuglmMMfzvamoXvXtLk0BBk3tyRX9AfNUrPtzhnFQIhABFbQP
GQ2j0BiIKJA9PLD0ScCd8MUSAJhZ8GH5z33R1jKuw50M9mjpDMBPJtEabtgHmPZ8w2hkIX5sl3Xw
Z2KCz4LxiAELapX11VeTi7GmgtGcdNQK8LEkBi7C7xQdSnuDZOnVPH5QO9+UYb7hPYWKo0k0SguI
/DSH69sIK1OC+5/idLjFnsqtDuhfHJkpYZTSO1x9nwcwu96KoW1mOwpcq1CH1J/TLNRp2LbkMrXg
GHsgM6woKNCgl9WEITOdzVE41F8xPJfRuvHaBwy58L7qfuObgEcIKezd/yCnb4QrXYTfD8CvNfWn
FyCRKNQ52h3GI5XWzBMDcudYq9g/bfDJaPpE7yiDEcw6vAFTYwW4PpscuozDJY4RcI+gvtvUsIsD
b2743axTXFeM8DBRNNd/lUT7Mhj5h0eH5ixgx3YZVjTn31z8otam4I0TFTUbXU9Lz0Jeb7Qyxf+K
lDEJmI0AuqVHtvt+Y4eDftnxRepinPXF3KHeF2864kR6ZueCSr+/7RXRHa6eYW3X1pDEsIfHHsDB
FpfVgRpcyPl49jUX5gyJ2ocwysJevRNEGFf7jGPbPPM/Mdi3QpNxM7D+Vpxu9DqSq8u/xjy54RsN
5FfX304a3B+jM9LUusgzVg/trjSZSrw1QfiA/WgLN8pfet2K0r+bjcOCXQIcnRnMYqfR0qs8l0IY
xKhtZvPXrDMjWnkYOIpJK8VDcEDu5aLgWCJ8hyyjWnkg/eM2QccyQJG+H4dqgLI7d1cxnvhpixvq
wh3DkCEVKAHbDG7xwA8IV0GMU5F9OY0uZO7l60WlGP55G1kiD10J04onVKHlQ1M5Eh4cRy9Om9ru
Zuds+hc50dibMjnLWn0STwuNJug1SDSD00Op6DorfGxAxkrZbx5CEkVxq2efMjKWe+cb88nBD47s
pvK5xM954I121ry6sRAxEGTyXmfZga4y3e9xqnmgqalkho5pG+owdTyeF8qFro8hQSNuErprf2NB
Lsm+ik3ZI5NhcfjNBa1ofsc2xaJrIxhLZNz8ht9CAsSCZHEdmFeigjW1NsB8CDLEFCd+3/RLDkwH
foZyPv9ya+vRRLGgZNTqGAh4COpqEWQyuobEZMW/hRHy7Pw8Zw+Wrwl4peElbl91p/mAPHuwqYYY
1wCTa+cvliUIDWFffoW3SOSrig/zy9fSssOvwjxZYdgQ2zu5y2Ni6wRcsXsTWVOGsDHsPgyDqsPA
ulRWdvBRI20U6DN6lNTdA2l/+v2MTr+9Fe80nmS9UHvGyXSwwHGm5oDZFw8DQaoIArg4cEq3uOet
EcFy+krAlNPQIW3JKUT2oV43d4E+LYLg3AuTSWIs5uPNLhIMr9HCoZ3PtA4ChWNJaa237R/mKHHZ
vBqadLyQI2ya8e2St3WqumEATnurBgAgtNPXT1p4vh5y8vNLyiOgXCWCunClgv+++rpE2b3lBEIM
U72O0WP4esbTcm0RISSzcZhPGgPnXcJrZ5TsHs8ebtukqzWfpLV1sDPMp8GKA4L56lgrqVDNqsVK
uFgKKYmAUP/OAu3264t0tJ8NQQsB6MarbLWDwsWbJZoVknBobsZ8LGUT9WCyKPZ7M/0NEmSghHOp
mgKdjRFi4jOdF//a+4DXti7nwACOVFUToBWnMk5hOwXO33wbYbrQYDax55Vq8YyJksIGeq6QH+rE
FdEzA9obGU56VfYGV0QOY4ZEIaDgpfq1ZTSnCKpGVALETQxegT7MeJVkSUq9xtflur1gAZfTrhm0
2z4J5JGAj4LI4hfrBCafxihOwWXoDPO4TCFJtQP+u0JfXfEeIz0YWDoQ4okwsHH6DedyxAxaYFkH
HL6h+HTVXAYVbhI8YyttgJSCuX5EQ0WTJQKVx0OQCW1kae6boQu+LtTVUmMqzOYHlHEfvTy4POX6
+dE1GWdrLA13aG9qVZ0sWVecgHau9JH1hsfk/cUiRZmbZndR6w/VGuXWEAUSbVDr2+rkCW6oXrf9
BilyoCjmnnuipe/I5LE6n0DfACqiTbPbGpBeQoY7DCvE3foVfFQe+zqcNA3RKvzW/zemODBUr0q9
GWrFKeCWu6tKtwMPu9y27owjzKvMS2sPlBfQv8E9zujEt5z9hYz1S8biZIGn2rGsjSl3Z8umHjln
BqPR2Z/VBjlKtnTf6YurgySjgeW73bSpVS8EAfJlR4FxT4v8zbknkOpStNdW0XwXhmKo7y5Mgm98
Z7/979VUZYMBovbS7adSs1vQvIYck/nw9SWobzpP9IRYi5CRsNRhVgOMAStTct846sjiOcwiJvhe
dYEpbhwMN53N8i+LDOpoobGKbYosAX5Rsf8/0zNX4ZA2kE51vEZtwQQw6JjiKVJs6kftSqMImFzJ
TnOO1aSWNEc2MsKZVTOxTCf1VswEgS9n+rT+Z7OG7M3QhfYlIt1yMZpwPIs8KpWOlqIiRBRCbvGm
a25sTQlMdbe/TNddl6kxBS8nYDfZi+K+WLE80fykIZizZORbSi4dfcEgq+kTQFbmPZLs65TZ57ZK
oqGnuBIzP732MemIdi8THxq6Bh/1+0yE2zO0x7IRh42IPhJhKFI0z1z6cF/OdlzOO+dlkJ9EQjaP
gdR5/vCrcmJGDT+e5snIS0rxYlxNHk/gA/aJC+NEczcmaOT1vy7odEu/OstaoLmmV5ee0H+iqM7S
6bq8PCcfab9Ill/VZxqEQXyux5QTzcBMfF/cMDuAZO5d7vjW9INAGGR/bIYvl4FBVVbhP7wBCHiK
8qBKO7aSjpxOHg3QON8+Bjny+r/kZhlKWh3XFgKWPA0NSOyLAE8Ge45NuKcaKASKMjkR/XFlLVhl
Ue3G/roJgq6ydXECzTi6U+0bXpFYQIaMNExgWHl2rhfYM4GzdRPif8RDascq86/K9Iq2oYYuTG4j
SEVu2VQvSyCtmrD71p+Ew2tJbdTY33Bcm1sQaEj0WJiJD2Fm2/h1hSfUTxfkBqn6repvP3MNuyyF
dRJu0BZRCT7RiQq9sM2jd4VYHRUhHAHYinORYIUlH192yLZIP9AEZs6MENs7mbahRuFwXXd0tgsX
ThrHSaJqtUUVf6Ukhfa66RbONACTRnQ9yAvY9x3Wnm6tWzg8fCX2B9/NKHjUWYknxVTTSU80DLi6
42L75ptk0SeyS2UszVDKP90ZP8h2XnCsEiZrIg13hgz6PuMUkEiriZLUJFOTi/Mxa5yPzmzlIb0Q
B15W1a1Zw8MvLVc3WuybisMBxEkahK4HIEw5ornGT/IAYQPfDCuFomNymgXzvEiJ/ddey3LXTASv
8SfzEnDP2skRdjpiwSUC4dBYdOHJ6moF2Xcf7MsYQOn4n7kJTVM9a94+M/1TBF8SMTBTdoFxplXf
s1WMrJK3VoQiisncU2zNruJiC8p92X/cUwcohAyk6RXnEktXFUPFrxVa7hGb74JONxpZ6cnvcl+X
AWbQ2HwZDpdfLqSLBD8s96NRbdlR7kOMwJJSgM+Xrgv+1/9F2F215yP6gA87S8KEDmlIByaEzc8X
Yq0bzbRf6wahRRuWv3m6fOgUYgcIKeE3vlwFAeslYxjm8/j7M/uFbp/7YsYOQWkfUddx8stz16ko
2pHCGw3HNvl6RpobV+HZhhPSFlABvYNVfouDdsSL+qq36WI8ZcW0FIX518s+imdRDdY331qEjIrE
eP+j6qNkCBrGNuFhWjuCk8d0OTCzN0O8y2Ja5HDABJ2re4yBvF96WPplRsTd6M6ZRg/yhm+mt1o5
/0/ZjTbo/BLpNcvV/HVYFGFEzuQVN9jZg90fHe6QyZ46CnUFcsxP25bpxyxfBBllUdeOW7YkQVE6
TLVb2CaSRuqso7m2NgYj6v6rgoGcMYScVrVg20/wxEuXZV5nlO5ghgD2L0d6xxaVwVQj7/y8ZESD
ax7rwKtA1Y9pHB/es4WLzF6Q0BRWrsSHEDhevgEdywUWtGy//P2aHaavFm3ddfhYHHGQjnmKf+OQ
9y9V/41WsgWA05mW7o0bgmkd4cYPUf0OXHXgzpRVVWldeapm5rP6YvVpYVMKIZGE+8i+aq/6KPq8
Si+EAfleMeOpgLTHMuy1Tyd9NVdlJmj6KtlurpBu3tzB71yEFAGgRk283suEz9YL+1vwSkawcJTt
TV3OvBAVpY1nutI71DmdiAYR0VpRbxn2tfGIHINx/eL7p19XJo/8JhxB5S2fdRZEtsOagy17H7nE
z3S8CiLN1tse/PNyNEooH2ENRNuCdxEWORKqZ/+v7GPsin50GjVRSbm/PZIMjV3VNdaZ0sg0mIk4
JsIYQ3SU8h12Uzka9n6KB6ESkaPqDzfLh+Dewm/d7lGeVVS3IYQoxOzRA52DcExTjQ0VG5BMgQNb
K7s5RD8NYYT93wc+WjsGWLeKfYpDhCAqSMjLSb7p1kBYtxrAsuUsH+0LjDh0x+m/j4M2UR0lfh9T
5w43Nznxe5davSSvhbVYrcRlIORPSrvVfr1OBdZBFbO8VMqgCbi6+XX9tHQWEMjFNsM35xY667xf
TJJwg3geTVJAcTKoHV3uvOBL5ZzvjlT7U/wJVoYGTBK+9EaTt/96qIZmYLgy36JyO2hdYe3DynQZ
J/erLrKLKU9pyRpNJoAEOw9wAzRXEr4SxpBJbUNslwirkjmgujJjDY1U6LCcA/pbUZ/YDmbgnwFL
PmRVpyBFOWrj4/9n+M9MD83BUl+YoQc6OWv+3h+G4NsCF/Zd1dt4ixMPCbJYr+TCKZlLdBQ/Wj0O
csX5MNJ70kqK12kAyKQQsaYpcqeaen2y/F2byFwMDcpB43tPjhiOgClbuz1HKY8/IL/pgox2twA+
WfGg8rCUom2KH9TgblpmUyQegSLTPmrKvHFHhE4HLOCbILkdtBRkSiRcSxLQ6FGYwWRmyKU9DNzv
cmz/dEKEpDBDMiLy8xeByUf4LLCDXlTcb7EdWZBHCihFtL3YL061jI/dmUu2TUCYXmNiUJLB+dZ9
CgWYRBt3G6n08NCNoLaBAi/mfpHVdqs0OPwkLjJxQdshGA9VT6BCc5PXP8ucB5imChBpxdXITFE1
xC0FqVrJR8t3/gEJXwQZWmHHtNcEtp6bwfkgl1M9hW9ENTvwk6yhnN7TSedn/ttdAJaeZvgK0LAn
Z8vBF9DvAY7CgM0F9Hm7t+J8s0IYSpkS5dus1KnBVA8sLlZOWVdsind+yLng+P3rRRAQxE6hs4bb
m2N46luh3NyQMuhOf8owBgCUOwEyMQ3xLUlR8TlZr/d9yHsfD1n6LAgZbLEkP2kOa2UZ3OZ1Q7Qs
2JTO0Lq+LKpzbMg+rZr2d5JHvBqAorLUKL1KbPFrbxAigbOUshs3K3fhe5dRp/YbDA1adWRXIPk6
n35EcLphUgwOWocuoWnRhL0fBp0BE80Tdsltnx2r4vHJk087F38fVbcYagJIRRQSiJ5DUSv3IAoq
1JnZ9SRTi31+hxLu7CJzUOzyRQeXVohxJs9NL7Ub9NjvCldNDKD8vhKGfIYMzjd5jI21Vd08BVQj
eACEysE/ugJtnK4QxZwn799exWUm3uCQ1LwCg5jZ56gfgTEBbmdakDUmdEmmLp921HXuIH2QZ1fo
VbAkr7V968K0j7M/UCDeoC+BToOPnTfJDVeOsmHqe4kbAE9IJ8OAaKfI3o+DhpbYnS/Ms4kglwlA
8YwBrjNvPY0b7SAlmymbvDmXOrrcysiaJoR0wSa0+0S9JwTRAgdSxmEDM/wC4rkiywJcEMGwvlg4
zvRimpGnLtHGbOacQ/XAwZa5rrvuE+RrUvW1zN3tKBk2F3BqjUv3rK7n1spO42JoqwRntZf98jCV
K097/1LhJJQYFn3UpuOaCYvvv8u9441q61w0jdMxUWZOPax5MGXcAF1e/ktHNI2lEwBM9Ei3SzEF
hLt9b54t7XNzaVFB1AjMfLo8+wzAkMQtrjdid+Mg7ynKqP6UephCK7axjiUQbbqcARMwxzH1vv+i
sWMhY5sY64OtWGUmR0CE9A4gKep6a4JUniUxWPWIO7m3t8BPD2FJCbGwUErlawgu4G4cq9zHHtdl
dCPZ2WzUSCHKlVp+eufrDrT/X2ib2V6Awb1VHp5aYDxaqke5jJavu4aufgnuXy7lGoe4rTQ9O+w4
tOePqZfpLaTz12HUSeHlAuImlq7KQjqLNerZxCwBiPSXm237z7QG0TQpPtRvDI1sCfmcsn2HApJU
XN8F3K3GvCn73dPGK23y3lDZpoqYdPcRblBrjCMEV7YyKytE7V21JjShFi2+5WmOUra3mn7v2DxM
vF2pSS6O8ovbfv8cmP01jKJUjYxyhkcnzu6pALVgyhIJqoz9nzVdM1xvwSjNZexgl9Olw73HLKUY
Y2dUDr7DH03T/pPLEIXyocR7AcTbrwFmhZFN5uH0E7Ct8O0+BiHMY1pnQz8oFGXkzXZoMi2SvR8B
cle7sX/m3AwoMEGFxNrujco7JHcdOur2a0Byw+wZu5h4fnAsbFfCIOpsnfZu/xFs4Zy5XkA0iG5a
bS/H3oon1PNNcAJ/wY/vFRM+F0UneQcZoEML9GOFBdMnpUewgKn+EVqnqvUaXfAt+wZXQolWvnqc
7uY7OSDu1GihO/TLCGNCDtRMd0ldZqx0q/4CDEHObdLfg1We8xAeARquH7inIrsYy9jnRdfT9uYw
JujbR7SS579zSSfuMRWCEOT64kJme4RzmzbYs+wWW/ExmAHjik3WELrW7WZ3Gmi9H4/YIvw2DcRh
VUkVNWuFCihjTaP3YySK16IanVJBOiQAlpXceCCoCyxghIuTccInA9FDvlvnLq0LZK1oxd3AfdKb
2nQsEvO4q0nnKOCX7Rz6W9FOMM+LJd4kWtV6PmXaVHwobP4P0jTXxlMFSA7sCNfvihoQO88K0ZTL
s7325vUOTT4E0UxYcrVvIlc9Zo/PmTZlYzY7JdFzpTVm0KMejUyq5bB2G5wz073OuoieFdn2BL05
1wJDwOJl/qtkdwRDGxCYfwsaTxvRCPXTc4c5zwur6C6rdsQNsnmYqjshZxSey1UymHnHOYm/BgS8
I67IL6iVM1s3s5EWkNXxCB80HEjHD0e6sAkgIesQhGNQ2lVqI38AGsdBtaJkiMJqjaYRiEXuwwgd
AJ49T7PsM4ZgCO6PicdbzPCo3Dnb6oj7wpH5SSnMHCIOKl6Gscefc7vZf8nTVRiN0KFBAuoCaoNB
dCvMn4RxNilOqEoCHg4C9INLImfbUSiWmvt7awLCluiFt969ogvklQmCnM2FgIO6YcLAEObAUBEv
wu0GCKFtq6k3fPpEIeuTKoHpGtD5bZkBvnqV3phlXO+EabskvM9kPEJqFN2NPFYOC0Vh/DP2mZdt
hTm2+9gC/jmjgkfbSQPQknakbZBb2CUmG5wcXHqV4qlI0+YgmmR+w41T1KYyjRcSoEJSnFeVbRjw
vENENHK7jeAAcXFJ9iSpHOHxpWwJ68Eq9n5npwYe+Bd5NE4k4m8+wH7g9sMHPa2JFvGyx+Z0mXxZ
lzWAsCNcKFV4h96rCwuV/6FQr+dMbMJxBtL7g4RoTIqNG3C4YlgFNUjEeEpi4GfBIP+l3RAz/C0+
TY1ImYWF91VnfgIb6z5KUd0lnrrHSc3eY8xMSWcOAhzFJwB47OfRkvjkhuxyHB+a9V6ixeWkp965
IqGrkEjtrlCn4TKgL3bQqwVXuIGGs4fnuI6Be8QFLgoMyt11oZ98JrZWBTdcEpPzRxSxK6I4CrZc
2ERmuDT+/Z2TKkfTZOQglqNsWXltKBFFnh+3b1+Bj4IL2iINFIV3psN0l3hNknND1kliOj4HO3tB
bmLXylqOkwQ05aAz+AShe1P3PBHigSCd1E+b4+NByIDjSR2TIEb8V/oemlLoBkbPoOENinAwqaM+
kekjXTrAT6IzaWrWKfH44/6m9duASxsIgDRR0F2SKel4em1+9cGIz7lptq/wBJV0obWrtz8zHlLC
F2XCDEBOxE2DpxU57Ga1D7BMZSF/FyBkecnuw3WJ9/SwK/qFn5CVNCIcRGKCb9pDxSoD3/vH08CI
l40P4YjWaxJtR94jmlVvsKTpJmlOhfBs2VWgigAKG18fgjPxFxEJzKnJqTe/zYl2YNRmjx5mhz7/
eJS4qgEetO8bYQ/c6rrBVG98n1dN+UbRmHGCM4D54YZ0o866Z7+1jFGKPN0b9assqVMMCqLOyR2A
DmRCHrn9QJwvNROj4OamStwiOOXCtONZF42Oea0zMjNrl2NpsIry2jFez4b8pN3Shubx4kipGycp
KYd7e6amI7jDqRTg3Uq0xsmXW65iQrVgSaWY8Pdyukg2P2eU7+m1CekDItFflGcxs2YT1+dpzxY5
QhbKm8bx2REyFB8hmbtNt66BDfqelTC3Y9jYVeXPx/iungB8xo/+7MUC0qmNYmdo0UJuH6A95z5a
jPnjqgBCIzjXWc1BPtJ8R+SeCpkUVZKBiXo3COFIFY0OZ9mfO1tGiSrzKulVGJKj0QIQvvYmK8yF
bu8eOq4MA97WpgH/4SNSeWrhXn9ElwZl25MtB+DzfR9n1d9520bFDSelP9zDr4wrsZPrNthj44zy
TTAf8b8UXb1q3dn9Mji3eF7LYFSYdNEfmRte7Rujk7F34vWaI1DX5sKTMXghR0AA7HxNeAYvnlap
RkSkluH7SozL253400zJ0oO6ZQgYUmgzzxaUsW/A9wn08xkxB5Ppi+H66APOpmygWRuF7+k2+a8j
fZWTa4in3JMc4b1ufTBVAsEvNdu+BlCoo2FQQNjpp4U9zuVWmGmbJuq+EZdfFU5wcNuULxF69p2d
FWUJeDaohDyCNtLaq0jfvl4hSotK6p/Hf7jmmtb/20Q3ccTdH0ynhOrBpF8n/6/oIalwF+Ik9wYc
OJWBol5JCUgS0KY8J9+J8wamCOTPhYtpl4bWXoIi3OHTaW001YLufqXwFpwBXviroHx1+CBX6aYE
A3Oph1pXyC0N1z61MvW8szY3G84nT+GpGE2vvsJ5sTDxZZB4RiQZRdB8imqD0m/gsKzGvD1bF12J
vE48mkyG/k1lSNHOyNpZao3VswFpHDPKEkfPbfQP5+rAY9Tk4mpZ6YxRnl09vmCmkykpw1cylhnz
uxtxdforbPPSIeEimIPgEW1b77D7Ye6rWEvC98dymigexJf3wPmxlzl/MTg+PNvGwNhe4AOI2pE2
50m/GC60ik95gCuWLrOgA1S7T2ZekqslA93di5DJw+A43niK/SEiw9Eh9MkxGTKHWfkzy1yJrH6w
yacMNc5jQrMWrgsBo/JneoDJm3zkHJYG5gEoCdSiEpfOEpPQ3ymRZ8hIklyWbHVL5NkZPtqLQDm1
VrUEWNFjtMBrLJEijppKn4X0oI4e1DxCB7B6Z7JIkzMAZopbkzE+QEQf4ZNHQqqBwdRFLohf2tM/
dhJFbCT/PzulBXIEHMwy6mSOnwHRpwEl8jgZoGf6QCvBshTgnOUYNELlaf3YIhbt31z4xORGDwBz
fby6eG8OZeAdlDyRvRPh9IvpYItNiuWwd4DVllUbKFSpLUTFJ0aMTqsLvJqG3uhOLEFHOLyiYKgf
bmI/Zug51Dcw3Y+kCeF9ISnCChWMwdCQCqctV2aXk3z98W7ED2xXMNbE9ad2minN9ixPt6r4DJSc
2IlpvF1eTfV+Los74pxdYnV0zQC3UbMZjEulojRM7HhoTyX8wDGDCFCNqVrIhZnV76uz8nBllJWe
MPKwgLAEz5giQAyZA5nmWRbO+mZzV4E0XL9D6i0KwlkjpFgrptqYfyveU5cMa9ozWO8w7kmSLrtn
tB3tKyovk+uGCxSdSOX7WKxLtVvdIWxCAshOe8uN4Rp0e7LPgQuBujwv3p+1XhhGRLuIvIHgS7Kw
HrT4BgjPbNWaUYolWqJ3RgoltKAXobtnj7liHe6BgRRiVtXP2ldpyW/kpn1u69MVnKtQsmvdWvze
GTdJjGgYZp54wz0dCNzXRxnMAoPBjShsJ0z13nEpmzIyp/o+/Hqrd664MdYaqs1HgHziO3IcTzrb
o9MzRpOEzF1IXIKHOuS3hg1KdDOdDCx9ESc7zGAownJQAARJJT1h0RStfs8U5Nqh/Mh/5CV3XzDc
J7RvgmhJWH+EKuGMlJWgtLj0463fsrk5oVW5L8735rhqvul5/eJSABVPnocqJrPcQ8yc18REXaut
kNyzjUtQ5yX+C+521L7LI/WqpPj84wstVqtpPZOgIoToloZCYa0Ko0a7kWviy984fNkxn1LU5ZwN
sbzFT7j4mkghFaRItwmJ4GAkIGKt++gutMJ/VM1l5gVzW9rwbfz5Fm/p8l4T8ssBU9+ot9I+W1U7
H6Fw7PS7fujKY8aS+MkB7fqWrmxhWK6vYgN5jJOH9jZILj1oa3JfyswjR+CtMyeF8C3tYjXNXKCg
zPXHScRk+oHFN511gYHjrH7d8wNUEPp4rgKwAwsOCwRRozN2ZIH5APW1K/VDTGGgVVVE2m5VwQLU
CDDO+jL4jqNVOVuL3ng+YXfSrwVxFuCXXPiHQEeJ/OrSumEfDkrn1lUZ/tiIvLP6O+WAUYLwP5mq
uuZMDEGnjT8iuuYZ8kYqKPauUBodcAARGOWZ2yyhqPdCotoMeV0POip3NixwQqtcTNwF1J9XTHbm
zC+Vpa5BlM81IWgPUxb2BW703sccd8VovDXXHAfeVFbs8Y6LDPPBwHcevkrXUDeUEmQtZ6TbVFYM
Yq34dxORtqlYMJ1KgmNg5EuejBeF2GOtjnqELmlhFyDZkrXEf1MbbSKW45kP6ThPaBicWSfjiOjI
9cp/VA8Sy7KRI+WKToOGRVnLlMC7rGTUCb60TZZbkhBIgqEMKGXrkegKsrW1gsuZQXBFG1HEQq0U
+U/XookzW4i28rxNnUBvOevh9zUOqhoLNeSSTeY4aicYUXq20M1JfBSBu38plXjRObl3Zg3lxRvv
8sGzi7i8C3GU2GekPkNEr6z8D0Il/Os91eFGr4HWVFQjy5XtgAO9k0fejDXWBzn6UWXA358Wj8WE
yAGOGmf9NX4DDlmFvCQk3PU7y0XlsOYlTRv5XfinguzTJD+oP+TXQD5An7shcmQ0Ris5/HV+Y+Qb
aKEQznmhQcoOx/sjTLk6CodhxYwdDhVPjOMcuCG8fLoPzhGchbJYgUeanLEQHo5CbBsCREW5XV94
H4kDG9NLLWVf7CI4XR0zh8I2piU0tqiaFsHPTE6YzEi849ySUM5P5LhVFOnsABIntPJZG4LyZwL3
QA5DAeevrYO0u3ML5qLrQYWi6ceM5iIqCOzvLYi3yPDCXAIA2Ldy/8QhU0LLYfjCRofih1vvyCvf
vF/Ml+SdSgRhGYF4DWlNKaW28LPIshdKNTVINZoVR/elzaqZtlyF3D9DSpEhxvejachrNU0OVdjk
Onpil+ppaoWjdZDpji3S1MFqCzn3AyylyVUyrMI9yUtB5HyR6yM16PvbJx3/xNfHewiY1vvfesPr
80sq5Mr5BP4dDOCLzreF7lNvuZnlh4u/6VgG6pl1p+8ZM5PmMp+bhTnkwvRd2any3bXceDYRRwCa
a1UsP68BEuu57yIdCMHskvbhIjCWPWPJbne2v+PtljTQzGGUZj8BW3xRGuAkkShEbCP5WuLrH195
6TjxiYhY5B/qgsX4zvr3kNGY8ztSMWy5/Tu/hc9TMMSo7MLAlgn4c8Lz/IvdWbXdSelh+jm2/Hwa
xj3o/D0rIkZkZFDM3M5HwwkLhmrq/e64Ppy5eOhFl/qaCQwDUlkjFh35KeQRd3nrgDsjNXsJygVX
b5lkfCu+eXcxqTWDuBONM9RgojXbglBIVnYNY7IgZA32o3/2p2P70E0xbOBI+sAVLRFmeDF5CAYD
sSh2RY1e6brv5Z3bDQ3T7YgYkKxLuzNvA36IOVIPpVR7kq1reTDTRBmcSD8O61ivSnzQezkCebdU
opPwcqQQbTqQsjSUEfJ0BRyHsVhVg5w11f5lbio7u8Fd7o19/+ysw7zu/W+7dU+3UCCNggIMe6I6
lH6/vJQklNV9HcMW7oxX1S0Wori1HOMQfcRCtXYXQ6e6bN+p1pjf0YCC8rGpjhG38NjW6QzOiaGH
ThJL3Sr+TiTg68NKMgH4tuLe4zeic2L3tRecs+I1BaXW3Mjk9MhHG4NEmvCFBtKS4Rvgbm4aUvG3
O5t2xh00WwYbXLBUMFosmhCNMU9pFuNqdgTilc6861aVrqUljNpREyRni0KkhoMvP7f+Pxdfe1yb
ZiQznxWnXr7FPKHYaPMKgkB4cD8hxaYsLdcr1feFhkALxu19//ObOt1RQE9BGICNchLFNWqEBjbq
8ZmTg1EGHhtCY8FbFlZnjMWeX0xXBCsWS2f7IEllgvh0nP0e8Fl8akUQu8J/bDAB9K/QL1vVlULt
F1grWmyLfsUJbwsc5CMuc+xi+H6S15hwUb6UzUK4VKq/0vchDQNkv8VTSjLEe6otBd9VI0VLbgG+
61VEUYzzqQc9R5w+7jOtLCLTvI9vXeQqu1vTOvo8YODiC7hSleDHdWsClNhmozxpWWnDR+u7qIaW
REI0Apq7cg8HsK2A0LQ5QkhlRkq9Og/3vCH6PEezDg/DYFW0Yle6aohdMQpqIs3GcZnY0aIS3puP
vQ0Gmvr9hMkeWaiY5/GpKx5kAGw5d98lywJ9t2hECzacSWdzWE/lVjJg57Ly23uMhTvApz7vcmxU
Gg5UYOFK5DwD6c6+r3/VsRQ0ThStK7Ra27XC2YQp31I86SlObP91Kr5sAtltxjlQGhVjHN4EpAbM
MWROQjYolQiTNaB3oUhRmL/z/XQruAQBlZAHvdy2dpwylsSGsgA8cdI33tqqrjt00BENBK5UbhY6
8HLV7MBVagmWeiC9Ky0twFw/W/2xAA2729oscXn+2M9spY8DDwK51MpeRyKsU5oo1y0e/IuHoso6
NlpuM/WvOAM2shaoFBlOJV12jMOIAvgmE+RDeoeSYKrdY4iA4dUPagmwzUykXeHxvXeijmrJUBiK
DTnHpVf8VdbNsu4zbREtM2D1ZbPrw1wAUNNJdx7xhzjRLwHH9XC8FhIS0wRZ8SuWRk1NR+xlPTKE
XHVF71CZZzYYtYYqmIsdQKsq/9Xak78azBlcdD3LK2VG7xLDzZlYH5pE0oBmm7qnd6eTCD4Z1MpA
UBbR1IbvmTDQHbPWXUM5i5Qz+tFyQ6o63+BmL1No5Iyioe59WOVOq3cnLxLxT5TT1SQSmnbNSWwZ
xDUu39Qvda4+Ic0mr0rzB9LW+AsHEgO++nYa6VDxicmioLZ1YWLOTKPYjC99vnOiNEc+kMyOP3Tc
np+QEQlo1eoFCnwWduoQXw+ckto9O3UzkxyfcOTTF0TmUNvIbyFfkcExQKKMURcGUP57dgNp6dcC
28XNsvA83pN4xF1O8ns3coF9I9QOWnWlMVKIQifmxNyKUNsii7+XPH9r1Jnmp3Na4Pj7S1wtsIf4
QGpmfqzvXGS0nXROjsvnoSUjhr/c1CYFrDNvUGOzkh3wvhRtQqJXufbNv6vBwLtmlLdFW67155QY
ngZFqRZjbqb1AawKZQo99cnYdlPb2y8cEAGL9P2X7ynE4qDc/WYyC0OpfGZnFkVlOEa9m2vxB/hs
SrXv/Bvx++ditz32gWFA0H3wz50zRLzUx8UMrSgSN+TFpIs8z11DMyaPPPCfUk05iUKqtixj0U1m
ItJH70BgIGShtXrE4xLJvkbgDiDrydrBOfD1Zlvgke2ZawWIMK1I2xdVPbh4vzNnmuScJMEdizZh
T+I1TWUCUk9tpBOXTQDRsw27uOPRGVBsoqFGOuu6uGT6MZt6yyIlAfv1HVRWaSkFYLqyBDTTc0nR
dURS15T8Itcw5x+M/SVhLSutWgqO126BNkxsrdbRj42cWQ3fJg64I7XKN3C0pRtbg3F53YDFDCI9
ASP3vlPPeX8sA8V4zOFHJGqltRIwNu6u8SUel8u+XlQQfh1Y5urKbUOCGb92kTWMO/6Ehnax14V4
Lit/5w0MwdzQOsjyyybDoh7uhvfWtYCRZRobgnb9JZiQVEWzCQKTnNKd3bRwEpdmXuqHkk4qm3GZ
ZZinYxGkExGje2eqP0KoAod4QlC1R+zp1y9kuYz65KpUOaygjM2lNuvWnik5+5TCOgkWt4POBfc2
LfTLmhi0RU4nIS8VVOEI5BPm1xV/w447ztU3MgTPbEdZ5WKvel1UJHB6fg266rYgBsOYwSvR6bWX
2Dt8GinVt8qZHsMhCZTTgFi/FfJtJA+LuKkeEeQFGO2iaHPLe/bMw5Mt4Sr7rCoVBm8ed5ENLBAh
MEO0RP9Zm7FwcGRLlpd9CJ5XOUmQLNs6GwPdtEmw1oo7/r9vSa5MpXScsXJ/WxARyo3D3XyuVT/D
OhkJTcaSRHsAC239ClsTJawNAczTtR0JRSXPcf1prW+z8Uo/daHhG/AlmUStkH/5rDYKma7cFltg
UJdySipjrEVTZ107bgz5EzsPCkHACjGbZfT+BrDU60hkcvAiY2w0lCy4U03UYld5xUMJqyj3aZod
fpa3qcZNEg64G+65FB/c7oWrDO2TYE4ahrep+X5YvMT/QAXkUZBDHWMyLQRudxjYay8p5TEiOeD0
r9ulgdLG0Ii7cdoK8oTzAxcLJFenxiZns2B51VN9Ks86AnIDfDXKGhERsyo7Vbs0yQUNrreakHN4
WsxAQN1YOAVnxyWhGfpxujZKSlpQxC5qxVHAN+TuZVanofaGiY7JnEQcjMpXbs9BwISrJwBDDfV+
jVSJKDqaho5uPEVt3ziDY8MreWH6RNy+2F8fet1kG1dpNooaN9mhOCkWYN9eGWLWJlPlN9LhKT9G
F0vQ3FKAPf98wv9Zf4684IpIqGzuv2WJRPeOXdM0grXSkbsLP0aRIXkd9f/gltlFDl84wzKxbZjp
raSRaPiKiDeHZ9ryVmzOGf59eEt5bMexxBSV0VT4AwaPOsEb5AzBp6L54u1iGyEQ/43LTn1fqmGR
f6xAnthnyXNLV2yOrtYGApy5e8LZXdwWsH8G/1Mqk4sr9vfynUC1P69LrMWvCdrBlM39fwOhlJAo
XlpjeDNQkdrhNS3jC5lEvxAqr3eK5vJymSD35hHxxau4TI5P8KDhkEaWc6AeZ+QtpLCTrjYq0S5V
9EDOkt6cEu1xf6iXrzY8QoZ4cSS1oSFSrpl1qTsziXgnct628kqemuV87DZRq1Q3yv3NCUyHmqmT
hk9uGptCdyLGIwRL+i45I+tz3j+wR80K8frOnpDiaelt2zYd3NrMYmjp0iUT4eJE3UfvCopGVMG8
esJ8MqmDc3gS3pJAukQrZQxEGAkToKIhDfzfqLDnjZTluMnQPbnwP3N8myIi0CqNIcjrEOlYIEJs
PLoxRkm9gfG5mw6fgfdo+szjQGkpxMRRFsAVDfGmcB+5nGNUKN4D1OM0DD4WG/NkqLkvrAsdRRL7
mD99IcFg56zWy1LweUaFidhthTTCxLl/uwKHQXIEOsfzI8fU3VeUYgi93fcvvcQhdSJb59ncnAjL
jKkv1hZmmU4T/lIs9eHgOHpha2PlXcEsA1dEtCtuiCdUnxlpLGisU7EhwavjuwyuuXbFYwKXeZIe
lDlold2D0KNejbF/LQ2HvY4Et+VoFaQdxbqrWqCgjcCUIGKPt/wPHa3c5RoncwTjXnmdmt/8bC/Z
ChSKSFSsrEmoDAcuSkGtPoOSSajBGyqXIYFxrXlydz6O2VIu/CK9qoEZ+aRNX6Y5/RJkeo0Hu1E4
s+fQpW9s6oDrHZlxX9HTG0HRfaVxaHbwrMk0Jvxl27CD6U+/UlLKe1MKxFh47GeizhgnlfzVqCzy
pXKQHcE/HmVfQfsnWe/EMANheBlTnCH/pHI5bQmqGcxLYKi7iVmIdhH6/PQc6e2+0+ctHsk45oEO
AeKZD7mzzKJSEEkmR4+35nVF1TTyjO6kwx9kb9VhI9H4KHhexfSzhkgy9vZRkzD26pJFG9fuK/Am
uCSpQQ5GmgP5mgqRbYfeonkGHngE43u2Hb8tX7K4+hXqqOTHjDP8bi+Nb23VrN57BMxDyR5UjLiu
ZCeG+tDkdog8FZk/OUAyldwCyYjmworX15jUdbWP/NdB+wCArbjCT8FB33htHWfqIWRTsswP3Nc1
qthsVWds8ItGiMNKv5yIp66Vl4XDiHxJRV/bkC0xpgE+RwGr1MBaoLycIhgKIkV67gdddsAiohk6
OIwaVdTy1gLXMDifZCHPMrxIWW8WUFBM8BkO3S1hGPFHpp0Dz7ygJ34LQ9zfhLo0tmp/vEtpAEAy
MFVVohRn8P0+gI0XxGMa70ii8kHjGfFmupnKwaa0xB8rEdGwGiLXe0m7LKSENGMUstr1ELEs4XoA
QhObPXeDu2c51VWcrBm6KWk/XR52IyXTtVpO+1mpspYR6ydcFFPPIOZYgSKHE22ZAMUjYXkMxp7+
955XczU4Kpmqgsk6pFJPbuBixdWkIjXUSFBwvMRk6Oa/nemqayHM7bfYCxBbRshUj/5zrGCqApFo
hUCND4Y6WBhGuvZ0jzbzXYqP9+LtKlHxYF77dxFrPZTcOyRGlWPERIbmOhBqPkdloiaHEWhF+BhF
XBXhh0yoiD67RwdTTpFCZDx/hGSBI4EnZ9a1JI944P2OLAcAu/rdeO4Z4sXhNsYQCGbh144FctcS
reCzXB4XkSNypNA2D6w+4ttiFw/EO1J7HS9TyYLsyoZuNOzc/g3JG8w2+bSx4RoOum0kvIo2TbQ4
dZPPEQB2BQ+nRuOQbnLzErOBMFmtAru/v7s4O0s0mBu6PTaxYgLU+RNzRB5WSeqwObnvBCUtOGdM
ll9sXE9PjpS/ys+paOk6NAPg6o4XKFWXDYCTZks/m+K+1VJ/OX/vixQC4WQHVv4FHAVc9HBdWljm
j4hIqwCuZ1ZOjexJEIB2+R3EtRkFYSm7FwrPWiL5OvSvnGu/3GFoteeiKhuACVbQ+5EFY2RBOPic
cdSccjqfBRNoLSgbD5Usmk3+4nz/X/W3KPDZ62DvySbdvP5+kkeyhzthH2D4hpRyuzLsmK+9r8cl
LcYsN6trAJ/29uQr2o3U3PeRGH9YHmgGn0Dd0WwexPmDHR+xud2IJN3eNyvxFjkuaFWudAGm4iVB
bIKnuQi979x0aJHwRrrcbxVcojfAA/zjeOUqrwnkQO8hwQWc67wxZEU6/4eY77/EEqPTLalZ5LzS
AXlEL2Vw6WjVGG8x2Vpt+SRn91V70e5UzJ/Wnf1j4aOK6hgz9aoGMqfKAYvMBB543eXrROjVo5Bq
hDL/9Pex70xqHAS073Eg3rXH7Xc0ahTannkpLHJXmCq7qnsOnTbgKDE8Ms58+5yyvLJty4vN6jGM
b56lvfRrQXHex+z0lpaXukLspWoaA0xDJfKMV1LHDU0hkXIaHJMi3ovfZgsOgEga3gYsUDGTfEqZ
SlskK2EtEuqXC17NsSaksu5k+3ChLxlRduIVcZQC9OotdIICG/M0XJMO6Jda0B7w7G1L08qkv4um
U0KRrA76s5yf4hY9QNfwDkSr/BW2RqVXIt6vij5yb7KiRPWVctPPFZPctQsxMFrY/ZlTPzEHDB3i
LYe7paf2LRTrHYwTaop66viymBcvO4QeDovNk1k5YSNj4mn7A7Nbe1r+r5G7lIALwx09OBu2krAT
urmy8VY4838vKosiK/tTHxUFwialxwY2/diU6HNqHEvVFvTS5aIKdUJCh17yZ9+bY1ugrHFsaLrC
OIU2hpHnylAzOf28uRFxFFBvtFfW2D2rFcxZXwvgPQQvnYAADn3Tt8PbLZ1QeP1Xh0YKwd/95EGS
abXVN8zTbu8H7daPwAZtGxrRusa/LufYyXJFFanbJHMtR6iFn2GeCSalpo8WR34rSfxPI7NifvoB
O7+gmPWPMjkDs//bRUiXKlMN/ibjTDLKV4jikoFqGBKItzTJZGfYnmjdv0D62mjVOmWhAE6oVTrs
ljL4A0u5U8c46UNUNl28L5ZQzXcLO16LaZPr+2JVn55+gDAR2i9dq82RO71fPZuxxoDXYVmIvw5G
I46SAZBFZiZY/CE2u6e/+TWQ3SI9PAwZT6t0WOJnD4OPXeDDszWHoAMyJhphWxY9tIEMSWvO5uQH
rCUbtxGgmKmtd72mnHns8AshHYX4aYSz6TEZdD+nW8FvAYVY5+io8JVHjcuFQcISjj1oZRSGw2U8
r5UlkY1fWdtn+9pULARni1mIX2AMqQTz3rwWKaBVFAAD2yH6pDAwQDqNkAWGpBCql1NvMS/JQ122
VYhUpnNGXZ8znyl21wEYWVLaa4J/PTaPq6yiWl3rIK7JmD4jxQQ6i6dJw4J5L01yweb77RG/GDlZ
OzHQ+QBaJSy1Bzd8uuZd/ZlcYgLWQartSpzatOwaC+IDCDkMHRBc5/hf4tmxjZhvozysUMWqlrtj
HspI1jny9rYcRHwQMm51JkSTNk98K0S4jt0AH9Li4jcgtpcKLx6MZMZOdfPcVwrLR2cgGgS0Q3nK
Dpc2H/dNArGIuczJDDJkpXXMi67yAFv1EShiKE4BPmPm/KNSC1RIRzSxZJ7vjkuAHO/5CMiebEWX
iPdclFipkb90iW8efZMErM+KKOpzsx45gW1NS11lTm7qT94xB2M/bmEAZ+O0wuVpMT6zUBztPQzg
A3hP8tON0BIbDHpTP/6i8tVsDxZO/Azv+OSIOCZVLuiAKrl3aPg+ua+7bq1MVcyPEUUSmE5kcijr
zB18pC+cKamhP9/mDXW/ucFp6BKT5WJg76+fcVPh34IhxYYeRQ1wjkdiO3RzvFfcYKRForWGMPQ4
EK4EQMJr96XCL1d0MjcxF73wuTO264I2eRhrwKKrcoRP5mGi+G8RqBMX2qXy2qS2psKfwcTFeTjj
4G6vpyVeQrF6+K5GGe7cjlrwiXo3hlHRJPhJ3bb1V9zcXeA7jAwSvVeVcSHgcaa7WEPMd4lb3x6j
RouierDAI3rUHtzWeB7d5erL4njtqip//ATItjJxB7chftY7IYZ82xPr/2RGa3xIoYcDNzmlnfNl
lKwFiha0Aqk8JWBQ4sJWa9dwAu/veQOH9nbekZZQSIoWm7LsarC6OkfLGr/5/3ADlFSuZhjbn+0l
5wZiX2jz1Wk01K/7T6suDLPqebLSxUJsJKTU5o+badlM9HuDE1Xt8Mj0V2xIVAg74BnGPxPgEBsq
HKfxfVTxLd1EQSC/WYbhtO7KEz5KX9+gNg6LoqI2/oIqP4zU1C5g2cLCxk89D7tkZR1dRjFrwMni
rVf8dMtrslja52YrSDkBvrMaXn49YsN+n51SUZMrHuwEEGpexJ7P8ItVde+mZWGtu/7qbg6fF7Y3
ZGz79qiGruKDIjeYFMNUEJ/9AbEtkvZ7VSIRCBubaiLJyxEqS0mTHLxRYHcew5EAn986E048F6t4
fyvBi6bUd/G0p6wJ7eqB7LUPRmJG2aiU4UwjsDWFB6132MN7BS1KGdwC0CjmpwFpJG08UNzWD84m
g2pmVP+zv5Kg3JCwSM4xoS8NB8I+3iFyuT3uplUpW2UlLNYQVgM5IvUmcOa0qwzHJFhJ/q40xdUG
Vu0nKz8kMP2/UngM9u0xXk5EpxodxnDyPqi3vEcXks76N5hFtx54/gMjqIdHAiegJjAmVuRdA/6T
Ka9M33USP/x3Zx8rnzx+YoN5fDsBg8qcgvz//sHYojcVWEs9cx7DHpBMkKN1pjZoYMdpbcobh7Ed
8g5mg4ApEuEQsNEbtuEvjvWlfThjENR6qiYKvdy+SG57d8FVGbartOR5QjknBZqFE+V7e4Pi6Yfl
lNTzDJfLNcMYniqMd7nY9aB00aS2sNlGSxLdFlBd4XUgYc3ag7S8rgDENQNODAkt57ltJxa+eclz
D0qy1nO3TJJJEdr2lo0y+4fTUwntViljrfv31WKgaHYX3JEPJrpHwIAyNdovSIdlbT30ZZUTEFHH
GNPqT+HLxy2iuU7Ksb3QG63P2GDZeWy2UXcPhxuHKPRMI9IUfujmh5xebriC56ecS9WOTP6SPl02
/4jONeW8vinhoyd4nn1nAQYsVc9QMeVaxirsA8AL+rIYypvq44Msg5AReGwY0OGpKIACP8OMZzyp
1Qj6dui9g2SMxLEFQF2BPxPKsO7DPtQAy7UJPC3ZY88QH1wfJ94jLaMtIJUUm1L7fJA0FxBCH6zs
OASk9GHfQnyiGfvufNgtTSARzumKNQq8yjheWQlraGc7GDOHaIc1CLUQUCaclHhFxsTblKP6Ysmc
Ue8ZK/CmnfC+P64lTJnW0Yyg1KYrlC5TJaNjqhp9mcNQsbxB3OdiEW0QN1Oj9hgH6vNgAemIGmrI
lTC0ra76aKX4SyoaWWZxldanhCb7mZP+2ta7C1J3ebtSl8s2qenRkjtse/LUP70wEMGJTixIQrpA
2P2QNw08k062ulBSOrb6l32GX543z0wl/9YNm6PW3inmO9iBok4b/nZQmdkzAZKA2wVZnIhn/ztp
K6JsHkM3dliAcU4vXv148kX0kCm8SBzEXrD869zPP25OA+kxn0T8W5xIOc5GRl5WDcSoVakYc8m1
Rwg+8EZ8hOO91O50E67e5ofxyeWhVQuPnVVEKkMwJRxBNdZ4FN2lkEMeZ8tU4FJIhvaJEgWazkyT
G1yNw1YJja6jSYUXFm/ozjwrUDbqasK6LxjkrUQs1a/b6vljszGT0R4MAqIH8dFgdmYB+hX+uog2
R2aMHqB3iBCpWPbT8gECAiELc7O24u8rBiCD/6cJcvsk5fH4pKS0MSWf6WwhqSUsmDJbYmVGfmtK
IHvFiSiJIvlPC+uSaGO4khoVmhzIhCN+s51iFU9w7iQgx7eLwRIYLSNQSNpJehgQlpeZqwiaY8R8
9hMhsnyvS2akUCY9QbVddY+IL/Ggey+INNfT+FzxIRYUU9ac+lMwnfcetr74es71zRNslyp/UCnB
r9Ln/F6Vck+RGoRVQpe+FqRCaOqjeFEuPB7R1VEe7MamoehFmHMT9wqJUhKLfmZN5ZgAHu7tRZsm
0jM9yYQwK7DHS7z3Sskin/QMZwTCo9nAHI0eL6egoBgIYzLvokoopGXEVvNjHjFEdmDY9W7AsxJc
HiEb1fJMoEvsB7hy4L4x1kDmwoq/IHNYD0lp4uvwgg5kSuJUdZuWniUUcCkD4KQ25fzqfX7qlsnu
ii4AgZ/SEsdVeymm0N0NGxCQcODSjl8CY1O0MdCp70c+4aCLJEIUeHPQUEOaWavIEZoHHk49duR8
kq8x94rw0pB49/8EGyl3jJrEvnlt122gEfaHAIfUVFRPJ0oAaasHx4O/6mSCLLYFyEicHD42lAxV
ZPQQ+RsEq44Wa0dDB1v2gxbXI/0I27K4cRFbuHXkcYhLC1lbciOgikjVf/UC4G+yr1bCEYypy7Z3
hPFXLDQYiT/MOSnEDpPipAblJcPB5NVX9gQqZWi7QvuTDp4m8TN8DrDJUPqOxeen2Ymg85tWkyTV
/LWN6z4tvU3Pe5vvqOfae/JK7EMuMg/jAkNLkg6ilybtXYtIhCPumPG2CqNvEZ+LyfR4jkLY6DBn
DEcnCfAZV83uBOr3kGjcMHSQ3oCCejOvGzoAd3//AdbPt4a7J0QTyzlaInvXzQs9cbj3/mO+ApCq
FYTwQVwmyMfnlzlYVL20L0xbG2uuFSOjoTeUEibXS/dQ0zW6HClVMGMvn6VM06o9I0Ho3L8LSw+n
pHDPo/pzMC4xiBGKNHlT8ScTez+YyB+4i37B8roTbgx5I3Jo0pHbmn3KvsanRxeuM6fAaY+HNl1g
JG01GcU0cj5On8Ld43WY4zeru0nDjLPqwTu1gje5q3k64b7H/fUJ1lMI7HjWfNo7mLSRHKu3LnYD
w6Sw8GEeESsu59Vz7WnYmtZy+cd+OBNnfktOFGD/EOiv/GgqLzXPvxpa3R47qhXYK6FRjFFZX7df
I820yNOikSxO3BUXkLPs53WS1zKLvjQeq8HiaR4CCNV8lubfg2Nu5EUbHLYlmMDNGaKWFCSQ3AgQ
sVAFTEwnccwpXfAPNKU87Pd+Ifzrj+tcC1LyahQuxIeZRrrtjfI4s1NZ0MoyK3HQT6lDvThYLEg1
haHQi8/p7iGdiq/E0kz6StNSV9QK2cV6X7mgnLk23/7GaLscBDZWya7Hpu2KkBtKvjhXQtdMv1hS
ac9di6QeDZtxdJAP/D5fnsdmpyF1FEPXVXmk8l+OIQLpom6AajHJZnswbmiuH3LxsRiIfG1sZ7MU
75NADTO0jxbQ2v/9pK4eNjitxZXzerWHkJijPuwHKO0zn0SUXU1ZXz1IapblxddR6Yc5dMsHs3TT
03g/q1FJHsUeTk21oADHJu/9/jdt3/2SO5XRRLzwP1C7pUKaXX1NI99QQRuy6xqLQh9sNJGQPJzE
yPYpvZFlWnPC9S4MH7zEVed6QN9jHaz90kip+smZmjI1CzE8IzbpHyof/PspuYAV8A9YbZDD5T5f
V+8jNhAT7wniglriPqUQGWjJHcP0U2EV8+5fpiJuxVHa1F4R+NYyfCqx2W/sja29qwWli3Cq5r/T
3ZVnleHNhBQvAk0QvLm4pENOsmK1V+N3cpRbTbeYk5JOa5wEqHcTzmAHQxb+C8uwM01K2oFsgOTm
nx7osy+n+WVmJRXY0C1CvffkU9XzMARBzSIapQLpiykWi4BHrNfj1tVjXFqG7p5Q28ZKHZHIiqAP
+h/KHc3WHLX2zjxkKYASgBHiN+vZIUE2PkNp9jVCRUfp7Tnz6+3Obk1Y/tqz7iBNO2aP2OEpWyCn
Rt5m7tLLsJVuMYoJdqrnuNKzSkE521ZZlyXUFzmX73JifLHGgC5A7DFaCKsOWXGcQXkBK7tJJfte
iy7SUMbFRNwK4dscPFqh6VofXEzZu3VIxuJ0W0WsZStgbK9RDa20mkFy0RrJ3EZDYtqPN07q+zy7
yxQidg2Zv5ue5kMUBTcWmlgB902m5NHXSzQSJqoLIVzD8Ov68xoc0XIveKIo8BOFLouY3KTwZNQe
I1U6Yyj1yHGq6ywWY3Dm0LfnmiPOVDrrBk2ynNFxfA/ggsjxAWa3j5up7ToOJJyMwNyhIl27qYPf
wmBJH6EJ39/Eyxa8192GJ1JxvvbUOK/WlSp3DMriCxTRAhA4yAhpCwcWYSCML6UWOoY6fuIvpx3j
mIuKQV5Af/i/tMq+nbhYZVZ9nx9qiS7pj9QSiWDaeBSgvMfuyGz7tXFBfBHKsW6e3Asg+32iJCBH
KiFRBL6GsvCpagBqmSDt88r4iegFL+qgxsuOhIFV6TNRGK8RL1adKFR6VFs3c4O4TklqHMbYNVmA
ofyLUvmv3g7m1p1jdKX8UaP43iRGXIHkP8F23WgAaHXGa5xAIcbfGlns1Yg4q/+o+mvXQ7YQefBQ
+bwCl33aMr26uuZ0LfobC0p7ze0hoTKKHayhzRHSkit+/GueWcw9tJBIFsFqgVYYLSQgHKWBdLtz
k4fD5D5FCfjuwrfJZlGl+BJmFU1wjf+owFFKzPEyIQVTK8rNhlPZGspd2QNGW5cgWjbt9U+/3Dm4
0q5jdEWCgFin5AfwMJFhj18VWUdtFpOiLEqBIA3Dtbwu1KGhkPMs1a4q+aP4Sjo4f+u/uUdxBXe+
toOUPWFMNin+ydvokalplbSKV88gtvvASvg/6bh6sF1Qi6fAv7mSjfZhHoxWMSL3UkCXQueLISRt
iOMaogWVFk8cwRsl8cGQYRHZOa6+jgy4at6x/4ZRO3KCPpIh2ImAPM/suXdqi9SJQuTlNOOsgsuB
yIn2VSmAjhUY/GIdSzY7FDEDWQJwtdZmWl4+U3eNkpHLgGmVIMS7jiE73+4XP9l2UO37t/QxoPxt
/067WlqVlNQehoJlf6uqjKfZdmD/az8dl7VMn/5kkVeMbczmffPz4LCpH18LmbpmKAYp/60vSsgF
5s+4WyZddzpZLrojRBR4nfP9IFti+bssVDPdHRN5Ku3cEaNt5CIJiZ9IcyyCDKb9q7yu3PE7ryWU
emZR2MIqpjZGm2r4foDszt1Jlm0A0JZPxJI5Byd5Mp9Eere1xDp2TuXMaggG/K5NMEyfiqmUaiWe
R0mO03YcoLqk8A35kDB6F5gsADCy3JuhD8L13tCbabc6XIk+OM0tLlA3SBWTGWWY9oihnxumi0qq
DhDAFqLmR+LPKzgCgz0Yz9cyXH8En7nobgTfneT/ULeBTU8/Sxy4rahSPUbCHC4P7fXonr5HdseF
W8HUVRzQf7dK5nj4ajWkgj7oNM1e6eoRLuejWBSQdws6TK/8UffAA5CYvIce9x8f57tIhO/UBmmS
sMXXytbJ2ovQ8DyHy0hSsc+Vc9xPGJMdNgUiLLNpYdvpY0OhAL008/HyK6Cqb6aSnMzYypgg1jVy
g9wDAWvFAAcHDPQYvl91LMEGaN5mL27VFWWY3RUHAKVR2NwPQbtL9k6x6Ce1WPGwkXTpTlvFENmW
iiQKbQWrgDdtUZNEXU/R3y/FrJEgTyTahhBk4WJFSSxbE7KUfALD6VWEjILPXGpDgnEEm3fM0TvD
MEb46ZyG0gd5Yq5jwECu8ZfO8GkoBySXM4DDrncAzmY46kPcddYpnLobG4vZJUkfT3PyJEsbF4mh
PpuIKFupPfC4/H4scSSGuZWGnsbdljZq7PdBpnhNoZ34PqDsWLKsJduX7fyCgDG7F07Tuu1CxgJM
rT6YJYRM1vRYMnZSQT1x3MowyuOs6pF1qAY76KEkziYxwj2MI73YUZWHMEThAARIBOnMwBGB5m1h
63YqubwMydGsEV+YfKIOf4BdD9zFBJKd+KR1mNQCnYuvE+zEc8KIyUFGGf+UC8Zrng5SC2U+kM4w
DhnosEhrdOVlIXenYaVtqAw7ZiR9RGcsVxxA5T7Eun+cuHXf3PweMmovIxizC+NTJXiTThM7+non
EzYhi/Zwxc5O5jtoyBmkO8YDyGnvj18LlifLUv0p5+Rv90v1iddTNQPs//2TkTgi/0g/760HMbK2
YYmJaaXE+h8JPOZweeppUPZcykWOEApRiErWvzPDxIpsXBzfZ2kST/A9XIb8xLCq2HjYwA4y4LeR
oqRHZ0gD9RhAc5uc8ukDedN+ekNkRFaXcaoloABa0SGz7+fD4oQhAdlyGW4tkRfzEwqrx9EnK8ZW
yfPhGpFYGFNznUeY6r8DUVH9z4da0GlKvZQbFJksR/iFGF3rDuNjdDeHGUfJH+9asAFo9kJgIZeP
BX2CpjT/Mq9JK4xUR10QcDwwEUOxtJBxl27l9VAkxLG1Q5qRF3m2X91HnQqWckfg04VEtvyM33xd
oCYldrSRFtUGx4wZYANoaCQwhOq9hS5WHXQ0hn2611ukYGLX6Q1jExLId15KrHNOQp/yZYM9rGvM
XX+FfLc2ZhpC4lmd67b8jl6H+mdOhj0fkEN53cDygo8rLIZPSlDlXp8AtczSI5qqg/BBTxTveIBH
1zd7UqB+yxqYwj8V5BSWhmyfZTEtLFQpqXhGqilgtPyiZtrbYO2hyU8qjhdQJwxZxjDOOdktU1Pt
PLwh6OuO/b4s4f7pLnKBkoaU6qMjSgXucyPoI7DBiuQkWLXJueYxY5031j8ndRjwKXLvnOgGRX1R
Md1kAToV9ccV0tFPrsF3ItxJwDkcg8z+FxbCmYiq6FCjwJ2c1SS+VY8UaKm/PsKkxzcuSllVycuT
FolcsOKBLHnD3xS42S3D3i6XYjrQPVFWv9N8hEsjTOQ9ykqSyew48buyYIaSbgFbtH+I3G5YrXsv
UskPZaQSLjkA2gYI0hToFExBmdRUFjAIoLMjW7soS6v/KhxbkB+1QjpL7nsuzfBD+KE6CD6rVUT5
Hih1Mc/gfGua2ohdIeyGOgE5r0bRFdApLDU7PjLFkuJOe2dPM9jaLSs3Ytrtt4RQBm5B5gEudn2D
YJmaiLiVOEVf4IGTcrkipBSzjjUqkIrseKpsLwSj7ChnoLHBxhkvreocDPPdSWkoVzmiB5ym9gj9
87wFrXnwYQcg/fdWYqtNsmdBErkrJ3/nql8fRMn+yKKMuNfAQ+38JwK4TmdzAOWqN23DrOVEqUOH
uztqVzkvoT+K0USPIAVBy6bTLmEieAsuhfNcJOhN9CBGtdGT8o6hnUv//+e+oWZWIYBFV7gnl/+A
ZQL+HciinLcrHEDcadnNYMLhMCLbnGx6P+yPrWq7UPiwINkQuK9Y4HP1lHlXZuApKjTqRZxKsm1g
XztabmzVPmf5ZE6iqwkRM7INQ+9Dc+uwC3+cJiuSUW+R73CH4RMypcg8FRvsofPhpRIuKfmTIHM4
BKlvX76k4sa+kcGd1Vx3mkJg1DVtnh18MEH8NXORbpT2RQByYEYN2nobanvrDPjs7cJIaD2g6U5E
cKtMtx5L9/OrVYCv7JaLI5Jyfu4Y0C295EhXaOuyh8JAf8rkij4MrmsCf34D6PDxT7ruAmkCYaTJ
9NaJQnudN+uDOkTVHPTblAX/ccmuP3xuGbCDwkpKPkOskM2QcciacSBhCc9hyL3Lq1n892lqukdi
XNPfjZ+nKQGcp3DokIahdtPYe4Tprq9dxBn4jZj4p0NFAKVCt7mErIt4jR9tiFNHYaR5Htr4UYvp
OEpyntEJxbdtwKjjBPgeWQr2eSx6to+KqFiDeEXlgSf3KAzEAa2lUhv0ouk44BtyO+rrEk1xuvkJ
kiTEgYN0PERES24nqZBj0jp7txNf0Wv3f+mKO8Bvx0sr5xIi2YdlFno23QsUeu8yAin0Euu5T827
SWWqcY/oSuQwOVfwTBYslWiYb8/fnqLrAcQkW4f2DQoNkuKklOiRZbhrjqd4gpqRMd7i+bBue6SY
+hA0RY8IJXgC+I6Ce85LLMhhmakdEHPOrPmHNR8fH+i0b9F5kEC8VDLIV+22Fx69OSaGbenT6sKn
LIbb1P5nDU72EWBpEXQ/lciK7R1hERsm7CLKKBiRIHojxxH5+G1M8fXh57/qHHAYvm7cwfx/u2T5
sumSx1LF++dUJ/epel2o9oKx9QOlr+sp8TCDXyjtABbVLdhveh2vuG9M1bJ2BcGiwQMTRt1ZQnwI
LZbuIswBrDzW+RBvSkDJzHn2nTWtUAZO94S4Sve0joyBdrpp/bsCNC5ChtDnlZydRY7G5s9wRJ7m
+Px+D8/XdeNCFUTgAf1NRb9nFQ0uRrJW7vRDLT3wdvQKeUOj7LqddPVFc2uA9sM8+pR3FJIjV6Bo
SWrIBFtqusWKoaj8mIetwE5aQud4LoAlceHUHHDERp2YKZzbRqvgimKDaGVMDsc5J/neS1a49EE0
cLwBqMDX2xgUfl/kQ5zancZezbuhh/bObHZVROauCyllKIxIVo/mAf3eTBT0rlZbOZsumEzNAQyR
if7naLEjQb1tdtt6my1SBf+UMQgf7I/9aT8GKfsROJhxg/tuwPPEHsj9uiJBcZBhVSqkek6Z/WUz
Uyb9RYdsxD+u61SBhhlSVNLbvqPi1sL9G/sLNXhM0p2E8umc1iJLJ0apAB92NQc+zOKeqR0Q2jgT
idCQa7wBV/rmQu3xLD+y9RWd8Vjzb3jGLmi39zkTqCTc+OQDassw39I9RBa8JnZrxXj+Xs2+gLyB
YrG2czKxD9HUPPrn3enO+B1yFnXaNoSfK3jt13gYESiBLW/GpTpwsYEZeTwECDLYFOJpxmk2XQJv
8XHQpi2XuxZP0a5MRHWZpfCt5QrmOCl7UlnGk0HREYaGIUK9oN9ILw7PAjnYxtUHjcjfU1eSh2fj
qgzlMbt/d7+EeyE4lissWfEH+39suzjKXuwL/Zc4ZSunsshrYJBm+1ARKbCzOJABGAEN3CecM2Ru
bnQuZsGEQC4jAjbE229hk+Akm5q7qB9PJSYi9eSPxQ58s4mnrgDpMLEMNUKd1AqmDcP10bAcdu9s
YbfV0YNoTf3cse574COUppsy4c3lq3lznzl1B1FP63lJWeYGApC5wIhjgMPIghFnG+z0Awfv3icF
jVzXtRiTuuYeEERtPdXKDgpxgg+JaUe8UiBlKNx2fSEoSiii3SGjbKlX+dIab2nbNu/mhu9zBN3s
VmEnFYQU7Kx4u942pv8Ugpa5WTIcl0NyCb2tRYFJ3h3SDUWc+O/8i6wUuVKWxyrOt+/3ol/ZONxF
opU80DtH6Yw/bIxNjU5Zo3vcb7c7Flom+aUEIex7WRgeMLFZr62U2xE9KdTdodCFefHSYf6VJqat
OIbGfWWR6lStyQcA3OkprIBCpyPng0/yh1A06hJZ/7KOfozAbmC9eaVVmXpbCap4EgqwSNkslGdB
PJ4aVxymxSdkkn9PW7Dvi0jutSWaCs+Qx8uixmLzbUzXH5VJ5lsMPVQZKqxg3Zxo2aIvYK7jisPG
G+T+E0soBQPQBWIVfU+SSXfH/5DBAVexCkFRrHYrFEiVlRcUBTbIrD3yRZSp/zoD2sXQFJLlYKxh
dxFQJDmlPPIiU1U+IEST8M22P5Lnf019CKSVm/Ebns2AHAth6e7eBDx2AtG2e6hrnrOdR9IlzTRo
L3fGXb+vijwqIkYXj9p78kr31eP73iK+lcNGbYUnGXW9Xbv1LsfuUJIsDgTf48u9arGM5uUkaLTJ
veK+NeOPdyNbRYkxm/3ZYOW63+3UdL209cwoahu77h78N/OFHeVSKQ4V20QITNLBtdfdofRYyhnn
uTmqlYFUkz/kLTVgW+kXafKl+5k2Yr9PBkKjVMDRxgKKtpNLixtXhQOfJcPj2u4rTGogN350es6K
/eHwrcig8GwnHqxdfD6u05KR/X8oEKLUcFjC52R8ZELoBrNGZ5L7BdqS0jxu/eqRmVjvB/iP1nqh
Q8fxUuLqxk2P2prbp2ghSpZ+dsSj1h60X0VyHOHsRbjokDrjJsR0b8JZw1N4j8bm02vLn8lQx/Ox
/NisAPGL3I7bm9KGlD3IQmTh0gEjeF7CUDloTF+6m+3hUcE9t6ICiT/tjSZ/tO++OGmBw+dLJBMn
7V624exko7QqYpUd/t7vqw6n5QFHIflqw1ugkvw+ZajvfkqBMNMp+26KMnUrZvLQDCjbtXS4uOr4
FnbBX9pS5nTV8qO2jDVc46ZybFtGRDssF1gSF97riPdrpJvT0n5m8D78JjsjrumXNaxEUuqzJ6aG
DYHirjbPhY/eE4Hb8eHlz1MS4D3sieopE6JXb0rSOFvYY86Wkw3SMIhlzosfYPuBikJCmaGi2s5D
jsCPNZuQVrBB25SM41dRo/eZVcvDC9dRLEYh8Hd/ECXNA2xdSV1+KmL6+jj24Dl9MTT9clag0TAK
u8FFa777t2ZssfW9AzUJ/CjMh+yE4CdmZlxEorF+MMt6F5jPSLlP+hsVu9wiMXhgYIwYjIqBXSmd
tilH6Hyty3BnCnJUhIgSXdnuRDaDalycUKrjEasiMVySP/AagAPrKOZs17O5pi1ut7lTrwT5M9A3
IgdwhBBusPcqQvPV/K1fe1Z9H+z16xRifC6+SlOWPmduowFXJDohyJ7CxunxW4+roxtd5S6JfYuG
0kNaXAxB6+ZW+YA9LdtIGVhFxsCwOSDAsMJJZYRtCWJgB41FRqAXN4uCT/MwmWXoMWCOEXx6c+at
WgpcwJMfRJp9mN2pCzPy5otpehpy2pl/d151t9XnlPWlnKGBHMbCxfNMm/V8cSX8++JeCWK8Swfo
oRpNDjj4jQsfrW9taN+hX1lYsVzMUvq9KkKVeKQssDSgR37K9xsDfnknXc1ECvjKT/dmSQvWGGbL
X+/2WBzegWdecdRrY0OjbWjpROiRg458YhVpx7cRWWCqNiIT9fc6On0MFLlrlbZDDxS197bpmlqX
0LrJ6UMBQcitYAvPGhHvGIwiTZzi5+zyz0ehaz93U2/XPxkj+uMMkZOYR2XoUtqSTZuf+eX/iCws
LB2lzcPgnEXmGeBh/8RMjC1rkIB4MwZVxIpUHFg5g/FyX4gBD5o6dLI3pazlrtd/XKcQq4g7PIDu
BMEz6TXRZ+w2BZez19UAwibvwCTfBmaDbnlU8Md/LTPNO9IHIGooRXF8+nOsTR+STHJbh9Oikx4s
neDIPzLeBrMMhNDNTLdTEnYQysgqWMa86mlXWxtrP63gqy4gI4sUoU8ngDy96cpR6oE4Ytg7Uxpa
KRGIDdlBkhrT6EImB7disFB85WkcnENCh+Z6TCA0RiRoITxuQbnHfkKtAp8CcdTekFhxs35L9iu6
yM0Iwk6T8LzOj7EBPD+3ale5zePNy23c/VDxhUVbBCcJb3R2Nyhp+ZFvR5Afm5Qdo0CHOwfkvRr6
Yxh/wUYx5MKA+pCNtKiIajJEgqZ63PLTZfrkJGVo1ftt4V6I/n29u7OD3WKIofR+QYiQnYj4JndH
nFrKWHJKnuvBIIFdWf4R52HzNCn4X6qvEEs/DFT0NgxQAQh9H70R205xF1o7tdncazS9muM8IkCP
KHQaM6ffol8hG+q/Uy4RnPn50V7sCZdmolJwHijIQ7X/eDUuqAUWpWSo97f/fWUspztuIzK6RQCX
G96jTLf3TH61mZguhlej4CMa8mi1f59YgDwl9V4ZxtGYl1z77Jfh9tgDuq0KUmNVVB6fKjcbgZ19
EoIIAyqFnxPPeeqLansIiwfGDKRwj1msn288lAH+8kfBuTy3tUs5lWn80mAZ2DUSQ6B/9/PPueab
i2A8K3oK3oXW7FwsZE4HsGEi9nmAeCJRHQuSPl67TYhc0lkkbGdIbJuMGQCvfrwalkjxbL0rai6h
x9egmXrLZdy2nENfJGoGg+dx+MyzoAAxczl3Tp7FWZzkxwxi/iMkGwTb2n7r08cuINvic6/F6TAN
3bqr787BAorzEV4R5bVg3jyk7U61dUT820X43gWIynJI0OK2hwRo+KvsOWOkZ/UqER81F8ymQtfP
XSSnvDL10PlHryQH51SoVNqsAG52Xy6H8rLK4j80GrbWTkzSPeg1d8hig6tsDRJM8ADTEYvDc66t
3zKEwBj6Mp9PVeuRwCpRFRuSn92nZs8Fa4SPQEbc5+rsnMWC80HFECXIg1p1SzUAwHCUL8mlG6u+
mZtaEhCZuASBvOlzIep+K5xgcNtQqJ/V5vVb8Upaq5FBbas6m0ErkVC3/FWhBOV2wCKcBhtZGoB8
aBnPFb4YrMFPELPAFbtWoLIjEyxxt5/SKAfASWuSBxfrQSkXgQlvPmFdMK8+KIDYE9rVU59TWKFS
q1Epn1S3utgnZIvf4vjWFdXVXcheXmiifV4VKfqiWtld5fXrjaHaTz6y7jUWFDufAZOzFKuDSa0c
S+zQlAK4nFMeB86UxwEn/CP7gPpoKyzTtlQt4GKclm3NDIJ1SxIKjF1RSWdfjgMN5SglEPD9uLXt
M9tkZ8Z1J7E+Ow8iC/I1U3I7/O9D4jhdX7C5ICiGRMh3G+4cOGxP99s071kJdh6NFQWmX9EmHonC
hm8A8U2FJEQoG9EYck+P2c/EE86ebAcygypc1jzBFOSrBb/3/4WVWnd3YHp85aNV13Pxm7ghUd7S
LCpExQVo/6/qLfArDj/OpaqmGsGNMWt3bT/7pMJiQZa8hde1qdwMhPVoRyTCPq7NBwht7MiR52+l
LG+pC38pQ9AzdwcVDMWFAWehBrhEeLDHwUjd5qdPTqFy7DtgLGo8R2cqODo61vTgsrKT/+abIqit
mrLNEDC8iE4seuOjHPleouDvl3Ryw947wtSJoE+VrjYVe6MkGfjqrIcrM08Amg6tPTNUcYfszq3F
Fx9Z+L98Xun+3BS5bGQcdpWnVDQWJDVthKvCtQTVIlVY9DWN5j2uUXDAGhwTYbZnBHzogQHm1Muq
0YEnmmtc6eTkONOxT8YYkROpS1E21auoy9WOHv0pbKMp01dIkX6MGicPYzDB4x8468E8cmyDadrM
5Jq+3jeKGbk7cuJygjtea99WUQjJfBIfBgZ4QWRa9HLgkWfNCmGqYwynEA+BhKyzkAAzSaLp/wqZ
eLZZdB1GfiIITh+eqedVE1bar6606ccbOQGoRU2sj9+Y+vCyOjdDxbRIXVSrCOKbS0l+0br9wPBM
7Mva3JV4NY4wIDEypzhwV1DzW+IyJyfF01s05d+0OCj2oMf305lOaR15B/H3GALsIBi+xnEp9WIU
5TK2u1U5tkEmNznOR4Q07w0c/xtL5BSM7d9ItNOzEFzUNZwunPUhb27w6R2NksUTiehCfp9eep2S
dxbCHlp67rMh/FKuZJTXNHwj1kcA/HIftuWY9ErGe5Q4qItEXZmiNr3fRQWnKcLE69f3ihhb97OJ
RU3jjGi6oUovs1133pMXEXrXIvQ2s7ldg7mw6Kpd5W7xXmdLss7Q9S78MNLkodZbZBEzofzvvtPd
5xTPZqgf1z+lr37TGfIE+ngtCP/HeJvOqaUp8VdneALNcMkn7ZWJn48ZL0WLbGTZYOemH43l9ahe
zwy/j7xTylnDdfHpKD/k8edVcCCUm3eAoiQkmOGl/FO6Le806RnYOcmt0OGf4O24fy6Vqds7o9vN
iycLhpLrKHr8hlOGIfSuXxqk5HAM+7A3jO5GIayHA3xlEdK07CV0BzNsWdEuhXM+1h7mnB+DjpZQ
8uANyuuJziO72USGi7ZZZ8bXoLs/iX0dH3E4dHPsPuqgG7Lb7oqjW/bqFw5EofilqUVfhkHb18e8
o71sTrwDJlPM+Z0AtoUy5KZrEkFWruaWD+yhUPaTJYIAr1bS3MXlBPOU/jStIbSINxpshaq2DKxP
+pPu3PGohbv5Pstsx/Glax7iw7O0PWYYxEaMy9Z4zgsbcVSWfUqRN8aL2ZxqLHTHKTjmZTroA3cr
eIr0dM8LqF4jlzR2KENUxwOCpjPQcHWbWxmiBncOjjCgLS3rpn7e8iWPvfqRmJs4EIhTRyBbyWo4
8A9RG9XipKmRox0KgpeQAjqbM6Sd6iSlfDiBfrKoLvNw/quGR4cuxZJVaskoSAvKN+ruw74Bm/sD
jGt8AuAQ79vwqOV9rnyHA9hmlTo1WoJ5iw6XMEvkSeUmLwEhmtTDgv/hPwS8szzx3whVK99se87f
Ak14O6QG+uI9C36lBn6nbkroWTxNwsb6Jvdd0TQ5CUn+QPj3mCQ8uzQe6cZvQn8FtjWaDwaKqQrv
XnEOPDXtZzixEMNNm+BiezKa9oBucDBg7Ek2puFLtaTL86nFl1jOZ1LuKybMN7bqgpjO6sZgsow8
J20P0fnbd5mXyecjxcd/asuoHf+MTFpDDonm29GaC+z5WJwFun4h3YxXDjmypc5y65mfW5mPP4+N
ljsvr8H3kwyuh4Mr0UYgiNCX9XN65uVQf9S8OaSvpmYL8wJTnIyC6pNSUYnauH4+0TjTVFlZAVmc
dzk5Fp0W+kqDyhC0eQyimn6rlif0fdiNTIg1NFt5yrSZoN8Y8XwGDfLTE8ExofXi73NHoggaXtXp
3NHnJUwSIYiBcLNp+mOVox74n8bPUj9CScc1AWlWGf5hCFHgBI9gh1zWXoQwHztbbhnQxC/yUeja
iGXVJy+UcyCdROYJaWYg4QYQ7GddZq3UHguq3ZK7F+LdCq2dhqjfRgW4ofRTiIAPjphkPPHDClfE
iXSqGL1abcBBA3o6P5b3VvRvyUj5HqPwoN6+tmYvukRxqJHv1TZO6HDapdLj17c3i2EBHyi4BxqM
pHz2O8+ON6HgwPHyHhzS1gMeU6nV4RRR+FQzH6Hf7gkzmh07Gd14gSVP/qvND4SJuJ+yZD8Xt19z
InL+5KRqfJGHpuh8DFI22/+qPZfFIECFqYHN1LZv5yCqRforHpUzZ2miv4foYJm4fYl8oGCnCYl0
T8TkHkpCMXlYUrVsFrf5tPF3QvovRrK1elTvNcDKn49WoLmx6aNMiN69NpmP50wpXWagO0oEA7xc
dLvrKWDHg1zcifB/ERGV1uilI2nJThmZiIQGN2wj87hBqVd5Nw/YBU72t/12h9qhHzNO83HR8mOo
63LbCMC/CO8sK6CJ/b65chC3O9f4+11tVIycXHoo4MtYo5gAD2RVav28GYLuHpve1cUcMLw67jRl
coYe8xiub/WkvuxXeemTZtURdOE+47/Cx6LMt75Kg+GQ6TPbtoFj7uz1jWTUf7Dm/v4AGttbZMXq
1Nks+M6E1rElLddsPcCQECyK5caAhZRzEZws2hurssbMdGhoYcKuGJ9UOIQoyMdcgtt/miffIIb2
J52XLU46Dpm6U1BnE37O02+7TxES53a6Q/M4GBT8bQuvErm05fAwXaJFSBClMPZldlVx39OKTBGy
Y1kjEKhxouci9jRoIdlmpU5xEfLEey8gXOCp+XAVaosTmejhCABukIMBEuP+OB4wseLc26GjwGhj
YydwFxOm0r//AYdfL55Len3c+Yc1ZsvMZzulmSvsQfFw4ntNJmeq7e1XUOvid5zTbMr9g3Q91wKn
yHhNwWFsNBGSDG805vWWk93s7kB04q0sTVLo4MzjDFwpjQKCHO44ALDnIHLnK4oYgssa+xH8DW2A
GFwvpxwh8t/eCdl/yr8p8irNQfRNno62+LBXyrYtecE528ksIs62p0zUAJnLpZwXcwdCV62hXOPN
kDvIijr9zRb1/JcLH88G9MzRVuzkWl8MAZpwG3PLBLPH2UrjAVXTTnDVHyrfcxY/ARbucPWMEFDC
Hh4zgUWtIMmu/YxD1pyoWIOcf0eNMzs+2lneT/SEjCvRDh/6GymkB62e6CnAUeZ1TN8L0mXDiDlu
wvbGOs077RKGC+u89zVmDLGAj4Jh5k0zWGZAuqZW32Yi+muEHgHz/YOrxd4A9ahsVxk5y1h8646C
n386FrWJ6UaV0x28O7CFvZNP7Yo50nBgj/m5XEEEelp6y8ve77bv7X21NRrvrH/UiRQr4sTuklgn
t1eCcpokXVkWTbTqSuQLissLUwf0bPWzlhQ8pIty0NtvCYqG/B7WcRifvzV5n2TuCfI2Ve+YPR5X
V09su1WicflB9Do50l70uCqINEl/cEP1gJpLoPm88opTaBAtYKIbyo7NSS1W1r546tMAgYENbKUT
EiCyjgvgruoGssbujRs9gB88OiLV856D7rE/lQ4LHMZ8SBQL4BecT7AcMXeJFfLMf+DjeQywUppx
13RGLdl0Gbt8zhHKfQzfQ5PNahFWKsujz3+y1u0kKvBTgXowIOLXGukFjqUV3/fDbfPdI0KUtnEi
P8SERhQ6LYQ9G7jtB++zVZTPMiR96CtTTj3fLQmS1BnHn9ta34gfQU9oWggbhai6/mEBGCxdTqL9
/9zGST+Mh5gel2CF+PwC2fvX7tTUOeih7t8K2M5JblYiDO5fxgeMzq1YgJYGW51RaLJeYXP2G7vv
QE3zbrtwy2F3bCncl/7WEeD4q0ZTmLsVr0BtJv8yb4U6NGZEoPE0AVSku2ZQ01K9gzL/y0LTPNWw
Sf1NHy7Oh7SCgycnIbryfY4+r8uxlp6SxXtgGnlTLlOWe2Je2gmttNI7SggqEVtJbvMhtm/6auZF
th7rzYEu1XmYcpoW1pF+Fb3i/ZfH1S8g/d/dcbeUO1DMv/ypvKbAh7fOQ03RBt054VnAXZwit3Kp
SWte2RWZuuMHmYu/j6+NCyzswzNBaz63nal0t6yWPV7NEVd81sOAVHIAfFdpYsu84dphbG06Ffa3
ntqUd5PyEymh6F4PzPKmYY++CilEWKJj64eQdf+Gt57nmavoaLXM2iXerKov2oj2vGrI1UwevHuB
7BHjpuZ2lN2WQlOX3pfejoGg/etn7sxk+RJ5xLjgNWsIRFyNF2WlGuo0ePRUVahlVijqWlEJn+fS
T0XlwI+2N7GOlr//kpZKG8SOPhSatbDPgFwOV6hC/hVzPnJdjZQQ7CvppLjNqcIE3IAkH7nxNaxo
KbCbo3aR/LstKtT+d24xkZ9W+Lux6X0m1huPDDal3APJagJgKbl4N3G9XkneUzacGmLF/hgDUmEX
e7T0agmCm8MsIiZw04TU8cv6rr3nV1ii8gpDlxU9frPG4EUT+mtSQW4h97/5ONfoLxNj07YnMH9V
Y266aAfmJjh5k8L5mxTvsP/Ri27jnv+F2guQZ3q4Jd0vX1gVZFbwFlWjro7of5NWvZV6100NSicW
qqHip1wKEWWTvyqIxqhJ17k067tlKEo369p889jnRxCvEHn3uLyQjP+JqKnPJSHxv4nJjj939jXT
F+QF4BZkMscOK8Qk7b72r+D+/ILPkUON9o+CgTBDXmms8poTr98ScpkaBsmw7Y5M2OrCyX1N3vuH
4bSlGDZ2ClkH5Gc9/QBS6Dl4FU3j/yhQtYS75C8wg6kgC7KVjL5n5jTevXAfEchhdNC42JElTPq+
P6MXdF9d5ace+59iOVTB8sqBExF6wNFT+ScS3c1M9eNUo6di9GAqUHROHIdad9Si9dEq1RMpv9/c
nzpOhhJ3riG3bYjDjGxhEGMQwkTBMDEcwua5zoW33tNzD7KxTUFojhg+IFTpaDlhgDXiSg2mfYKg
+bXHMc0dS0hWwS7JYXTuAYn5UT++fANbhY+QHYGdFbxE9EhRCgJLWnGgsuC47g0VzqcWn1jOKFjG
Sh4VUXR3BoKH3hZf2X+DvSwt+CvtoZ4Lh9RITWbWIgDAE+Nibl5dEDn2BsihwrCMUcCCjGxr3XG2
/Wm+4UqLi3q4ZMzIFBHUxviWl3zlBIYt7rNnzgXVL6FQmHixDVIEnLtyMzKGs3rAMn3NWhLmBGEX
BwB+nK6z01u8FoWY4hTKG3CHrpeoPj1BiF8cl5ANz7bsxpXyy6CqOqkiVp/v3YxbI2Lfw7ABL8ai
f97+U8Q00zLNcxpHCsXQNM3QJzAgV1zFLM2hljMocE8gmrZEd2qyAJzN7RNRkknwPDMP2AbXGeai
Dq9syvOlqDdXEAWYZZhtHYgP69PtmogguJOfqXbcqL4wPdMQfIDZ9S3B5bTxitkVliIhHdPCVCEM
JQtfO5aU18e9itkUj88Ne6xhNJ7a1JhQoOI29cYAlRWcGaFTmYbP9mLRmG9VblhhEVG4eD0NfkrK
7rxJtcM+W84Fap2LN+1PK1QuFV1gvuMZzeJShsdMMyUrRsDJ7zBurZr95FClgaSg6r0ocQh6RAQx
YN3+WIAvVy0R0UMmHbBUVr33j7xwAF9wTesd1BFIKQ2Y6xLgRY1ewyVLTeiKUnr1raFWZ68r44QB
4Y1M212+NWW2eKmfafpbL5adUByzOpCGTQEx10WiecwD1r/TM5QP2XF8G4+uunqTAaOpQOd0wAp+
hS7+002IM9V649yTTOKMvQw87o83Yx00cpsunKgNB/xKu1Ne3VQg0BDnQnSDz/9p4PEer6FcNWV7
ZpcCy6MRKlvts3Zque/tvdxip4PSmqGuvcrMWV9aY3iZZHEnhnD52Kx0fN8fmAhpX3nmytECnx02
amRXz/HSG3cytXfM9n9rPCY9oP17jrMmfUcOH5qnxk79MnheH0pJM7iwspZ8Rzj1VHnz/7SH4wEf
FEojeB87bw1plAxYK29yQK4UTO9feuvrXQ1vfi802uQR0I1o0LqVzhwZh+xIrmB7mplg45za0/BG
y3THCyiHl3NhguaUtIJJu3WRKnoNnTqZrom+GDyETVj1bcOwEPzRWfRuJNy357XoLdfbsSApyeUq
GyqHzM54rC3oXBYw3X2qTCy7ncPSXAEnU4Y18jE+cxtczlb4VQ+J6Zmjt5vmMAnvt4TRdYALiitc
qMqSaysl9jejGW5zv8pX6DlqI/sdhy8hUni+3Uq0z/h2GzpuAkrX9AhJjIN4xxEjKV5cyEliHj57
cGuKooYbCvmeeczZNupSikDF8ydiXsv8e42v7Qk6PWNCZPvhaWDp1fmgLUDZ6DAb0RMdwpURj5mT
1CnB2FKXBkwEgUAITl8qv+1uwua2fJM90yBx0nGQsqxuYnVLYFgqROH2q4amuZBu5Jb9n821Dwbf
CBYflh4/elx5M2lC5NgeXX7nzy9LY6B8iAt7jtGKUg88LZYoFa6RLEji0gCyOjFc9p6jXgbNpoUR
DvugEkbPewqE32MQql+1EA149REGCh6LVe4ZA9e76PZN2kseFmcY+tBgdEb6BhGPyvus9nqWJvzv
Kcb2x4X1HoVNZCCtlJRBMMoD4h8KzDAb4sH4Opn42nFecWAMGLDBO8JS0OeKEfWdoOG42thQaLcZ
PbQ2LVo9mLTklDynYtZ968E1V6FS1fn+wT7w4zmbO54D9zLP1ROnYSbxw2yt32UkA9/YEar/mIU2
tHh/GaFsChtNM/Y5L6c4ujhDQrdl5ReCrx9dWeINzZzv7xEH+RJLlH1XS0EchEtT69msgFhcfxxa
CssL4tpzQU3Q1lkKdx1EfrQYGtS4s6KGucDuqTDc0c5R7JmT4rQ41fVK7GzGQ/rFvZZ1tK8B7fq5
+Y0gb0NJKpK2sWFxYK25OAAJ26yHr4yVxAwinsK6/bDpOeZiEAF1d+c7ben9AvQLe9UclZiunMbW
1uhsLN1GStUj47s/bx2zrxEXyEhUzpI1k3m0kvflGTu4yxtq2NatlBEsqrV6JI7dALpEXT82hh7q
JVu8vBvzY5Cn/HKCE0dvZcL0gsQLyxXBh0TAo2Qogo9pKLGtu1ucCeBqcj1eHEqP6iBLI8EoWxU0
6Aw7LYImQZe1FZ4K0+CyxMPQDP0wE1f2kvKC5AakeEhCZoTiu7wzTMUANr7QV68Vyz82/yy458nq
t4G9H/NtVD38wx85WmIWE/9jDHWDGe1ytfzZjWMwzderjbk1YfN554WNqeZbrkSUXIUfzNZQOn+G
Kps1T3BTsGMuNSVTtsc2R3jmx3BwhCSSbWGcOpq+0EXBIQ4LI9TYAgsoauiNA86IIdGG215WYbIG
zQt3wIbU9+SGcysAO6iHgbN6uYha93C7i7/FKSBDgalkNvtDCFX1IhiBN2BBqVbXkjhY8FSE8P4v
qxXVSwCpJlAjZa3HUw3qyXwEOtef8cKZnm1YwQyiS3/O4AGSrYe94aZX5ehmDC6BIA+NxpfktBPT
e6t16X81gamg7wKJYchec77FUQpadedrXAuIPi7TnChXEY6g6HJdoe0MnQ18or0lu/1dt7PUfCpZ
ZpJAWhjKd6pw+MsGTFU7PwJl+E4024kI70b4F8MMrS8cC7SOEcf0Uz1vKf6mN35Pro4lFg4LvBK9
Rn/nhS5tG6tJaJfBz8aJDDj6xsg1+KXGj4ZdBmiS9+Y1krdbEYna7QiPaPmA5GxV+mTF6k+l0+o1
LSJ0oZOdJe739PpjRbmW6tlx+hvIJcl81TyjXLNAMHB+lYuvfEqMRRmlo9nSalVyIwkFnFywKbgr
BAazNzplr47dASXd1myOomYRjbdMBLfbBP/Vh2LaViJeOO1sIbWA1BA5lVQ3haHSnM4aHtjgLGqL
Sca4+BqZtJDiQIeq8EiJ+BQWifJBY1joHLFJ321buI1N0wAAlvT+sr2q7eobWErDlkHFdxJXgiEX
YqC6LlVtMFRaImewtDzXPANWz4VcuiOfYyAy9PsLopgZFMAGk9fTqSCFVYgjaONl8eIhx0mza1Pf
p+8LehpQ6dFFmff20IJABIbVFHMshahwqt/+dpKkHsjZllMIOX+Ry6VvTp4SKPzN8usH3jjrin4u
N7dtJ3Ydd8oVW/bfHzZUDVIqNRVWGSoRGmHtcxsbtGQSCvbioljcVNimNlCq0knu++sfxnZfFimK
1IVgO2U0Y0pwUNdi3zWWmTXewW1Z3okscG3ig7C6W90t9RR3ni30J8gfW5WUq3BpVyHL1lidGHcB
aq8Jy2ZgICAuHJoKRhxeK3pv5SFBw5WUhEPowVBO9jnCTYwjt6rvgjDM9UJlrp2d1EH4frg4nHCw
FvfDxWvV75JzWv2vwBcTQ+dRSBXL4t4c8aYUytYyJNCcFeXRfCCuvUma/GoKN1TardqB0jnZ0B2L
s1idqQanXhWnOj9sF3by9Awnp1MCUk/xWIXwJn22a1pj2ZyZfRpelAVDEJcVG4vaVjvEhk+mVrP6
635h0DBML+b7L39EtKvvnQXuenoO0+8i4+F5Q+22wt+GeMD6y2Mv/MR5y2/ie0BJgWHCKxabC3cj
/FF03fWHbT604vngLv1d1fJ3TJCXdXKyI/jMYp4tUwyRsd0RRcJ5DPBZFf/ixx/V31HaHFNlg455
a7TvcPmxtnK4LkSU1OP4xoUJvLaWE/LamFW6XxXqOzvXDCY/pqVLgwCg/HXLipad5REyeLlGwdv0
rcV2lhgJd2RU+Jo1k+/RL8m9fKQG4Yst7g3cNHz4ZIJc3FPNVNSS1d0PcuWz/DuevhJ3c+a0cm3w
aksv6UVR9Z6boFCjynDGBTOdXz3E2YmHOeSMoGl10LOCsi3eBJuzkPrwpEDgjweiVIP2E+gncvMq
3YZlxemG7YNTFuEE7Zw3v2W3nHYV6TApBsHtyqjSuiLxUCfoFTH0vAG0jnyf63vSWMn1at+DyluH
UIUt97qH+k7EgDkc62ZrIWvcZGWKxtl9EqhdANr4LxsttL6z/iicKLlHs0+4/+Dhx90/2GEqa/8T
ykzzWdxuRKZKeMVaBgUYttM+jksBaymUtcWxoLcoxgknwSl2FJQ1otVUjxt4vb+5rNyxo2kmvayn
6LuvsubT1mLUH8tka+zt1ZSo2VxwKqsphl//put0jXMB7z4aDBqnpUqF0nXfDU7syMP2g+HDslUr
iXnuzx8ROaZM0roKShJoZH7lQBYtHOcwFO1br5M/FXVGBjW8pnJeoBGWZMloIIABrun+7oPrJn2V
BW2cZqLRnzuqoJoVB1r+M04RLfqKrVUqN2u0jO2QOAt1Uy3Zpgln110Aa+exstKIFCb9JOxbvRMG
ok4TwAOgVCj2ELDH4RCDEedt+teG4XoL0mwm81l2UuYwirltCGowWL8Y8W5h40lyywaRhW8u+CBT
L1uEopSbtWkFn3joFGI/K66P9Yp4V0K7/MSH9sU9pGHQdwe9Y8BunXqJCBlNoyZTH/yXoai+oaXl
C9I1z1X6am4DPnBL3L1BMiJqhmADxq+ZViMReqTtTNj5Q3zaD9U0PCxQzm9xaXuOr0Eotz0AMM4W
14ptOdnY70QnDwYsC5Gq/4j+IE3aBMb+Z6i3WmtDDxhsUMlJNbzVeZqPYyo8DhnfS2tG3qJUslpY
+bJnGAxgKm2OJyeJAzQZDaneSpdLKcO1JiksPKd0b5iCq3ournLrnqN4fowG5XJaRHWcmhpITktv
A4h+gQUsNp4TJLIZigxOLW77rkglRI4H3kwcQ8LiXUFgRqk++EgQC7YDVqKH1Lxq2okMHso+A5/l
SxduPkvM9nh1WK6QMGa/JNbMgHS4ECa/1jdJYXp4a55+5wmgxn9AGTUhvOhVMA57BEx2erRPL/RH
SpVSLyODuvEHIK8m6LfBzr6vmwqIbWiNV6n+soHawDu2jxRoIuA+m4rYHa4XP4CL79Yswf0VzI+G
48d3WZbDPO1/PjgfjR06/7zPHKOpl+cZhPbgmXWhqzSrVsOuq6DgC3910MrRmM3tdHFjThPWHA77
dAgtCOLV4EZbCSgO1zuAiHpsrCiPwijbSipJV1/lpZi8tqWIxqPZCxVwsksc+bgPuOuLRKYWIIcp
mUleej/W/j7Emz4Z12bZLoA3WX/39hKNfk9gaiCxQMpD3+GWyuLYsXm5OLS2su9rrRUkhUGNB+U/
NxJKOBOM/Cc9IYtVv7VIix7sbLmCLUhoqOK+35xKbr6wgzJYHC5fiwlvDr+PYyfVpKJi85kKT4Wp
qfb0x6Cb6HxCXFyH+JLtAaruBgwdSupwoVq1bKKi091DGZUfCxMJC27LphFiJGN6AFJHSrzCF+Gv
xb/J6xErQVXyBx8aGKnDUZ19RqsTABWTrFJZd+ZawtsvN/4EDEQ5tQFYKqd4nd6+jaHUXTgHYPej
wNgocYz+G38OtvomUcZs/xxwNi7PW6JgKdLXaeC09RDGyRI0HM2Z/Y+sRxgX2CWl/UESyU1i696/
zCug468kOsMFeTZwgFeVbB8qiDYUWnr4MTz7Q/cLJqwY+8GqWZZ9PFKpPZDxkPBOA7thxdk0GF1j
y63c+y5XFR19KdZoOD9rksLF6+WVUB4XpVwbq6roelkkOevkhOvBKXofw3gL+9vpulk6eyEjse0g
k4mKoLoxTDCMJaRKD4IbXyQKWiP/ofNCc1wyTPdyzzxcCXSvdEFjXjrj/fHt+qn8jz5dgxcovkWs
F6JzX4nHoCz1aJteTDP55vM70fDT4hbvxidUAs1RGgEb5NcfS7st5NY1ryLi20AKGYcGIqMq/d63
J+1SRauo/KqY8c4dnYottS5Q5cs1GeyuhEFZv/+s1XDZI2e0ifTqgnQvD+5xG/f3frT87BE3JUCc
XMt1oG0kk4frA9J/bq8zjgPgSm5A/bC+wMPxK8xaRgXUO/GB3NzccYp84WzW47MpQpvRdCUKcrB/
R4HgL+CrFfg5pmbe5f4vi/PtDBgP3bj98D4JER7rdXujh7g6oE9Lo8FpJXbWA7Qp1biYfmrqifIs
M3DP3wSDJOe5pkIDLUN3HB8YDancWuy31gll8sg+mrX8viDNw6adasdgAlNGp8aib6IklfWbbENX
zDKqBeVzgUPjHSBDxiBYsgNpSpbuIx1T9x4oaHuxQA9Q09Ty3HZ9CXvNFXzl62+liH/h655Jpbwt
x736HMZfxBX7gQDkI72OTzHsGpPdMgHDWEwBm4U3Ut6Amn9cwAq7D4Di5SpCBWKWdij8lLwGd84C
jlnqa5krXj+uRektGAkzqv4icQB1dSnk91QRzMf56SNSIVe4JTLQzqcfJm7rpr9nX7L1kcq5qX04
M0IfQeN/1ow1YuW2lcLejyCYoIUpQp6OAqxGjzJMd82e2eNjta1nYKxmcffjErs29Du0nHjpjrwk
cOF7c2fTKST2gC+5bs9KEdce/uwF9HuFEWCAXhw0TbQwjDh7z5xCOFmaGr5IUMv7yFCYWAYgv4Xa
eR6xhN4d5993m5ZTfOwPuvzzn2BzCyfCF6lujYHhr2lkdSf1UpGHt80dJ/vx8IOMWk48bL9LzMjN
Ns+UPT+2Ivw79VKh093/Pi16b0bIMrDysvCauRHgK6bEfvo1YXEaUJ0xTPunvrk5s+WgBHG5dQRT
ns1bTeI4uoIbFtkWSEI90kW2MY+v1fVgJKZJ6/zDR+a2qzxkkh5W1AM/p9/iGmvkY4i3atpV7mT0
J+6REGGa4o6fR/c5Jv5hIR3ONlgPA4E+9UO5C9c5O+aGG59jDjomfjulbWmLQGhmgSRnbIemu1NB
uKeSpZT9zM2NevBYqtW4bq0dDQq7JQIDksAzo+TD04Z/SpJxW79tJ7ZO2BGcv3YjUJ9QES0HvQkG
6MrtKMcra6vg/0L7DmMH9b4kmQcnLpgS/vGl5OSAnfBXgZQJnGLp/85+BbBrnyLJL0eK2ueoGCFa
QqFCi4KoHYwempeQZ1xsCwDfplNttsD1hopHLkMBBVHILkju4QeltNYhHO3L/kswuLnE+X0gPn0b
xEJSFVyrvPnAXqeKlJ+dNQDpAwQ7QQnquXHsxMxQbDSpButwRycQTEY5o/Lhmqd9OwCX0fs2onYb
EPYja8dKEHSh2ZmjE0dsOx7U6cUAd9Ae1gL+X8UHuIEF0d/TG+SyBhGWOYvZg4PQ6K0hB4bKhf9e
ELaglxiRIlgN9p7Fp/2Km0YBFbT9pEm1TNkWDdx9z0AHiUGOPniCrOf5wN3Nyu/YIzipaigMmjo/
W+V12o6W8FnmuCQiL4CkuFwOee3k0EHK9PTxfGqD5SHYQ2O6vLHKlU4+qmw2KuKo0YoaPXVuo8FS
bwJ/lv1hV1aRiCe4vdgR73oYZpaLnmjrWDHN3wk2506S3a0PPDa738xgLXygaYLpTl3QuzZ/J9b8
fIUGX3RQRlBaX+qCkP4nWqjaNvuuZ0xWMB9aSeIyXWhvvS3l4v632pQQ87evKsSXVvyYcD+LI7cZ
DUbLDSdcUMFuQzsaWvoczCoG63+eXAdwuCZL3oyESYjhpOqK19mEV5h4007yvq16R5PSfn5TWPc3
rH9OLknfiwUyRSAr5APzkUtNyiGFxIe2sDEcamAykEmzLmowgbRxQytVbZEvSRKboN40kFUODYxz
m95AmJkE282DOiVJbbCjYVTTWHL3PrkvazVKO1Lax+vZn88gFmE5QmnFlkddpFuwbBHATevo68yk
OINvL9G0Acs2FV0L9jfeCNUEaRdVikHbWxuWy6LY16jk/nr7kyODXgIX0QXRh1N2277gpym0nCbn
/+HhL4Ag0AordEgCOhHYo/OU7/AIzotMB4e+ZP9E/5WdXSewlc3U2s6sJqH3QNspIKuoN6mmilRn
an0u7bJttFFB4/TZNT/QCYHa1mCMj+hrQI4uNS7aocbMRkZLGwSoL309StBhew4IbcQxE0B2hnD0
GhcH1PFEX+s1LDMG+aSKNMSSRadIqhv0zd9QCRqabwx4Klkm58erweqm0KrozJ/QZ7CiBmqm0eGu
/79cwIpDN+B6AC+kJWEYUkG4O8ph7nWdA3x5K18l2Gqy8loeHyucP8DVpki7k6xhv7rWFNZ61mtK
igGCI5BVBHfpupzq4L6l1dQUVzpkVAT0UWqeEA19KFu8d57CFZk4v1prgMy6btcikk7FjLualUrO
1L3BiODulkB5DCATvUn11NzpMk5IYl/ICb4edGdgnfL6mKaz3YbDknUEv2jrruIzVZ8OFsnpNmEc
71ufd9Txp6zcz6df83zHZQc4qnNCsHNUtAvyTw5ep0xUZYfedbw5ZcLAzBBeAwbyMvOhIGf3RLsY
g6rzdhQrHeQ5tDxy2huBQ0iNwmKeKuHsxmGxw9UYvwayxZ9wrQsr60ZLXf6Y4UyxY/fX8vY+n5tf
HGDPJweKVFRhh/J5iuW406lODZuzUiz5QNo7eVXXZK4nHhyB/WJMDm20RfvK4NHRTZelKxrDNGu4
biEdTGPFl2Pr16kzWN+ixbK1CTvAg9NmkgJ9uYLDgt8cDAYJ88FPOfwtBcsV2nYHD2wxjalEiUb6
BhU1yBl9z23LKphZIgH3sROVqSMZT+AQc+osGyWOhmwHV2kbLu5gCsTsoUrqGUE+w0phXOrOhRAp
tzm+mvxmm2diknpNIIhD7Z0Z3yyHpszWOZsFE0sOrWfooGQqZOED6I2UQj3O+w/1q8x3/GlKHGkm
AdKSfdZ93cMcakmH2/kvhB8msfAjhxOH2ZvkbkyuW3B1qkq5F57RqVtsYMUPWyVfOL9zWJxxqian
cUce27E1K+LyL3hzLsVbUfwB+i94jiuu+ABaO19myhpYE8aLo9EaJtJc1hQAYA7E5QIVoN++7TGy
tukano4cqnIdRMb6zl8K+i4dkhOiKInmskJz4Nscpwwh7Q/sQxQCkWRipwpILzywgV1bAOn9n6C8
cd7sVA1uPvtJiLXUeB8iICYiY7xJM7vTurIwY/JKhcWHGZ2aHPbrHHtThehVrHwiWBHCDdEOWi4V
1loJ+U3tC+lJmJUISTYfQSiLTlEL/seDfgkGUFldQXB6EtT7Pl+ukm+ArQ0hbzTijtCEPKja+WT9
CFAfwnXLG9uq9cVFWEeQIvaXBC72Ps7gBgTsRAV71Q6nhEjJMhNSol1n9/9rdUmY0X13P7/r5X+K
qpKGVzrrT7t8hATWrJWbA1DggvGMyIUKYU5MnEMhb/BTwyEfQeKHde8ha8lksupXn9NkSRq8f3lI
BL4XC8h6Ji2gHNX9gRtEs76JgD42FC/v9WwW6Ur7TNkvL8iIJNi+uoR5V4AL4vuHlIlDDEJXb8nh
t1q1thIVLW1Dzo/q/FyYgFbCZQpReKRIb3UYA7Pl109Jt30qcKvct3Ys9+FrohD7tMbdgM2UQIda
Z2enFMukIhYnOGs+Pu8hxvm0sJ8v2vKdRA6U8Vbu5tCZ+lLMVmcqh3jjB+MUFMy+CZs5xtEIizwh
XdlHYDJF0GZq1feQlKlP7eqkv7zhJJyF3Ka+kwMFBVbo1y2tYgkbKqWBTUtV1doMn6CtZ88fMDSZ
l61MTwbZSEw8wP8WUGzVYA5KdrPlJ9iOPCUTcrRTDoNuWissUSXWeE6rujUQZDSSRK6SBL0jiyUk
WY5N1yIJ4FOISw5yPdNY8Esl4lrSPzmqdjRs8HA/IhrJafER9eeP3faAX7/x2xqOQxX1fOy5Tu3S
GCimwsuIsYS91BDgjPG4cg/sswiPIAzNApvVjlE3IkRUV2obX/9aje+QrXOXcIsUKBsMC4FaBUJh
XpOaQkjEH48RbadiifuXDdBnHXpx/uSgxsElaexiyaKgEXwQ7xtL6cNro16Tq3hUDXg3VQXU7er2
PjvoNRf9drLkXnLhpSshEMvD+zLhXivdaIxFHHhlAAiPXVkwjbELzb+SS8fsfHeNjmXX7AmvMnGY
IwY/8N+0dCiPQeP6Vf5yuW9uN226kOFrY7oU02i8e/DaD7oleYvV4tvXsWanUNG2rXRoAM2w59/B
3r0CPpD7qUhORK02+V3MRDeJd2OUo7BqEnkVK8A+LDkVghPrU8wS2kbaiTE2TjAZnCYzytFfAfxe
VWpMffsPtgX1oUbI0+NktlFCDmpNzeW1loIYv9fvj0VEAFuSA/fIxSiALK7WLmY57/QCzqnQEO9p
NoeSVcwLq4s8hHOH1QASaBv+GPdvtHOuE8wzBL/TSyVitvKWO1ooTUYC5mWfLw9zw292j4Xvxq1e
5l8sfNR4n9pSHra79xl6xmE8Tw71jrvL1IOdIAWEAIi9oLjJHCxPvPqa6jG5t9N+GnqqByfZLqTw
VIlNgnHaPVdu5zA8hxbyWWxp00UjAEqo1Z8fQ+w50ZLqtr4P6LwHfZYVPeg8HtyLO2DjHvlKxroD
3u4Ri2wJQqjXvwDo3SNVt+54TyVi2tcN6V/ygcsmWlS4XaiOYaCDdO04jSJ8DFqPt+z+GfEbmbD0
ZqAVZ6wjjChNt90N4JLYNByV2KlKnF+EKzF+DmTEwhyGOHHtupoMZO4Fkjpx5nkeoVNLOSA+qTBO
4rWkPhbczOMgP8/fZuDzdSwVEyG/g+vvpe40xdTA50JQRh6iVg6ISFXSKoDCN0SEWlmsWPFAkrAA
WNHm4dX/y1EhRDXwZm6qjbznP3LzR0fac2uruCTS6lG4lndaNv0AAsd7hOgy9Qi8tn0sKPMR+Jep
t2F/PZkUec7ufEGDipIsk5c0mSPTSfqrt4Q9p1neqDE6z1MES+vLff1TYLNet1zybVk5xM5nBA2i
i0vcSR9/PzWEIH078CUbbudmkub46J+jxch1Tx4PY+dwaI5kp96PBO+pn3VOHlI6oYrpH/WwZNrT
NCYcI8yQRK8voRmD2Pn8IY2/4Si+aY6TZfpjfkuOdutyJyD17hmAke2c5S3rYS3VFuLJ+lMrqK0d
c9hw4r8v8TbWDjB5exxomEfeYrZakzZIb5+NyWH7E9NIC/xuhkwYMzWqwZ86/j3XE2n18n8I2+2B
V8qOHE857C54n7G4nZR+TJW/UmQE45z+HTad79R+Ngo8f5IujzAJad3lbHb6ZbIVq5WPP1tK6uLJ
1ksPILTKWIkd6UWDWSbZ5xcHBGVwrknvuksndVia1JzjVkkcBtXaukLd8jvmIkwjBIqsVAfiaU6s
ER29+fm7Stj3oFVq6AjAnY7hXzAwDra4UJn5b1yWtK3eDQEWbKBbE4BKfih3TIzyVTVSEpNTo6Sq
5NxPY8whflqXku4m1u8oSmzBKFVcXrH4aOskTP5AmZRwFwwTwdmF2uYggz6Udy5hqIxxfHuQmz6B
qd7slqz6zcGmeKBU4EdNwUVTH94hF8TrhhU8xwWwZGxYJr1aFrXcYDxj6Bbxh17/+a7bPpd7peSv
3BxYZc8BAFrbnumS/IyBfxcZ8lnnYn672UBMWaCyUlhn2iue6Eby7/jLD7/GQ3QGOhDqIdh/uUig
qcqtHHpi8xNXoyhIq3S5+SI6FmuZ6YmG2TMdt/DoNzFWOTfbkhkPL6zhngKxgLyQM9ANLrancCio
KvmjzsVYHmwov2I6HnO5BL5+tJXuuJHWEmlGq//hTnKfGkqasSUr+C2Jf8xCOZ3U/d6jU51QGNpr
aOG8RTQmPHwUMMf4zprMqC78tt2qAeFHkf2PtjjweQzNcAH67aOq8mz9KzaUWhbwJykwymYnhLQW
zvMTlqOeaD6oonOr+TFTEDaRlM0t/mQzJw5g4qFe3yeP5ZWbgDw/9zAvEEv81J/qYo1IitDcuHkQ
JuOEnhznWikpDwAl9RRj0RAHpm08afo+ccVnZ2bzoL4PxyGmSlMybaurTRk/CagLtfioEytjvKPI
52Mf5t2VtB2rtXcM4pO1heFnd0CLiii3slnk6q/F8GOLLNDLtH3kke7azDtc3D5Lb5zKnL4Y0CP9
IgHW4ACoJgVyShEzSRQ55Mh6mC+43k1oBtCXo6zlxd5VpbGeuqmrYPiAiPlFpo3wRTs2JygJT0nY
yojptScG/BFe5X3/lsYnibp+QdiYr1NskDQgU7jjNJB/gtpHl+5Vs0WhQukaJn1iHQr/o/FVIIIl
rROyOBal1kbIvzbCELwNlvgmJVvo0tvQL+5AhOPwC2VPpidA+vX+4AthpXObaKX7jSJmnFvtd5KS
He0OFSw1Atd5op7XOY1G1390CF2b3D0/ISb8SBFElkL53hUxojnwXDj0UMBVGnx9EtwZGmryl9RW
SUVZvDUzKDYb2RS/e8NPxEPrsM2ScsBlyTKu3EHtKMKMYX7jXzxKjgIUQSihUVM3r9H/FOUvlbri
p38crPPBF+2iGJgToBBuYZ/pHkZQmlE2rXct99gRKGnTKSnS81+DV9E3EEhYCw0Osu9RLAd6L54G
khixpYP1D7Aq7Hod8ScKKdfh6nxNVh4KHIFocBEYq/91eU6pEPKo6Gq6nH/tEkz3RwlBX1xOcKf+
+avXeinb8qiGb8j9HdqhNf4IuIoxGR5oia+//JhFoLJpb7lm3GdjeeMNvrssQyeDQZPfZhgAmYWd
dNDL8B9q1fw3Z8fiWJPFwvQIK1EqcS6pF+6kNV1ifeGt/atYCWwqov1crAKeaX3nPntTvVx/HM33
gqF0XPBXCQq1wjq1IPJNd1Xm961r4m/X/lBhSKlVoDB9WNJ02syscyuwJgwmShxYqnQ536NoMSjN
gYkehMT9bgo7kPED7FGsKn7Qx//mj/YQ41NBaf5fcsvLhgU/k3ZyRieW984GjmxbAkZjsCPjJjwm
8f5HHjHkLZcuJSzoioHFipIO+aLZW3ve2PmX056Omxqf/wG+CEYSs0nnX+iXO2QdgNf90Rm1VwCM
7n2xwBd2gLdV3Yug2BZDWMu2tt5Mw/z5kV1xU5opM6DwSCjjnTmb+GaxDIiVnmwTJ1e9KbJq6K2k
ekBFh+PAuzvS69V17gEcfisUWIzvjEkzRmWSTDF4aidyG4AFQbkAfUdhGiQaDP3iVqat8o0oWbv/
gW9+sjuy0Hcrsm4SlOcyDuMTjg22cjSCBOQRdNJ3wRY/He5f4i7wro/lEIvZ/0wkp9p5kv9HxVUJ
LUrNf6fUUdUDzNyc9I50+QmT+IGy98Dz8fJCrhc/CEl44QIhkzSeimCUxYttdKiARS1uUf9Ad6TW
QGccIX6AfyXW89Kds60BOTex3cAaFVlK3I/ca7iMW7uNKXAKa7E4o8jVgwHhRtYWNr9sDky0xaG4
fdho5maB2aQ+3yOzaw5uBVtuCDfg/2+OZ/H5x3r1TBubsqEf9jXP+s4jffa0YtgCKiWrIjgoSguK
er4+oQvAwrplyK6mtM03VTdgDyqSRSSXHWzO8GCkMko/CzqRLIZZ0UE3mBnBJZP5FuSSoBKAjKKl
bP3XNuAHUGzTPuf2W6CC+xJPngYTxuONgutKAfS2lOA6zq2Fr1dIQU4TZXrbgLbailnbYJ8j6uWq
DZd0NmH4CtDspXBVsybkHmuoYlRjI39R0jHI1wt7U7ieuTsy1DWi7IVAk5GdO2/aFEXBX3WrAzlk
plswSVGcyHfRz81s52YGsNiZUwpx6zsqVdXaqeVk3o6s4Cp8+UbKVuz6NaqXKZGGsB5EqgJPuouj
WS9DnohX8607XetVquf7QkBV7V2euTtSwhGR/PIV2ZXAXZGIm3w12y0bxkrI84kmoXbPSf7td39f
MD1u/MNssNKqRE1pYt4z6CRj8vcKQ9Oeyybh1XvjzHy4KLdUN/+/ZpcBSqu69voTX9yCRdUVUQHm
AHZZfGfdSOmHLQ7Q9AshLJwlo1vOpa2wsJcfJyt1M2MQ/qOFwdG7nmhhG8OwkmEnDFgoRF1PkWja
I5BCrekEkTX6I61tAvmclvkoQ89Hj2ErCdTtSuGHKIaWZiW1IuXzBZenGwMHXf0RGS1UPNJMKQtH
1tYFLalhcaxdGgkZ2WDXTiUKMqBbK0XYEiiNFcbANwKpC9gPXixzwNnXscvP77o4cASXzNMi7J59
eEijzGm8NMTU7Vz4z3gwTy3R41SVJrdLrLoMRnLmRGjH9V0Y6/lrpqFP8gggCZ1Par667toaNBIA
ys+LluVx9aM7u1++s/vavNlTScBFaP6m7oPcv+Ry7XdjhTwlDo6qdFWT8J4RB5LON+g+TqVhqkov
MkBl37M3F6RnEOJi4LmAPb+mZMi4ufiC7hcgdla4WYJQCTK5AC2NHjVIeLj1X2ln9sLOYNypChTx
3EP4wtUXqcJdrW/DoiRVi5nhv6+Tz2Qr1SdMcWta9uqzSgMyW5sypP00e8cLUb/J60SM17PyfsQz
DhNAqB/yqmpP92CiOWof22rdAFMaSpVbNffXN6Lvmu6snufSmLhzytFHZPEhYgfTVApysg2hsIWz
Bvm/j3iU9EBppJokDWF+V36Ig9Op7Dsq0WGQy8aSXyPbJOHYJuGhHXW6aXnmzmSXxywTnNHR8Wwu
9AqLIsGKwgz0gn7PbNpPDBqfhYhhUmiFFYT7R7fz03z52in3mT56Gc15ap3DY6IYLQxNwxRW975L
VnlzAaMA/8vS+UwEV64dnZfKn5CJFrYNeNgou5tbeT0SS9DfPSGl2SmwN2/x5rlBGPj0T4BgSm9q
WirRP7L+U+oy0ekc2eGXFMTML6dWTbXeK2XCgJn/Ccv/jDoruxqjfYtAg5gi8nJ+nxDneZ090Y8Y
aujAGlqTEEvx/p/AfkiLhKiHe1kT/crsc1l2YlG1SQsf5lmlQvlK1J6P21ZbL9mKO1FivNYHVMnP
PXuixaU7NWm5BoquZTOhZ7Wn/7Mkt0+LSvYd6EDpWj0UkGiK26ZuWDCj2dDfM4GZsxBwwmQ596fk
DEfKr749ptB3J+EbPPkF274FBwKfkpYINuJmdYz4C7Az36Af9VorASzaJuv8PqmoVn/JaC4aEJ7Z
imqasdgQAAFFP+LLBrdaH/hF6LXjIdG5RitW6VVMBa79i3i4EK4E66kGTiubE6Ct3CtbfUTIG3A0
2mQvpw7t4/uBqeT+BTisy9nwFoiR6+V56I/l2RRjKWd/u1nYvHIxJ1jjm0k5a/tx1fTc3rznZfaT
8/v+fDM5NubwXqnaDANf5GHGrJc1Trrcr5A2cByhS4NNz2iutldFoIVtdJWjgkDmF1/3upy7qYSl
Vv14Ki/Z1qfNKKIM02b+ssKnC9hyR8t+DHFPfV0Et9tSVxIwMA+DW5+vJxDhnrHClYR64/UuZ8Nc
EJNz46e1lBbUoCbdn5bOZGXmRHvhPwOTM+SSdPG0s3VhhjqBWo2PLbiWYPgpimol4EWd8gs/PGQB
Fh4//lRXCwM1RZNFl3UODt1aqZvfmzaIdF+csucszxOQ471GG5NpZ2CZlmw/le2kuL+0i/cy7ZvM
ob1AIvDfPQ2ym+S7HsLN07PG1Fia+pYLjKX4rHOaASHNUms0vHSTkDWFj70IIjHAMGT7C9INLpKT
kLYKPD9BjfyhttNNmg3xOf/Tki0xcSeuqdjQ1E/UQOzsgnFTzu7rJh6GrCcqi959DcGvqaSR4Rat
SbgktnHw6gC5H47CcEe11il84ws1UZYKlk6lbD7F1LdhwEDECuXVJ5jwl/8ASddR9qlZtg7+w4/C
jnmXV7fluRS/P25O1jrR0xaxcm+CLuGpSDVR63ENktZCw2bmnlAgqepsy+qyUFDq9yZVvcNu507B
JoJfuvoCUkjgKJmdQttAF2H3le3/7ct+3cF0Vo5iOK+EOnBPh9COTjvxt9yPFEGsIgkens7k9W0W
FWFtPAaO4aSzZk4gvl3WEXeSum1U1iJFiGxfv3AT6Ujrzt5IAW4jBM4r+1MXQoRruXB1SSW5n4/u
f3qcFbERrpMqCANMnZz3xl5td3TYBouVoGUcv2UT3Efd1Oq685SBufHO1RooCrE6itWig6xfzCTv
yNABD/sNNg4o/S4Tyz5qOlcjC3WAomNuUCdLrLQdwRXfI7LpTTJzn5iYKt7a59iErMZMpDjfohFW
68AbpddT4oxndFtaamjMb4NB/61Iqo+HQBitYwaLExMIFYVjJ6pnGQ0Z0VXQiCMhBW/+ZlujYUmi
yMxG1J8i10SqlURsLRFS9+RNjg9GYWtef8FcPFcGW79pywqx1HAzCkEIL4bi30UYh5FIWT6Zitm5
0EiuEAYEDnoWdL+MVYmqQrgKGtjgdFrszGaQow0x8oNsM3LNpUsAhELLcc51raucyPyTLQT4zYD+
zfl11ZbnNt7kwYQ3UtVPD6mKv6+6FLtlEuesCXj0n7oLSsh48PngWgkhAhQjB/UxaxPut8P2PjUD
k6n0g6YJxvPOU4Wop6r8aOFDic+EpqKQnhQjgk3/GPFlQHVsqE84W7jRMDZE5sNqZGGk/tCweMUi
XUjDSin10ffCZWuM+KZfdAf075o452FcKQcAZpOlrJu2HPHkNyoZQ4D1881AOavTxWsjzM3SrEKO
muNCvidmSzHea66biMiCWQwB29Obkh3DE+vmHZw1QpCwBWcu+qdZvAfsYtQPWClkRLuo2joMYBTO
kfJIwhdFDNGR1XhEnNAqZwYr+LSaqIXcYAtwpRInMca4AFp3v6mGCHmUR74GWP0gS4yl9Skqas/Z
cdaYWzRaPISPyA8a1d3nshUWbw5w1D+DTl1YFLittt693NXQ2jCjYcrVdNn+9jsBBUzDeoi+cKrk
2nR9xrx4gq8rqO12Wny1Eg4HPXsD/GnAfjKsJj3WJBjB6JmVIxD3i3IjREw9edRzl5EWxiZVf89Q
WJyLa3/bJAttC6pDj7seMPwNVMwO5qrHSGMY6WNtvAeYZJZjyyVFfGWchDZSoBdZSO/Y7WntfQgj
zYSPIjrcNUCFivmF9FZWBofzzJLs8Sz6hzyJq9FT8eav5g7R0pjIdijcQCOTij4xXbZuRa9rsmAh
76GEiUwH3k5zXaHlZYQnVThSv28ZbMKG7icpj0PIHAw/0XCiucy0/RJ5wjXbTMnsD338mEXpI7A5
djot896lvDITIktvhWsO9OBCf7rW7RuKPtqKszHP6AXkgcqMOGH0lSfBR/6N/0pOQqX8lccGaxBf
stfkTRdrgVCKSreWbYq8fPKw0O7YxFZF/YYmvr8cq+EGwmOQWsGZ/TciXlYUnkMnmnztssyTGPhx
D2w6lcD/aIQ5z879eiof19/6NQ9K2+59VnBx7JDg+fDkSgn87qPpEHuPf9Z/smXz2qKmoV6c0675
0r86UVtVruid0SUfvJtZGm5EEzwzPN79oL7xtpMKF3xLu7QLwl/Q8bCYOWOlfYmF7WMfsAmT4aD3
jmMD7ETLf+TPKz0eHlFUP6UfR9utlSYLdL+XbVcWzFeM3LDOQiQIslLAbNkWEdOCAqOhXwN5nClX
8oCqqaWtNF2DZ8qx3624R0lB9RnJ5w//CuG2gWzQfN8hCJdjnQHhKZ3RiNCc8ofZO3UwUar9WD7p
MsT0mJW7Yv8eXaUz9kuoMHqBMbWAknIgkGXuwzJPHtvRDkfAu7AlaDfsItUfKAh6q29Uv8mkdeaL
vBLCK8fVIC2220GNxf0O7vXV1Zj2QQkkfKz/bt0Nvgm0qoEaU0XJrcgX6lKy2rCRURtC5uc/N0nn
zd1hTnsuptlgLsxcoDhIUmjIo2xHP3cQbDB8jDZstLC+cQ8nc9qsTmfOfoppojOyvqHPMLlgckIB
cuAHuztJ3dx1qUL/D2NIm1Xwfw3u0COCh8jnvRAJVwY/60BHq2uor3L2On+YEGgpSUsL1+7r+R6G
FhaS9w7Oel1DBw4neYWleiaXzxP81d8eOLh5ewHFdeR2/RTzVTR9sY4FMDetCnB1FxxXluIamHCV
t3VlpABQu6ZRT4ZXRqWjmLgDQ0bcsIFa82LsqvVoLb6Nv39YTLZmMz1l7alenwQ3ZEZsowH2SBJO
Mb+s5Qs15T8AH6LY207rbtbtdx67rdSLfzLvZHUTX5ZhRJs9eRzD6cdmVXZPbcklHDmmBJlQFyjq
G9zjqrDv1lrSs4EVYxAw0l3LzVqJPr8yLQHHmb+5GkzIkkztvwuaPgIddBe7SzK4IcBBQjCnnkcG
qTH9RUn99OHGnD9MopDLIanXVhr4Q1rUHJJsXahwm+11fvFyOcUwU9jdG9/TSF4AiZdOP/K9wBIF
mC0PxGKYT2PY9TQf/YJDW5H8iUn2QRdM5eeytGMPpfUl/VXjoGB16EJ3Deh4U3YFr7hMoXmw4I9m
WuH8Tyl2ZYBntzbYkKd7XpXepOai2ADjrH7fKJsOgzzS86AyKanELvfWaumHvfw/GEEEYCQa26TS
FT4+3V5X9xie0+HTJWMdcelLnTIy6iq+HTzppJFrMyV7hEQboKVuWVXHsbE9m41lAuYyKrWTQc4v
liTFsD4Hhw7UGDATbQHvHPcTYO3r7NMtKiXn6+eVs+kCCavgWYRcy+kTRlebmk7aWfCqjckiqjot
/zv9Uyi1rEOB5m/ubtQ6YTuMQreRW7cvAbxGBSjmPVi6qPnN/HMrMDGP//SN56wURgH9OuvKIOrK
B1MASOJzF3oWVX1j8TEIJs/7lwMe/ry7Ak1yZ5X9W91C+wZdePyW7+Xu+uFgEwbSX4fJODnV40fF
FzXQqryA3d5dhB1M2KaZiLm41XTgKIVLZZ7JZIlwlcZZ8iRzjjuie6KDmjk9iT8s86x8jAQcdbKT
fl81t9oj4lMYja56ffvUOq8y1ggrbnsmxsoh6qhfQy5Q0lMY3dCbPmBq8edLoSpfzQK1qC9lLzqA
MKRRuF9/PfEAw3LnsXBEaJkF085vL+u1tUEteArUFh+MDGjnirBH0RgXiE8KOuGJ+cylc3W22bv4
N60EULv9l+YXJ1RrGpTMUm+GqyFPr2GGvyf1iSbKFeE1248fw4ygjQC6Eo8+g63oPuu9onVs6Z7m
FY6oN4EuawTLpK/1JBFKKMTi9QSJId6l//10Cu78GHv69SV8nZYCzfAwIwVf9Oc/nFsBd3UIwfI8
OltIr9BVps5Or16pUBrVnBuI17r7bOTYlYSAufhn+DLGNvh0YWcHK/OeywaKZPDxV6EejcxKQTpJ
oB+cmdEOEo3cQBcBtgrjrJmPNHGGcmF4de5NB80CsGZI6nhbBNJMAwKKUp98Knpex6q3R5m+RPPz
KSbiaZZvKdmR1M22tYcMJzqr/cFqi3QC1ggeU7zmp9YfyHjQmQECInmgbcY/o//qyFSc4rEPIjsV
L5gHBSPKkGRv9fTSrWv3k0K++fn8oBEYIEsl6NM5bZQyzP+KK1wTpk67Rw5OnRNMTBpUaZ0wk4HG
NZ0dr+3eb8EWypplgTKb+gnplLXsMko6gnTM3qb1VLrbdtCWrpgjxpV55iB7Ud9sKa47iUoFWagl
oVcBWJiH3vVxEim5YikankdZ2BljcyDiSQ1wLWI+SpJZ2q0AeacLnvm8vWfrX7NuTGiPYYnhUkrJ
Fo+aOFLDOoen1eLBVKujVpiRzxbZsEBHJe+F6LpqTzJWZqTnQJaBAR/LwSPkdaTGdRYIlCDeHMWo
9oSM47wvG9MUeSr7/uKMl5dBiQmxtT5V8UQqra+MfvDmKguJ0cf3UFIxjM/0KeDLm1Ar5NnZepoS
M34BfPhkDBBI/tQUroDQj2yyPz7Dj1I4Z3njiwsz+UpbZurYfjzaKAEvzCUu+KTOIDoTLGt3Kvgq
lY7i4wA2AYcnkvepOGAEfEVQTYbsv0P35O09jIkZrExb5KDzACETHdKn/KrQ0nCbRQhg6bNjOtGn
K38VAUdMyZeDcAkT1EHTnKlo75/sj+4om0rnz857WxG4Dk/JbQKZPLO4ZyPKWiNI3p7cvZrmD4y3
tewqt+Tc1ukk+ugVkT8PcgW97Xm9VD5oxQpSUcPlUkjl0aejRYToShBOnmJNi0NyCyQxUwYwaqY+
vYgu9uMpCfdy/ueLZqpzR2z2iL9l+TRkhomFCYdH58XAgmEYkPezoWIGxR7S3cGqZ6f/e7yX/H8V
pc3/IwcGXxREFu11YGE0JKFCiJQBlvsZ3KmUO6YWIbDWTOpix3pTMWYze/C5L1W1l3X/B9fiSbll
bFJoBUs0c7ppMkEmR7djFSM7/7QYmavrTglIN09yOOet58ct0y81aOlZrHHKL7a1+wAzz58OYw63
27SPg5i6MQ8FcKBopAkISW7RSp2zT4yxp7RVF0k8RwVpIoNK62R1aB+ayjDWbDaMdymRCHys+rr6
UlLV6zNHAeADVjtjKZ+zbJ8ezNmuezgWRK4HvN7h+3ZcYRzb+63GDrBX2dg4/H1st03ltPbF1sH4
QlJq0Uu+qcGDUljqjDnjTUC+k0hZbrvbKlPNTj/nvn9LfOowIJBo7JzhOh/D7M9X61Av0BiAlsqq
P1x5Z8bQ2mZWGINrm40EAi0k7IBzzyYeT50ee31g+odZ0ZS6tIfXbk7d5BVVd/JlW9T0LGGfQ5ZD
XLPrlDKqV6ox52ihGrMAC+JGNWvQPK1lkh/CwEo1j8v1voTW/8VrkeMN7wrZJEQzfYr/yZJXxyha
k1W6ncU0Q/mf7lt4XHduqHNSFCkHtuFkkRelvo7NKiBaAf17Lrp8hNChcNnvpvJ3SB7rNJKbgfr2
i3HcRhQljqOVNI4hNc1ladxHG41m/OCsfzOEEM12J2Fa/JcFdSS4ruq6RMbwJr/uPnWg1Fbud1ua
bVwqSdhKmteNpBDIQWWngKrUcGT8h894MZplkE8J25mxb8+3vyZcx8DYc9icsyNpkSpaWJsFd6vk
pN6iJLYTNKbqoaJVxK8ZFHc8S0tU8vxGLUNPq6R7g/lDcTLZ8BAFY/XDGd2Q9O39hoab/RTA0f3e
D2hEWV6OhuruwEfTca1sqn/Fr0odDAG4NS4C5YecJbymD4GNL5H3WMUtf+F+XCxeGUP6d3Bjrjvr
7mtTvV1O0fmCpneKZhV45i4GpNseyTPCUAc5gFTgRooSYihuoNDmgygJlHAvi5fge1kw4ZBNGXmH
tn0mk2CbRLScnSbzvID3As5FpuXXEXOggTKzuoabnIIH5GD26JT0IX+ze05gLuNw6vlmZSv6hIOY
fQd3U8g+30+veaiJUq2kdl/zniDh5EL7GzIKK23Xp8cEcCzYm0ZHWO0QDA+4eBK3Zxk/RJ8LlzB8
+uFLbZgdPyuMuTSM6r/lR+pJTJxc/QcLWCldpJFFmYxgMTMYnTezW0VwjuzJgznPnlICPV8yt66i
gP9MY+yBTJJrM+f++r6ck1mflpHSF90m5kP9+1JJMJuXkGUE2YnioSaFTo2LE2e8SCkvL7+YyBw/
ZbD2NQI3EfMr81CZgAw8keDRSydzZ5KjcHF4kmP4vr50s4uQ6Ri7DvzLeYNIFzZ4Wd/EVvxKXVBn
jxS0DXqNcZjdCFEUCVdF6rqxraZrluTJar6GlTEgJYj4WPHuDjZUftMaEjZfsVud6V06VphwM0C6
BhGGdiH16Os+gMQh2jsgIRiAI67baR1fBATnJAgtR6uUdC5ZL+A8lwY0SfG189ObfO4aj8uJbW+/
uqIl5TjDPB+NiMmmtkBkK52uHkxFkjbTaprK3OYnkdRJCXOmH0K5RFrK/ZdpNimqcWAVrvcNUNgA
mGtnuQi0aFOTLXuwWEVZm4ufKWzkcaOJ47iSzVHjGzl4I4cirL0q1HdBlv2uOYVJYAkLhITdYlm7
OeDGWqFf+FITgBLThEdsVPHgihkHpb1WubGj+9U3cRLQbEYoMvNfV9F8Jp2AR7M1sVNBUlN0V7Ub
GZM9Og+klvKYohckKCNL67UnWM9KjBTCpfyjtxXXJgU/7KrfzF2DC04XoP8G4Fgj/UrhP5gCiCOu
FBlUMkk1glUGBR7FZSy/oGF0UK0gk/fOyiRPGgKMycRAG9PNNmPw9XW0i7QzV4nGWZfEuK5WEu3C
0YRC/tOxDQvmeGR8e7jL00+2EG9Uq5ofN5/0cKMtKbFYKmJLmD22L4Qd+6KP3IqFGDU64EU7fjQG
RVpItfY39iwe2WBe3G6hnKJrToUT+g0Qj+60lvJW3a1Y72a2u3xkYmr6bFiz0hwk/ag3WpKc7kfi
qJuGPQ7FyxmeLU3sbUMeOFPbChQI/ccYDGyKaY7di4CaLlnYDTA47wr1616NNWTuWnyPml21FoMC
GIL8vEJ9ykdGajA/GPfTjqcGhblQZ+TLRYlQBZY4mAHvwk+L55mP6mmvQg3vKsio2urpwl4RT6LI
+QPC2sJzuiiBBO1XUgcnna0A6/uUnpLt9dEi4lCjShWdwlYSl/kGqYTcl31hzn394DUXDKSa8lAj
TuX0dXdpCUrvmrB7PmK+wUKm8kgaDizYFoTna8IzE78E+u9b/E8vdhmas8RNebwEAorqWarmbr/2
Xd4uTcvLl6syumkRCjDzzqQKp3f4/1+7QfUcs/jwM+a5APNc7qoVkDLD+jIBuzLrbbNVVpIh97Co
zO77fPZbKuIYv9ClRuvwsl3YEeUCLOEPABZD7FJu8bLNA6k8ZF3LIgouF84WXds7UeFEvv3gERif
gn3/Kl+RfUSyAdutWS60D/JEtelSa4N8sE4GPSZF2oOGXCtQjSxZf8MUjChnz1NAL6nFOxMUFtn/
XUPnXoP0dwquqsc5W38E6FMYGob/GNMgpq16ui8JE9mbjkDrmXmnn/7oEEDT/htu7DOqyr+AIn2Y
TnTvJ3zogdxsmGOL8iTPlp6JPu75CdvTvrtgkWTIpaQg0ZssNqb7pic9JXtqCT8i4oR/UqcgEitU
IaevK4DPpFJNTk3syrSkvHGZxDmvuWfUpcA5TBMU9OJ3EOIaAatAZNQoxn3kSt7SIO9sURqiL/4p
SVGT4ytDu0NPVSuyatyxOD0kUcqD6UlFJzwT+cVgukD+Cpj/P9gvzm99KQvEo15l/SjzD+3SdAvt
93mKI4fH1znpCqNGbjia1YjMslCwUl/sH+eHHF9/hM/MkudPtHXu4B31tDKimKNBfygBnJpUT4P4
y23m5+XdpXm+PVpEfVdUpKo7iQxiPyLfZ3BQ3gyHO84E8dXrGxStUxQF2BYS3EmZXQfjig6pezGU
d2O9p3pa5Etf/Pu6F6hZMsRG35TG7LhuIr3QMahA56KMRdPZZeJqkYr+ps5I7m977DQYTBSdB0hA
0IIKUXcurrguNcLQ+YXRVDJbpsSF1XOwO+3FC8NqPIL/2txCsyE9a0eDWehYDNVlLJQRh42L2IOk
/fK+y8pGJdDFVk7thMZluxvF/cnC9OYUsVIqyVOvxDEYU5nnc8qsUrY5HYkcDAh8RN0M33q5QFQR
MDkXWStsPugLGWbzZOxoNSQpnnJVB9JpsVovE/teyc+CGEWzJpqNuBwTGzLjA/wuqWvBnhBv+aK8
CMnL0QMpS+7iAR2Qf3MNIzcI5eTZkPXPrDsBr6A6oieydj7ukx202D7+m8jdisULVqDYyRjrihgT
FCtCn+u2luQKGfyDvXHbPjI1E5lF+g7XpSfoeBmFl7Ib0i4djTF/nUZwMtgb0Fuc9ookFQJYEGLE
paP+9bhrcQxGtp4q2GSxxUDtqy7WfpyxMn93WgQi6rj3X+fR5IuOJ2kSZ6c/0BJola4YhTLZ9HXc
frZjgABknzzymgHWTQCphiffMxp9WWPbNQDeI4sYtfpb8jsMaa+cRdtQGrNgcPkh/eSeTjWIvlEY
iuQrOOIzKFt9JdAhDy/+KQzKaj+gp+BH/oqoX2FJzRpnCrY6R6/U9TUR2xToDrbMfO9j0FxnsrUI
FB8GSj+MP5lLPFBHSaB9zrqR2/Y+oxf0EfsFsp+7VUIi0kw8AjxGsBJ+pWL3rOo1pxmXBbyEddwc
z2neLZOORBF9gIBcteHOJ+AEiKWAEwnSRK2Dw2cAbopwiwErhcjW0FmSinAcuUCT5l22xOebfUyP
2ogjLtWAyagXU/I39mLMkmvR7xlWbLs2ZTNcAAtoOI7m3J1PsRxWvuHXjqmSzkXrBiY3mCwfy/1Q
+raM8J29LIDEtunII3QeDbc2INX4vd7ZIJp1DLtV1Psz9N5fh81woyXWHfEt0ddKCdP2Ylk9M5n8
1pB7SK18s6PuO+FI7hjGUHjxjmQ8K3pQklxrf/l1Enh+w6nTxe2sR0rh1qFIf+4n+0etTSbivLZQ
nm8qQJJ/AjVZfMoUMY1tgqkCMovuoyX8Fy8thqUq3RN7n3sAYOrMXc9N7npYMptLpXPzaHBqrz5g
m1XIMA4vOn2I/McO+FXDcjvpyNYteTRPZ94/QdKVyPJL4i/EvNYLNC9DGxxU0vvkNsiP4iLUanhu
5BRbsCUXE3YIQbEgwHX9wEWkADsRFEjRQi/zK1PuwEuLAIRiYeMdf/muUKtPm+7C1sjwZDOhXljL
/MoMVzZcSrC57e47mEhhzV0VeYinftjwEx6tFMtEdyFfNepNdxH4KAnvix0jXKlykhYzLN30Z4yj
DhMWOcmajp5X3J7b5zCNI2jbvp4iOxlowErZrWzl1kkjS5GxBbnBG/KZ+WSGjC21uND//VNPiPXi
blP7+pMryhXqT4CCPvUwu7ZsVluU/C17fVuWxEY6j4gkY9sIH6gBEozHxvvTPgTtJh7nVMqaMRr5
Sne1dx/WWFP6lZiH6s4B+NEyHhnBnHjcVnxoeCVaxj06Rru8IDhWldtmAd7NcRXzphYSO6/IIN0h
NDrnRfgQmTQVUCRQnoqLV7H+G8gcRfvRkhWDbi7i3D0hw5qpxT4XmSf1GCtNIO43AK8gCWjtw7s1
Alp6NUj6bdPQRdbEDgYrlPAQ1wmS2oQH1TNHvLRES2e47b1lvi/C1cK9HfB4cQR9KD1jPyllKgIr
rFVx5wLXZzeLEyN8WqDzbN58vXgHO0EjsfNOrdgQOh3+B9cFBnd10ysR/FaYH+lhjEUtss0OaYUc
CaQMhZEvqPy5mIjMtiNyYsRl1QFR9sUS7w8P7BEb7pULssM4RTnnA7QDTrgon/aPkVnM9vn+z5+J
2vbCPlcSR4lrL/SpNpwqzY7ykHoeZTbrzGVmwmRh1UEZYOVcvcViugETkBDXkvQri3ZWXAY7F7Rf
wS+wNPHI68c4KSg1yUTZWU+q2gIKpu2kO6aDx26M0O1SLReSk577fm5hq6FSUnam2ASBx7AeE+tq
S+wK4KRFwS4F5L5Vr4rJm8aKx4rrUo9XPPEQCezSfx45ScixUW314hBWKL7Jt8LraPc0C4kFt3kK
iHc+RKXMUPJUTGnprHSOXDpyGjv1icun9MuLQfVMwxKN9Ociuw8tZcHXHRN3jpdtChiDELLXRmNc
a1EU0rnvUvr641T234fDb59F1L8RgR0YqIQk5GO8I/A31d5yz9lGfoy6pV4RVaBX7Xpfkof7MKr/
KiNtxMIxeLvhEngcLJSX94MWKSukKs9tOQW4bCuqPEdxLw/6yJ+NdDYwQQhllzP1lh6rcVSXu8PE
Gi8Tfwj+KQa0Vhpgs8nVOaFuI/53/sb5j/bgZj2TStzLICVWHDTAV0JtWlyyCtSMQg6CXgjR+Xsn
0F1neuBkYXwCIzNK0dDDR3WvP5HfAfZQpUZy5nShhc6dZ3psAY/k4PXrlnsvXcPnGmdJumfglknG
KtquvY2ZtZ8plv8Uv4eu7PqbaMGAFJnmzHVUUm93DlFRO+dyK/g9gFjiMAzhSL38EOEAu5NEkl7I
n2vpK0evUAsSOc2Nt4oRXG6bI22XAW1FHIbpizLNHT+FExYYK7dGixkIQwUHP+9C6c2sVPk21Ckc
6mp5K9+IER5bYoVayZ7CQPlmBN94ovRD4awDCQRpoaKarGgxOxAailXY4+aSjUh20zMo0hDoEIYt
44wXrE4eWvvY+HM2WT+YgcHkRoTSAGywyWdDgAKUbIdU4z2b+lZm7aAjvCvUFno1LuHAhf8IuWp3
M4sKnxWDODCxxk636vNcFtxLZgELJizHQThP9RVtdaMFE12WYFyL8FdOs+o9vkhuQSGKu5edCexq
tMyL4pmd3yymnKMJrhAwFW3IOz4NyI7TjEieDehdxnqLQXWmPHBU1EvQ98ndAFXx1LRZ0E1u744H
Lxcrm4Z+kdeF20qhpKnAQWk3JTKrCsojQYYsfRulnh0DbLP9rXukd6xQflhmvaLo29osLrq5yQND
zfyETriASc2wKazo1t7EwRCWSv5dkvGofPE4rSpojxYJWVSzQ+wfrqizmTTNcQfAEyCJt/Js6bF3
m8wXgduATIrzzMut22HWPOO0fiKi6GxwljX6yxtB/fnpLXZwAeRidzmOtek8wVUdGMBFXhq46vDm
+2FgIz6O4ykv9mElsNr4i0ZK807X6c5dcQMq+4f13Z2DIck1i76V4i0I6ETUhvYi3Jt4RrUK6v5Z
LV/UMqexF9Flem8fzx7okWtBL8t15ke9/+xa/UdE67KoCZ6UM69p/8tQ8CjIY2dYjcqB/RK0lez9
qi/KUJxz9lhOHCam3f2LGbqi3YFuSW0obXxBLzmfoxKTz7DnT/0GSi24mmHJ1LXPQgRzgGjwjQNt
E2wFOc+yy4cPTaxaoOQu6kSk+As4yWl5U9fQF5M2Wan4sraGvZ2iQhbRkjXhF7fl8r4RVPaBCWq9
VNV684oGUCwhyIGW4iJuhsEcbqwF6Fh0ZlSKUKMC6+zWtbCIZ0eWelgfBhqH9gFI1U9mVODikJ8W
R5NLBQtIaNIONJ0A8jgg/XuCr5iY82XPsujIkmcHJ2Z2JocTXmFXGFwXFa8I93GPRjzWNwPJWBYh
DanHjU4QL0U7iAnTRQyzJPPeFBDaFcYxfNAtkRHHKHn3W4MzECwRK9im5wJOGiDfoCg9ILNc7F72
7IIZKydCGEXviNc0ECsMQivNbq5YxAfDDZt00l5d54RUYHZSeot/R+O4WYh4zYYrtXfEti2/0pDb
HC0FVn0e/p0c9JLRbVuW8shq+w0hxpb6M6WUEC2KD9Bk00w3aL5YKuZIxNNTZrCvEDxHXrChNwI5
mZyu12KET03h3eKlD58JgfXKXNVeKgoo5cVFdI9L1q7+Xe5gDyLbkUGI/7C+RVoFOy3wwxZDGLLa
CSQ8c+5MHoO2PFIa6+cUc+xZ/KzQrt1lW8QFFaNAlz3frOTMvOfFLjm7VAyoCo6VJWBqvAIr7KrJ
p6W1Bc+DDoPJ1XCFGDqF8Q88CXbNxyOIwcULQ5/MPoHBTDrBurNcxJgqVH6nO9ffwU7ppMouRgRD
14IVLaQRbGoJJY2exs+VSIQeSOQf88bHsDiTVYBew07cJEs6O9bhgYc8vENWWYaF2UNUI7zZ+DJz
kMhUStQiPVy2xeUc/9YxKpYIbIcwoS4eERQkEBRILpm4LbtpgzVvOtUQoz7Zrv92dM0FCuhhIKLX
4OEbC1sY7Y2E12j01k22LiSOtCrFIq3L7GHjGdBrs/aWWbF+SpS1St8XQd9eFj+8I5Ogd+RQX8XH
F7lg2/rAnsTMEjqG1KK/NxUgAhbKo83utYshWm7ObNOicAJhUqva4Pba3xyoPVEwTRKHjlvecSRD
fbn+OyDVr4/Z2BH1nAuGuHEobDUkH1rJouLSVWqAdGaJ0I9dyNChvawKcT2rCMOLZXwb6dDYJmRf
/hKKPsfSCEZ5kglN17OPYezo2n/FBNXSTQ54UArZr/LmFPijfH7Bun/QZKDZrdNVZAGuPPAaS3Xi
wsIrtVRjKCTAiysmva2rip5u9y5eYc66nl1ufJb9E3lYYcjw3dMslaklxe1TaFDmJDecMUBIxbU4
SIJGwyHTzrLP4v7SJflYWARD3QxOlxM8jY5WI1FK77yjdPm9ZmQNCGK07E6jsukkl3O3M+Oh3PPS
c1VlNJXn/rSAHg9H9qz9vRCLRVIA/bNwEDPmORQzh8fME8lS5h2jRY99zGJWmkPXuCXTUb1AtiP1
9vbOybk2KHnRZKtwestA6i8Syz+qziQaYBbfx280bkj2AC/t8iaGEXc9Ou+FRMuGSw4e9R/BXKnN
YN++xSFBbZszM6C1Kl8QOLxQH6uoCoXDsDfISS+mwcqyxz9K2psPlJeftTRVNhopFQPu6txUMqCk
t4FK/9mWkPswysON2nBuWTpO3PwV8ZfefuXpRTrIGo8/r78leipwvkAQLtMc6otMcpFzQPB01ljK
bm7Mi40ChHkDqMD/UrfP18+iMBWLKK9oZkIwq3ZWC9lyGvYa7trhtTbjEY2IWECpiC/pzns9lSMY
SLh17jGZvBvkwBuQg0Ea5a46ngD+AQN2lHVl0pqviapJ1KY7/06fYQIMiwVGLl7nRDvxUeG2KuRw
WMrz4kHm7r2dGjC9DSZwg1bkRV9VloY2brUjQtSycGi1B+C9dUe9cSYgI4daGvZZH8wiVoTqqIGY
Fonap2O5v30xozlMY8v4RQjm7HRERSMeQnpDt6qr6lqG+xXx4D6HNfoGUsp0lZNy0Kozq4dSXnz1
KegMk7kvo95E8lJ0AnptCkF9zI/Mxhg7zyzXnmbIE1ZPqLsFopPdF5GhxsZ3FP6q2kbkUaAVydnb
d01SEhd7XcBoidGeIC8AYo0VRh3kppduEESzEpHF+lLVLCL0QKzE96hUuhH0xDAgPkDMrv5QHwx0
s9ZdhcCyIzTo77ZgqqUaoBkI48JcBNS4A6V6Z9GQAnxjzZHDFCIZFrTLeMciuwa4XzkXKnHyRKCK
f+qUzCic49PkxRWyOaQtTWtTPq3hG5DTFVjf3rOeK32nKxcihY3TIZdCV7BSwZ0k3QLRvwVgFaDZ
Yytz8i439+G+9EwFjZP0bugXZlVqDbfqXqUQT8YOequZGHAlQqDgC3umYU1RiRfNJrHjY6YgZHnI
LMEUguLTJPr83B4Y4c3mFh6+KXl51xMjk1Uhb0L8RhJtMPv7TIQLs58iwPJ7wA95wMH9QQqF9WuG
yhMz5bvmtqBA4mdBQa1G6fz/woeng0cGDm5QhRphF9JRdez398fVXztycvCSONK66JZyM7ffcGa+
jNgjwFxbq3yyvgb7jieUt5Ze8oC1Kpi8WLUfil2OYV0mxh44uv+oWQ2IEy7nVw0wEuhvOHxpgJ+F
vU/VnTKeQt6pPCK5w7zxvs9bYTBZJr3FRq+gqumnmIkGINhsJ6qd4TaNlgVyv9kD5kbjGZUj+Zh2
ZR/dlFmMaafJOv/4zqvDM036KdlYcx91ok27sMknGis4Zd5r054No+cAl+AD8nEeV3Ax7wRPpcLv
bXYXORSrTrztvZqQjL5nj0yK/2WoCSvCKWKARQat+jLMbMyQsjfVIKYaWtRJ2mzUdwmvCMmom4Cp
sqf/FRed7ptq+XenR1wHMI7F0XU2rhcTQ6NaDfPNDqh45F7EaKP6WxflrERXlWZ1SYoBMfsFPV1v
tjhB778DTJ4LEVHSkC0LuO8QL4z+j540hcKRSsnnmE5r19BFGiW7O6QkHSOu/HrHOFXlerkCiVkj
csWbTd4CdrjFHNZ0IJgrXoepmiCQI3IrZDEb8CmYEN5GmhI0U4v8u7RM+0blwVTSbrslO7Kbo9Sc
g+mTs44dQdef+OM4rV4PjWBy0kxKHVKeuzctyyeb+Mpq6WbuzBCZFFuCNza5yaEFe97MKpvUUH48
vTm1Ubo/5NPTioXn8QDaU9j2cnXsG3tfkqpfzzBBTZfFoxzwTtuizM3hpitKcsi1flsyajYPSSvH
qTA/i8fXA5kQ+aIihWT+79tTPz2yxPhWm4/+u2i1UjDua0vfYYtBADfoTcZb0uO8ZE8o68gE3H4w
ipbLaiMM+EDSBIAlXmzVCGM1WwskohjWS90cvRpLf1XopczVT+xRaCbCCZ1Miw3iYfDKNIuOtfNl
niaiRqgsxV2fJd4gSC2R5VfO0T9LD08Y/+Cvb2pyvyKrg771YECW7abCxXc+bxHMAL5wHJ12ZCuG
FGtuwJEkq+21rcP/zsQ51VsmLNwtVSefrdyLpUW1sPbl/blmSsp8iRaLTdQPcWdU/Rz9cXs11rYP
EaxeFnTqKiOTC0hH0kSCQyR67tMXP0MV1Rw5W3WKdTn4fEOEAMv0aAePmy0pt47kPJBAH6l9uSxl
TrOCco35EBnwd6ESVupF7kroY15gQlNS+g2NS/otQitONqIRaC92ZQPArxClCb5VBaLkhKcCo7Oc
2QWuqZEkSGaXQIFURUFV4wByhGNvxgvmXrPEWUlqw+LvkCJHSDqiYdAaj8KrIAzpXKg5b2TgZc5a
JZgOzAyLpj/IGbrzXkmEKIqSeg9/Rg3b9oTfOZHitsKWhi0r8Rmqku4bQyQcj9kz8PogO//vLpaS
D42i+rARnAMJF032b/TbLk9AVu//vxLEWt7/e+8drW9h5shHseEjPHa7YpCA2IEQ43gouMGosrZC
CRqgw63qGtgNZbit9h+pfTCxSmm7//z9iFeUe7kz+bV2yrE8R2VbONe/Z2fHS4l9D7CqLVxqvrUq
lhVZArB80CrTfwbNMfLc4BE8et68kX7HjE+iG1RgTlfpZ1b1UoRQnlx8QrdP2KveoZFCEPB9L2jV
rDWyS5Zz8p+xmFGB25PjapYRSiRGT3LLVii/rqxq42QDhGBNNVzkcqA3colM6TtY5otJsJts58wL
zhd7S6Oz8mf32CzBoNd6Ng9mqNtHGbgTZqjTabSkoZGs4w5bOCgVykBsDm9oGWgo99LmUWrdoKhw
lQzoGO6kchIU1QoilukNVEBeTJON5lM+EaYwDNX/E/8lr4pbHBNa0DYiBePrkUSnLRCv/ULL6GEj
Lzt6/Dg0u/0MZI5dF/qvJQo+fOmCc4JIoTZ7XciHIOwy3+cbGQP606K84GyWqGOVmRTPd3Exa4wF
LsB6Fmd8KANMoPomEGKwaiKfr9CquaNuxFPyFnATHJDPLWHplY2XKUoBJ3iTWLwq+OQMG6x3sVNi
hY4wl14etNPCGf/nr+oBnNYJHmSx+NEefFdjaf04xFvuSLQn+Kxyv0W8ubITIw0hlzttCHNjGoc7
pQ1/7eA2NPO39PgyagaC4iymXBrLd2IjbFGqxWkj74vVrBB19L9esU+A1wc4DGYORu0ynr/ZZXRI
vIxKOPIrbU/XK5drhLHNBYRCFdh/Cdvfl6FTuKE9u5GoSmA75tg3/dlS/LXYUGrLnhTmih0Diln/
OSCErKjNOwRbpwOj4ICiXor+CxMvek8w0ddgijPwjgm0qfTYbQ2hFiZlzx8L52pnF0bJzfk9vv2f
ewoMi/YeCJEfELaq/8apzRZUQd6dWKcPOLAs5FsswYv4pJuDhBcnfBjhXP6BBFU08h4MLE6MAcSP
dHJb6luZPOGhcNbBS2SqQycSVh1wAMwjNnzJxMwdajvngDw5NTa+0AMpYFL3JBzR71g+vFJhvEV0
rwz4KR45H8R5Mf5gk7FB1JEdg3vuKE410JrOZYlMAHNBkEcSFDZUAd278MDEI+JrvuT5pIVWioI2
chXhLF7rIhMd0cmlDvrxkar2DNtOCMj9rNSghtdzpF+ocUnKl1hthYvjc3sSG3v/JBnd/s8Xv9Af
spc22L/sx248TCU4aXT+ABRGahCZ2E+QJgH3LRxN59whGnKuQLuP7IGrTZW3KLBcTtNLwH1QZ8Vw
eL45NOdOs4hWuZlpYEAYI3EPq7xOHsXVxo+ch0limwiDQdjt56YXq1VeRXQkuLU0qzEynAPaxyp+
XQFxt6HB0Ttk9lsHsLOuKxQvBwbMIm+8zWqlBFE4WTCl6XTweUs6R2WWW5B+St1LDZe/tYDhsp1f
WgyhH8HgaUICZ543xbwndfR4lCFOm9bzDO82jPWMO1vFEJzZUiq/d0unD4BGOuq9GyAOMMerkq6h
7U648wtiYI1y6PQhiZSFQPodsTXVXSSNKS9okwtCfoxFATtH+CVYLtTys5Z2ja2XDW0WntY002yv
ozPBxxjQacY4pCQ0zgDx8PrOB9UwDkTTiHngUEmB+csX7cUWsIbu4yKMbsndy2ISgvOEoiK4nw9h
39DhWL/QNyQpM6JJoIKt9BrJsvRYRsOB0r/ZqRpEYGSabaio70mpPEL7/Ie9qHornb7oKczu6Erp
zD9cDmraqak0ZLeTfwhf5m5w9wSqbntNz6HtYKrP2sAGz9kX7ZcoBpaGd3090vkX3BaZmYSqx+JB
466ZbzOZyOs61G4L4SXGLlk5+bCHJENxlCjcX3VNK7rxONuAqkAJ2EqfDqdAHpgscnWfDEozXcOi
/Cc9vW8PCRRyJ8ond1zbmtHyU46T9/Kh80TYkIYRbAblim+0Irq7WGnnuVtVB5vA0GCRtNZt//ug
t85JWlpYdKvyCzxxcuegdZg6Y+cK8Ewer5ZcapRPctrgAEAeSYxPaahTO/jUcCOOgu+7be5r5mKd
L+HqDdfONz45gVN0AkUJDLwZkYSP9RQJV0FXqTvH2dxhPxy6rnuqsmmMGlfccjA5yoF82InZkMkA
+xTHblV8O/zz74oFNFnhbZESqy0GoeXUvVOmtk6pf5L8U984XCbdkAgQU3C5sdFt2jCVRZcP80c9
QvFQniEbSvWlynt/uUgRKeVaL4VauLRzywwnA5lF72eAA+zz6K1yDZj0x3Pv+SME/+xoGr6dlXZl
7GWuLfT/f6Mfm9mty7aejbfA1z7rvSUUV2Isfo1xnA/6vnEMISRWbY7kGQwsbcmAszHIw8ViWizB
8G9VbbUKOWBYEPShjCzWYScPX+F4Y1z+HJhrGdkv1Ddep6L5BHOZUPEPwfb6Gm+Da6RxXn6Kd1LM
FbViWH+kbxUeTyGnNUzxzMBsYqX00zP0JEDkQEdMoZJS+GVEYn7qz0we9Lw8xs+Ud4KXzXsf6V1j
ElqqyeN5XJTSNjYUIWMqhvxgr297AM3uwFMknUelK7UhwmBx5/S9pwwuBXE8VWfWEJbfE9JhNIYE
Jk/PCsrtPJhDl3Blfv9BmS670A1AKBrB+7x7N71dUUOeyqVGJTzx2YrRKgFMktl47dWlcut+E+7j
lezFq06KBBMEKA5y9N6SURkKj2X97JdrcdP4HwsMZmlW0iXH58l66aDcwA9gJE9MXILI7SB0W20c
lhCW4Xp8culx3MMrxNSlvAwvN54JxkdY6StnWVHRQv8Xsxx4IDCQEKQ1EB+S70CAPUcCRpQNs5mE
7lFa0PVVHRIS3X22VeI3e+dBWuqp383V2jSqU8184uGuMWyS0r+kwA5ozEFaGgO96FWKTD1y8RFZ
/wzYzIgtYn2ToT36+qIW6F2BDuVMuU5/PzvxY6JEkQSDcZ5IKtNpZXTmo5gyzi/rBtgvwsKlPc6C
XIBRspDJaFYhVnb8QQPLULfqu9gVo0zHSOKiJto8cWpJBYNTVTd0A6686D6R9PGCmRQx2JkXIdT2
yur6Rl8L8bM0MVb7a6D7Nnz3aOxrpWQvFcyKSpObHUbeDs2FGArD0fHK8jYHn9SfDGTLurY/t/P6
fjFwXeyOdVF+RE/W6GHoMnXx84c/MEvJB57vp4uqkDdAojHDpKaSNtMLT5L6T44hDJMalA1MuIO/
Fk0LnKWeoYJxbJYTEQE859vB3/PI/2gZjc1uZivKBOlEpIhJ3jyI3y4kVPzAQXy5rSE4/OAEeVQC
1JZ5jyvGuSGeNSYyrBGBFf0mGuaEwfIVWKs3mFlYn1JqJPfbKjBVE+K0Qzjy6mHjexs60VDR5JhF
okVOMsSJcLC4wcExyjQsLkHZDvYXl3dHZzAWdKlKuib2wBBVCQLXtO+teJJA2D1APAdwl3IUJyEP
GLoPYkswu/vzBnWUOReQuMlR7DeWYoZW1a+t2ST1skApst4rqy8I3By9DBo15UGRZfpBFgDQ+7HY
KDDDF+e9xpsOxyYSdZzkzjieSa2liNGcEOeYDkCJwgCCeYfECz90vYCFuF43mP34LkFiV4r1bKFP
KAeUyZAlXPNjdbtJhi8d7BY42PFCSVkVDkQJv4VMYn1jiCkhAXZKTQz7OwqJvYzL+fS7uQn0tE/0
lfrp3pod9hhy2EAe7gpYjQ4iPgjmRCui8r4fwKuECn7wybuEVWR83kjSgcLh9vxQEaO7hmerLlHQ
LKLn+G8N6Ra78YeVIHnPC3ZQX4Ra4bDDmwA1H5J8wVdq1VssqorSR6naF6RC92gnRIKeXUGjl2eS
dzkQw0/719xlVgce64Tv0Y1Xwsa5RNnNuK2J/dWk7yQmatGjEkFaRNhm0AQMTPoLGsAEm9E9a+O4
rfPA1+LmDPCQ9acglODvURXeqs2ZPq7O/ssj6C7ZsXXYZK6cVNXigPGS05Ct3W6XmZAs0WBfwp4r
pqAulOcIWVLrr+fxHmUjafABus32pMcIJAqmwYbziBNHuRFUTtROFiBhCLyIScGO6v55y8Mgwukm
r87/9quqNjcjJcMt/BQLT98AgSnwGbqRUTrudcJWyK1YzoDMRGEvt+7FfCIG3VxCHVQ++l59zmlM
ZBrrNvCb7jcuuGrSK2p4TbS9NTVkA0UYVVH3yWZS9nnbZfsnPR8TQUtS8M9XENZxe1r/DmPmIDns
6hXo3tBBG6ai6y6v5VQm0G6nXG1ZYBslENdmovWREvDp+YvUQQ0JAeynX5fQkm/e0kMdjIyrMO9S
45cpIVt5bOkqsxICyhyCqgYgGM4OStDNu6eN9HitAAzynssFvmzueUmJuKI4ue+wgiPg5qm8zH4P
itPSEDS+tNPXXVT2SWRghkkIQ2z7zGWc7lydZtiFEvFEpvQSXew+8bDwQTC3l26+tVY0q647cXZL
Woaew0ynRE64ANMD6bGjRwUfAT3UIfCVEMy+WY5RZsLwQQL6h9/u8hoa5TLAHnMCeKmuguhPOFV9
9q4D/h/TZd++O5p2SixMr4Bp4qADgrh0TXsIqtsm8GQGDpPNdAia1smoUZH8HqMBnSqRMmJ1hWMR
qZq9YZe/pEftGnFhbJZ6y/ep8R1fkIKxhWQtl4ivlUEeWjy+HONbjPaSZhWFmYe60Xlq5GpJplqb
ApWAe8/TAyBmpR3XGe8iJcGmzMRVY2H1GP6cjh3QWmuoJ/+nzznsMj4MmaSouOu7ElQ0K7/Yc9n3
lCFs8VOXcUw24LWjv6EL1R97bB6X5+F4d6bvgwYPSRR63eZsVpC3BGtZxlZruYAwIZVOOaJPRZBY
vrqkyxQOkU6cRGzP62s7AMzGFTN4bqk5u7TJRf3miv3ZMjgNKGwXoA9/ned4azl+2bh9ZPVoliz3
2ZnJ/5RKcE9/XPDNuG/RQyGfLXJpJ1Vz5cZK+aFlhV0ua8Zd3uQmBnH5JLKGVFWjk/rMq967pQEI
737GjBQGaKVMD17t1viTLfNnt9W8+EkxK4UmmvUZvf78plXnTpUMXYonVqFbGLY7FWdT8rvDLu79
BOs0l8d+eB6NfucsZ+aUv5NU14M24W1HoixRMRWYaTlIFhDPOhCpMpwmZ1owFW4yKIMGNNCb3Txp
PR8yne9/dVsyJhYYx2GmiM8GOwjqnfJVkqFuHBJA6eJazVDQgEqKHslVATXluL2MqlExN6Ht75qg
xYlV2U/yGE/06K3gGOrSHkhvdhXutgB1GcIpOiHuMpQDtSsAfq8fkFOX5sn6tN27+X19LNw0H+Gd
P/eXNl8IKHK/nfjzLRjuunfIkKlnp7CuwLHSCARBYY0ZomXhT17vKG6cYpwv5es6tCkdbkcS6dtW
iFADDUenfSEES0Wm+39qDaaNawihanXuTHjHcASGyWbtpmywWHB7xTIbgaZf5FckYn2rNgavLPvZ
5CB+K10erUncVLbOTit7MB+0vTfak7c5veRUezQubgK2Xp3trM+paLlTM4rUeqodUlc0VvEnenZO
imhtuZESoU/7eYF5AtiAEhUFFTZN/Jwsh90pWSCITsqeUdvCHHzOh08M9/JYkNtmfRuX3k/1Wwyf
RW3zZ8mF0eWh9mOkbyMnJvEIYcsb6JpkBFJbFSM6oXPX5uq2paxnUdh1kM8Rx1zsaeanxjzBPew4
DDAVZ3Nngq2T1ddB0UHamZEXMvLiHK0HMJ3PkZfulCBkONri+eIOLxRKN90OiyOeAfQJX5pLk70z
pZovYXrOP1XMLwC7RuU1BlwioHJCPC2cClea9EtMVbyOiqzDvITth7MMRwOLeKzxGnKRYvxup2oO
cDMWLpur2fUUmWFgB5vvYjh4j5oxrN56qqV6z805i8rwdVNl2NS1lhTkztgygQwjCZt/iA5eM3Lx
s5JYUW6NCwiB3IFZvcD/QYVIZ8vqSlWQ4lv0VtNKyA/andt5flp8B9ujO64tKQzanysJGUDEz5QH
MFZyNs6nsnSdJV98iMw1EopVDLVdetOLRTeAi3kDkRB2CkypVbNL4JfskkFK6ijRNvCURiTQ4/X1
FDGmEQ4OLOslCPFfu+e4OZEDDjEByt5UnfILl3rekssbp+rukFi90uvp485o3sO85m7lpoQgYwjz
XFrzAA1BxG2f8g7s+DMVi5BkOR+rrBbtvZuQiHv1eD8m08akLb13KU41MzZic7VX2Jh4a7olY4A5
k5EQ2WeAloqhaYbpoX7VUWNK6zTpK5qr4JV/6MV7cPhAxnXAe4lzyADLBphrxZhDFCekR+23E0hk
6+Rzops6x1dtQIJhYFOVxjdntZnJgdNxpVcWNeUbpB9n1xp3J185KGs/kYOrGW55zlLzxWLo8cnB
BgKLAriEc0v1czLZpOvHmbmBRofTaGMkqH0B1n6QrCGTjhtwuCJd30j/XJ9PT8h84jYxJegXELgk
yHIE86CVHYbvnAg6hT64O765GGG7LwfVn85Mq2On9lNggd9luO/YWpBH9DAzJP4zeeae3Xj4NDoA
bNxZIPeQ/Cs5osfntSmXSQwfgBRuLd0h42lJ4qikgSbCbMzmxpzqrXn+rh8uNK7v4ZWT8NOHLNKE
p5EjHzRKn1tEStcvF2wNDarpFsEXeHoYGZSN4OTuTHtcCD2Fz0IYKjvwwVXRMju2vozU8/+xnw4S
FFBmyShWMIetMl2pV5SqLRKY/J+ODRYVNEUppRFjIIrVL40J9GxED8EL/RPdOlPd05EBJjuxbmh6
DBKxBuHvPOgdHNSh3ZxaAMwTVvzkcgD2HPLuc0u4sqjA+byWHtPLqAb7I/Oc/nJdL6qlgysYwgFg
AEF2w3rPcjLpuwS4xVRtePYSE/jciUIQ/UrVlw2SDrdMPtRcM3mwcgTHTeHH673jH9t2cj1d6xFp
4NmKj9SsdbOvOjH0fr9nQc4N+bY60zhAE/7r1up+D5DsHvAgA3so3rrXDuetPqJZQ6sL1tRit098
vUPsyOaQKt9Mk6uSSxj7hnidbayx01We+tkdOPtf91R6GeY9APZavVEoFkjMZX0gRtBpoN7TGHZ6
xxv/caKwlbtyHiW1C7JJyY9Ees5519ODXBGTJTb4a8ZIX0KAOmLKgKQ8dKFZr30LhS66+ZfmfzP6
OPBukbUeGhI6In+DF8gfW08PggYJZ6h77uJE104hdeePYbzgtFnDHNPcmbKp+k6uOb5jjAjMtQco
6x7P7iMgvWSWC6rBVJ6MmHq0S9KldNY0FVrAXIj/IR2T1uj6hSeDYjHiPGZ01bDLoORdCff40b5P
oPAraklT8ITGi/lGI5IWVsCunVOHcS7egcsQ1VDFbqkxaamh6BjBv5AGTIXW3EVzaqeprlCN/kr5
9GrfiDCnrYhHOeb+IPDds2H/FHY5AwMyC6rnHQhYY6Z5lW4tBSmO2G4Ii13DtIFHP3vh4+7xKLdB
xEkqheYJBImP/PACjmaVT8RYPlnJKaqMUgL6vjZl5chQnT4eASIXdETR2SUKed5UF3ajQ1jfkCSR
HvPd5XktDBdinvByLD67KSMXQ0i4AkBNB9cq5w2sVIK7Ri+O1u76M3A8QqifIzigHG7Sp9/7EunE
IBWJDa+3AIhS3Xd33Ca4xghHDY9FjVf8b/e6oieOoNKsS7y6+jr8jZFdlhZYEggSXssXTi0jqrHE
QIgLqfvJqDwq+rY0goY1nAeWeaCx1wrU2yEoKYbgGIO5H5dqcD/+qNrIk8ZB/z8AKIgXdgylv/9z
Le3uM87nc76HO1Vezl/q6r3yEwMniHFQz/8a6nxDEjcMVlNv/tJwT0xusjWyHYQJycCwoWpB6H4H
935M8/i8q+Bv/qV2HZRiN7i3+vf7eFiLim1HzwKwQIPnlzUhOICTZHJPQNc85UCqZj0FM5Z7zk/Z
WP2NY0t7DF+TZttIuT9lmtlvPaqz5Br5pbVs8ZsYhh7LLTtsWY2YIPgTabkEPDTLI7q7/hYOq9jD
kWxUgNFqoSNtoV3WjxJxi2oXvusIomQTLqnGUopkJQuyDWy46VKKWi3fFeNDjR2o3ObjSJ89pz8m
0nA02N/HIWYjm2W75KoPkmwZ8oVPndRHyoX67KZWAXv0wn8TcDjwV1UuB4lOGNMj8sA9QqjP+2Tb
mv0/82U2qi5b3qt4oV5JR93j14BHmrQWlsC6Vxka6aHN4LAXwxPmm8xod+hbMGHMWC59tRmIr8Vx
hXjJzn5p3s84/vETpJ0/UAX4SHReQ0hMTUZqSpVDevJH/5WeXWg1CcDJYe/od1m/Y853kG4qnUKQ
sBDSYHTLGqb2dCw74GVUwEsGrx6un4ejGJtKaxf9ptubp9n7Ob+eT2N5cQ9OKDcbv7kbvzYT8GLx
BAVA1nHm6yVNTsy3WvhsdLI4LBvLPt9g0ssA8IH7Vo1rbBW/lJKzrfvIKhDKMDgQHnLF4MVe4Iss
80tbWcbfrMuJh+QPjatHtEd9LsPSlIpMdKUg4IP62A6ZTAnEbxVGbJcAm4oo8HottxvGU2+89VR/
i5mGevzkYmBH2b6S3JpFf1QDlfUciaU5Y3bnDpaHvFuy/a1vL7ZptAtuZKCKLPieH/ZBXw+Pj3ly
vm4yX0XdB1iCS8OI3PUfq8uMkNqqg7FggaNYUzwUKsIn9WeF4HlKetmx4FndE5wwysQ0WZRWgo1k
GNxcOaC8iF8WlqSq8B1ASuygiiemkM634lKpsjUzt4OHc0rDtgjzYF1+ZRuRweapHKbE82Mgvsms
vHyUlBDxxfxTe1JntoyMcsPIk8pl81/TXNH8IRpw8Hs4KDNU/lsR9zqK7NWbnBfJR3W3PvE8+zvm
uV08k0c/P6xU8/pakErbqAye6vk2h7R041j1XlKeLQmkDjrtja1ibY7RaTqCou6nQf+vXuXOWxPb
IhLhudzmZP/RAZuFeFlN2cESPlX5F9qa3oLD7h4+8OwfcsYLMu8b+cTTs4fISCq6Ax3Ll7+oIOv8
lwAQRc8TUdQ+8E2QkPo9Mn3L64QNDGRz1apb1S91OlMMcIPZNGdJmRdWQtJlGjoMmgurfF8lh8nt
Mw+bQLg42r0gHN8QsKomdXHrzaV3MnJBbmQfsfcCbuNT06nvguZaWxbs9+BRi2cDn0ENOpB7vvkG
24x2p4ot1iJ6cElOvGNdvyMzU/Ye5Q3pPctqzWDaw+hCBkR8sqTwFj3ERXqrob18PhYL9aZNqTl0
kE+UCT312JaWor4OoI8ANz+Wcjw8uTCTstQMkJNBrBi9V3Rk2KGps52yeJEl0W7Ei69tsT5mzRu1
ehtAyt4kJwZR9XszO+mqWpXxSDxfEXACjuZRUGMrbgYd/jw3A9Yo1vGp+4J8WPrRI6v2dYc0V2R6
Dkwgv214+VnhrxG78EPjzCr9oCesR6vgepjylIjMTMrIk8b0pEICHlmLqDblEf363avnIMD5s3CA
EFJMGXnoBrfrB9oXjdhy1/XcjmQGE+wCTRejG4rFpd0Ft44S0kcP5N5D8+MU5tXZlZZWPWMc/4ir
fPYI/sPcrboDoa6wjIr6+d05RV4c0sB2Eu+8NESRdqTHKQOaT/yhtrAV+ZPeQOIpxtnXk2l7sW8t
Xu9UdOyQF1jMgzqvc3ds+2rGf+AcrjPntJwQ9pL6Q9Q0bMr5+MUH4eUTdOCY1Vt35tAT1Mbg0CQ0
YoDtDJhRVgrGcA2RIvrPobpuuR5ivQTLDn5F6RbHlPElEIJlTJNsCYHfD1A/iKWQxg9+cQeFaF6Q
30zsG/10evIZ0WII3F1vMjaP9qAKnAssrTz/GCpQ22Nle0xPeg+yBDSnvF4SrbJitN41HY1yqXhY
yIR/pJHV/pc/O52KaPm3hQb6xlErlRsb3LPxVJI/qO/FyzEaS3N+gbKo5iNBlQ4B17dkaVmMmqEm
6UKXMV+Ucg9bePbjFW+z86TDT/+G6kFHp6dUVhRzzcApEY8sX0XTBLw1/Hr1CO3a3UAFq79tcc9V
qqcvR0zu+Iyj4nf0wOBRyhxTd3FLr8F9/kIVkDtzAKTacTkYq188Q8LpqrJhDdA6sT8PLmAkVjS8
T3hPgjLTUKnptHiKrGNhxP7I3+6ncGc/lghyhffOScn5B1Y8W9bWk36LhVlWsN1mSmXuuUnZY8Zr
emDI87TMr78eZ2LfvUJy6Kb5SpAEQQ5TCSSTku9uD5aGKeyUsQAOeiB2o/nJeKFEFIEkdz2WqulN
n3h9XiqrXhlqjqQgkeqit8YVmnibRw/K2YCPAeXMEGzpqWRz3H1EpXebjhw8Td1ucCFyi3sHVkN7
72C8cpRGmiEdITX2+lUEiqJwuGWk8Jnq/Lix8Yl06pMyiRf6e3SS53HQyIil5kHQ4q1YWYdZ1Njz
Aio7pA6WmV3Tsj9NfMYsqqaL7ZuUfeQ8D1Voz6LhEsIRTmwtG1QN/LMmZDCiuSvztRNBaftbpYne
G/aaKt9qhqanra0pvF295roN9TjIT7YZpomQvbpxu3zoRMnHcDUQPcMbdn5Vxq6jUd1exuNndX0k
GatQCIuy/CbwBzXodShWMTxvEXhkTZEuQmZBboeDUR8snz/g1GZQ+k4gNP2xsAbnNNOY3eTUgvwo
sNn3f3ctl9WDNUsJHJPN4ORpWErMPk5IyushayHQq1jA7NCrWksxArOYijo9ZMktmqw3r+k2y/W8
gR1MS7XEa9IY2ssBGHReCYITja4Xm4L2NY5Byq/Cu2qyWLEYtWPyh85shutHwNdIN5wiMSCnSUJa
UERapLfhAje5hUUaGR4kSieN9Xd77yMZMry2y64ZmU47skJh8wT+QSn3PteNj0eqCGlvrjLIk+hQ
0M+SSqI9YohyKTUeq1m1FidVl1qLBlA9mkv/LyMXiTuKwG3TfB7A2xMkvToYnnh8jOOmebauktnq
62qIAVCmIezpDK0oVfwNNnJR9LaTOYdkH8YVZrJqZoQqUo4R+rS6B1vZ1At5KZxDvuWJsjPDDupm
0yVvTBJFVqxON6vw+9fa0cqOED62bri+INJm+RamJ9/kgbCRuihde9wEzqL7mAV+A1vo0+9IVxDd
fAq0tBgJkvVwswisMUydIlh0eVDqBtxQmAv/qlBNk/lkLy9RHbmth2hRmTxXx2/mbj10XNwqquTE
543zQkcGaeinr5sMciS6dRjkTwKll/dk6pAU5aomMFF80hQBwXiAz4mE9ZgW0j1wOzD2NIYX7s/8
/+5avCFGMNIdCx3qng9VP5xDsbzZx9JWhdCaqbAlqkVQq5aNvZc6CZRKJM8Z+mD7/Q/owaa0ea56
eOL/3yJOnauAq6m7pJIubQlBadh/+6IlTh4bmN6EB6pcRoy3oiwJ+49rrcLkJoqpKMKNbyOUP+7/
rbyc4NDquBzciROpmCGZ6D1T4UDo1/h/xDbJkXwCyXaCcCc7UZjWzQL04Uo4qlubcxcgFyohXFZK
Idp8WxjDkZH9MdAlr0B7zS53STQPUfHPh6irsg2NrhUG58pITfn+S8OYfuqDv1hN0gxZfN8K55Ap
WrayYqoRa3jn1fGBMcBJdNROXC7u/H0r/zHUH8nm032lRuoYvkgk76grK+QxUnHjiUvJXl9+JzF8
IX/vgfHZzlOPUvuFLecmI/m+fhDGgM0Qxxojep340vo7iUrmIUAsZPiUykmx5j6SkPDAzy0A9WOr
r1mN0lb23rhAvfWTNPvGLGS4FPe2kGdDsbzSSUvSmvIu56Nln6jJX+dqq8S91Adhe2Z9BB04RDox
tH7si7TRCWG8KFDWWVlU8x37azutXDygxLPqfENjSjHjdjeu+GwxCuqEpUa0a4SzI28XSgPhIj5P
CJ8U+6OukdXrkl9N3J0vSCAJ0uahyTRFDnVfwhKQxCl4Ttnr5/7u+khPeQF9sV+uCXGCZzlZy5DN
Hq2xGDmUqCx4nayE9nsJUHEZ5JcK7pa/e6+oh6/Ex/RgmHQUqw22muRxt1ECFwnTgnu9J30Y91ko
C1PUVjsSan1+SPBBinHhDUKD0XhXC6myiV0+r/rwDRgJcDsNuZIaW87yFGlHTjlzpPvwsV8hb4vo
uDQ3j7BaKRZ3TtexsylQbE2rH+46NWn2NrcbghYJIdpvR5Yvm8TH91RGxv4QldBfhWTWRtHzNyRp
KiH070Ze6gywTmAUo4CCeG0eL6rfB9NyDngtBNq0Lkj/Roy/j09DSZbrq+1innkvjjNh4VD2g7hB
NqGtsFUgQqyXvTIiNipEm45kUgmpofajWrhD5titQxvCndXuEf/JGAE0avbMIiiKRLPmLQdKPiYm
HlfUIQUFS0rJVshkYS7PgG+48Mjywvt5OlIp3gYIG6piANyuAhONfwtXZy5natqaz3a0hMca3WcC
dfXt17gnlkNZJqmy9RVsE90BC0tA8nbgsVIgXWUqaAfNQ2hz5jl9I2Pt78M8IlhMgesqHOske2T2
6qiR4v5SXJR1j17GJfweJvtkjlW6Ns2tYcq8mIum+P6j7QHlT6i+ByUzaW2s1RaIAjuJHbEHu5fR
meTfxljPC7/W74mWKFuel5eVw5I28q6oN4ZRhIsSSb8qnhFmfEAwC5O41xn3OPm9mjM5FUqOS3nG
ft0r3EEfjU+lb0bWvEEFW27oMBzFDsN2TiGgCvefJ6SINE+I6FJKh1p4qmlRbZEbjS3khuwvCuI5
mnhK1Mzdr8QL3KWrztfI5QXTiLHMtXPk9Ieahuyr/KDv0W98/PfDVX/rViLBaEmhKBayOrj0F9dl
VxnreaZffg54qHzl58ZWu+WnQT4Z/YR5nHu81fnpI9F00HQpa3cV/sfC7fDGPGoOjU6kNkPyLD1N
5b/dJuzAWVaibUlrVKmjqof6LC7cgetKCkvb+1gyQr4YZDJ8wdGLx0IjE6Wsc4ahqdjMvN5ZichE
TYg5U5/Anr5anke299KsxZFeMLfAp6/tt79hrsanA57YsO5VHnsmTMO6f7cdpERB7jxgdvls8WVQ
/3AfZaX7KlVLWAs8RUhnhC8uUhcO1ckKVkpUpLUqtC4dHQUSI0/6HWpL2TITr6YofXjfPrd7cOxQ
4IBTFkSUUXsAalY1fq5HUiEWSZ2R86j9qy/fhw53t0qrBWdjQ2+IgzcRPIEFGCP+u0GmQ14Ki22g
JrdiIYxT6ILCputckedFokhHNdhffT9NoGtFmW9sI+HZ5uwCXGgiaEZVpQhtWiTkF48l0K8Fo4Hn
YLXb51wZTHe0Xwk0xTX6q0zvpcyz10D1bRDfX9P8Kfq48DzgGCcNG/BYynTVfPwVeMx944lfLTsk
iEXj+hpYLRFsG8MF16DzotmmTno+H8CU3iLIJzdpY78z6m2sUGWYRTjiSJ3g5aQWj4dp2bwcS4eG
Pa3y/xuCnebkyqFnBD3LtOX8TcQzjYOov8aNu7EGeKg//DTEcMv3/mkeH03MfSds0AJWlx9WH1Ou
u1oshknWCGHBJhFUgqYQvQagcf0td8ifHecSD5hx3/s7KN67HV9XXMtXM0YyGKxoX5xmu+5CU61z
YPLD+BRjcgAcCcfP/wpu7bZzuaLSP2LXp+GgKyFekpcTfvK5CYErecEwF20p7ZuzgUgNB20WDPCj
5Xhd/wDpx8xF4UmPknWTzoVAufmuYah6PMpNvKXXQfPTfdzn4iOP4u7IASY5izjPBb9S9Z3Ld2dH
yzOd+OP4EsnP0rnILZ0ptsde3cXiMbIzT4+fsj2jPcUzBbFmTsdG5F7YRRgfeq+N7OaTZfNB32UU
zErnQcXzxXJ9R0N4zYW31/tNcA7zJHDbfxPq6s5uMZ44z0YYcpCsuzDKDNY1u3RgTnd62zV+YBOI
DFuoiJOnZf5qIEwqNq2QVqyz+BYxvmhkkFkxKyQfHY0JJ4lyEHfglwGvecA7seLwojQiRW1gjpBb
IzYL7C4eF1o9YT3dIOzvPPcYVahNGyaZI5PEFtuBgY/ljgrofGUq9i4SKmDI7R/KyE9A82ioWe1S
nRECcwSB4hgndjvn7ZyoTdBeP2sxPa4q+kZrjdSiPyNFevZ6Q0ilZz53PUDIgVv/63ZGY6zmmbf6
u4jwR4MT32iPDYpbbRcglnPFgFFhTJ7/QFF/bg/9kc7TP03tl2nrJLAlhhuCxaipeJ7dZL0p91wU
EcY15Xeu8iP/fzIDrJN0KlutlzJe+m9MRjarwxvdaPOVvfJQDDhg9vdKGoOGN8WPALmyiHZQivtL
eQ8DrT5rUEzMEX/PHoM0m80MRDmNhCXV0zGdphsL0Y9PNJoZeu+IQcaTUXBnBmrXv5U6ydena57s
ACr4XZ3DXKoC4I8fI+zZ+yI1BS2eDvCaYb+nKeUdiDoOtlrSesro1sXxn8dF1vyb5mJvL6W5vbod
2VJzeHrOOShlkOIQbVbDBlkTYgUu0l99QAG9vWTkwEAet53Y+h8uCVZE+Rhs2/q1bZASzfNCYgqI
s3vxyd8HXACtIbXep+VeFBr2qOUOE/TYXHzxmvKWAOsD612AgEkJ1okF+KTKT7HN9Pky2lSG4Bxa
IZl5n+3eIu5XapXBpw8aR51P7GlfM4JxIxS9iTubywYgv/MyVlI/7gFG3k2Gh4VAd+00zXLPyFdy
2zWu3DqWGR2jhkceTZWNAQ3Hs6kQIqOv45/P6I6H7JiIlEeJiC4JBwRNcNIrw19YiGyu+6FjDcc0
U614N8E1YwcybcSvLEWDpdyaX8fLIZAT5akStq+8jjWWNyUYScBDkkCNcLhyGN+jiPLEWLEyKiSq
Im1o+U1m/fDvDpG0W7ni87+dhfXJmtaQ8ruVLt5xw8hp5AxVePy8rpkqvZFZPwLRADtULx8tOxTU
tLXMBa4+7LOa9mkInoNQABWsWRE4E90gdZpg8ph5wh4LW3RXwnJhH3Ut19njW4l9erdk/nZ2qtWL
jvJtCrvs6OvSa0lVVP7IY+VjPrGohEujHFpv3FnbkATnpvSyfm4+xmLuRjLDrl6UoRoq+qosKi/E
Q9/vAdYQpCz5aQT9wzz/x8wRsB2CG+9P7OxwBfS9Yq8MLqd+Woe0ef8lauUxbyisXW7Yhi0/hdyw
FxS+22sKpuTJn5x76xO6oKFJ4Yii8VPzMiTbWYK72TfwD1+KCN6N1FNgK5YyHamiqATYbPPBQkau
v3wG76HHFAwrDaedqExBmaNWoJHYKJdmhg4TTyKL1wsehLDCayulqySGfqDxQbT0OBPvBpqTMNqJ
K2oVyDWN64v96KKnI2gYdlsrnxMr8YwIKFfglGvxRX9ZAMAaKOrtSY3lIjnsHmZrtOuUilrVCFDm
6XWgjsofbg9lwX7tbtDAan8BVPgWflaocwCnvw6W3Q0kZUQaV6VIy74CNisj1MK6sPl3ncplwJ5E
ep7N9fwFO9Lke6/JsJ0tZ5Facal+eJHNyszpeDF2UJ7xkfGkz9DnXNivA9nMEhwNbxKrl2RX67A4
3yOV4o3bzKdHBTJPOzLpsXlUqio36QMW2thYxIL+RMf687JMfCa415YYpvYlRJHVWZOFsEcv3yw7
EyCrN+yxH6WWTd7yF705poCBEwcV5bfef5vZfrKgkPbeQ02RLl+kaVTIl59wh9hz0DKMP8pCDEIm
QXpWqU0d19dDrINCQaB6UIA06rajrcrT8w7XBDcUwx9dRfalT7AGh7/gD16GccJHkA0AOUR/RlVH
M9Sx0Bf4eeRgc0n4yU3DW+L1CbqBkh/1tTEp4LuEt2F5YYIi+5RP6wo9kYgpQ/o+dN09UxEk4Hka
2o0gKgph/RcEaPIpaBJ6MnVrWjyuTVu3BAxObQkHyTCGQ38BMz9/o70JHctUCI3go0r8WsLgchHJ
zh332ZYf35AAo2hWpdbGmjAUdynGPMVGusp/VCU9JOw6qw+ir3xgWJoSwJVcElaMwu5UwHNwr6ix
1Lwsw5u0+g3q4tu28Ce5wTc6TUfJN9RxixQXJypGDi9Z704uNcE94orXVJQ3kipRyHApQU/LlWw/
+AVpgc1mq8SIjkO9sDw1g4JKu3pY0PAvVRZl+gZx2mrcMNZoP9+8R+gVtb0mxfucHgZGUSEbpVP7
3ZLYJ4CCRqiLZ7KpUNlfF5JUuVZNIcwjKdp2P0vmKQbJArDoZACUx9bWCZ6aQyVCUa17E4G7xy9P
qxVIJMWiBj77waZ126Xh9d8PYypFZwllfdYq3O64BiMEqVWQGFd9EidGqTKlF2K2GZYtL+GaiCyz
+Vqzy+ZMaJswCEzox4vcIbcL89qF0jMGyr0fM1zgogg/BOajkey7xuc4q8GPm5oqzMuvijRYuYY2
bvYcyGMzGehYokVWR/4jArpMS+/biH7TqhxxAZLau7xWOotkMeZ9WCkL/4M2m+H0cI4fE+Aj+l1c
r9zv9rKJ2NjxCX/9coP4ERKA/8Oqui2TyYpn1JDRTM9Ebre9qzBVKAiOHeFZGHOhbwXEJ2toBdT7
NwiL2QxStH8PAWY9tu8VzamAFMwML44nJ2qpZVcY72NdoOULNJ7ByozeacDhb9/DMIg2MbnTnT+V
rCLkMBdTewq1MIMb8HpLmu0/ddJeGPlfVTeaeQWwCLYt0+Cm68O7OZ/aDcrYRzSWDOOdwkPjr2Au
VjbaZr+tjKX2924c2/WAz6ZJF5cAgozuIp09gchRs/Inwl1JNWfrLz1cNW+UIp+EMHmZ8bgaRgUv
09RAXi3o+o7NY3evUejepW7PgsPic3fMIaWD3iMSXxRqbZwk9+RmLJQXyiwjQG/dEMq9SA8tqEkE
GPyXsw3fr3Nvprct+ejswfW8h3CptSXIcSfk1eEi5kT5MAdShb4wZngV5jB/4IcA7sAC8XKBWb4+
yiqzVlgFaRJ0PepljgY5IbaHQUArmiM3YMlnR2yhONeDzA8LAyjKhbFWjkDcUZYG6JqjZQoUanQD
pTDWk0d4pEvHcfjEl5FMcPj0gU75RZ/M87aXqqkCTDvhc60kk6NbgZ7v54TMknhxUqEfcZB7EZmV
ZMeHGErsTUGxNb6g1J1PlHcdSs0DI6i18enz1ZUz/eMwx89uEYFFSwbFJ3wnPUgs3JANOhhmnKMe
4cag9UPza3LezvWC7P103QqhHyuLw6Ub7UsR+iObH9K8tZcn9V5D1C0RDsxSBUDwyK0I5CPKmdot
HfXsES9zlkJzu5BOETOS5UfsCkrE5NlI11N74t0aUgSoGn/pgsoZiEzfMmSuaVETjOVSHXLU3V7y
eB1p0Ts82qNdQqAtJfP/sgFDMcxy3IJjKFSVB6NfCMCLECIpphV5fKBNvxR0ckBoQFrF3vZJl+Bd
75peSSjNYIPXMKds/1fiEiV9thQg68Kq2dC2Lesx+Q24Ha+50ZxTJk/mgdePaAPqr2YJtDQPBo+4
c4u9I2Ck/UH1ScU/7JzY/tJJpzLu7tQXt9oYTn3P5mdr+b5RZATAyK7yUJwxX3lKTP7sUz/iM98n
svTNLMkxQuVTHYWyxf+It4yCGtA9AeY+3i0uXa+5lbvd/UCxPS1qAsX+hLIsUOfhf3CCbfRPC+D1
wCLoIozpQmgTSSXkzjE8u/BLRLa/nGXyTiRlEE/9ff8UdZx9W36ZwTR8GnV2ABXnHbXA+XtE0uBc
29eURR105xdn1aeiAJLstZ+Ms5fvp6Ma3z6n3X83nt7Zp7ewcvlrmeENwK/MWtaeYJY4a0YzTLuF
iFnD72apmVP153UCYvdFq7d6MtA12fr0XzeGeLjY5bCFwqQ0+tKUG+fH4SizK1Bx/rFNwoGSe6IU
zi1MgoztJnt4zlfquVWM7sA8dEHVq+gRoEiDrsbqHYsKPg67pZZxoUuzTCsEkAMCcbisxCBf9c8A
CJiNo5df0jlA7eEwiltMYT6aOejkZNQIVLmRX27QZRSeFeyYeNaaxmWbykY4ptUCElj9n0acm19g
9GVxy/wRabHy1v46EfUU8cheUpUJvylYaLDdcSaZ/4M+bYpQYeZBXh8L6zMr7hX4fC5xi0sXemws
W8Jlp2V//C9WKq+DWj0UyhilhaoqiwIaYBc5CUry0FZ61rWuA5qnkdFG3dnrOWQKjFSZnMUjrSJ2
0FmSHa8fzlp0btorw+HqFQtgYheukEY8h36V3QeBb1J87+juBgnTJPjSnVR88X5rkLjMS1fbA8iT
5+90Sn9+dTmc2MAYIcx8aJshT3ARDd0FLC2Nl0MZz68hxuqRtvVyBtppZdKd9XX0TlHclrZgrxtv
Vav7wC9A1ZYncNaKcer7fFJv8TvwX8ScFggMQtfox8rjpkpdkvG0W/DKbZMKzFovYclzkTVCS80+
WwuPlNXLrcxMw827inj82KO/J2m0WupU6Fn76QXjwfPnhXmylBuITVvJMd6CIMZYwZorlp99z/YE
yBEcegPdw9HNDzVPlgG15Hj715Vxjva4rImKS7iiUM90Ne89q7DFVKMwoXft7cFmu8qFZhri3F7l
Z/5Lus68dcEcsTbX+A5L4ot8ADoa4uZZ8kL0+7cxBFZ1pmLElYLKUErXrLwoxIV/Dk/XelHG/Ctb
kAylo9Mhwo3rVeXO01ieWzUmZbq1KqKl0txisZcMFL5Z45QpzNwFBVfrmpswyDu3BFj9P+n2Fh36
C2BQvOaykWKThXedS5OR1B20iqHpJL7Nb8SE1y8geuCvfGB6uLUYm/EI9arhe1p1Kxlw2HQbZ71x
UqHKCK42+Ub/fXexBJtFZFXqgr56FwoVjcVA1Gxaia7qmjzFERNnN1G5L3/e/QczU5uENCRQy8iA
PP6dRJM8/kY8cbacl+6t9iShT4R8WlBKF+HqsjcU1QTBd+u/Qr5dcI7SSG5FVjb3X9fHGJs8wtPc
gYI1uctEA0VPICmyOQwZxSxNaCCyVWz7G2ti52ZxFFmD1U+8vBo713eaxIyr4bUB8aytvNYThi5t
vsLclF26KZDqSkW53REiuNklI1/xq4gLAJst48owlTmcy6ed7t+Evgf4lLJ0gSz+ASSni7Dw4WmX
hPNQi1LobVrysSuAZYSUg7xoRT2ApOfCbjQcVN81jadLC2Oo4LUrwVAb48a5IOgT1QvI/qnvNNkq
Zlp5PnZzfvrwoFtbf+oQDCGidCJncDORFZHOCNZoAZXG69hgEo5BN1qJttwWmezuDglmnBeARNvW
MqDgBBgl0eed+ulTS7mt9FNVrEjnCba0kZnPzWgteQiN1lAdYth5q4McFQx0XRHROV7ptOvcOEwB
+KNvehrwXiDFWW8NZYP9adIovd3+oPSNuCA9d+zPkYGWBcU8gHhj/yLadyZMqH6VcG8aLBn8pfFV
l2Xr0KBbqm/FQCVlCSS7/51UuULWzTBZjdz4XX4UKKQ8+c3D/zL4VEBawlqtdE1VlYEGYa78s2Vt
P2csj99oNGtXjCG4Jk3XDsQCvyORr2pHsFn9UPVAN2jSye3y5IXH9WvdOJmml323jGT9FuquOxG2
BTOfRAw7rtiuPfXlFpvZiPdEVAJZsbiyjV9IU2d0STEHuTtRxw6AAubbEEdQgbS0pwElwxn1SYJ3
ZrWxFSoBlQ7S0J8nXxSf2SwSD5rApebv0+Ryus5LGey6FCglpA9ihmbXkSgU53qX1/bvPfweJoqt
j5haV9U5f2u0VkrMrwDkDDYffc+BOls6852gAOJSRRpVdzICBbSkhnHQI+GHEvYYRurNy1fRlhuI
2684auEQzd2LNdeV0K/4NSkuWk4V5vuuxY6VRSXDs1CxhaZOpksJnpVo6dFs1r17vRE4mvEtwqzo
dudSgDKTQ7o0/00a6ixv7hgR+2Iuf/hWh9MI99NqzDqw4tzGiqxbyqzS0zgEd4rifpAAi55GWtvk
zAr0Ss6mjf3Fv6i663qVFe+0b/EHjk1SLKRCBFXICEqdU7ps1tCyqOomnqxXy9ivifnX9mXm3yIw
P9gREvFiEvJMYwtgpSxh1pTCSZ9xLvBI10rGoszujKz3HYwenn7dyGVfwLPxVM0a+nzdumFZxwxO
Xx59Udg8eYvM0nX/AbfkTtl8DPpsettWDJOmMEjKRKL1LcqU7O/PZnzIo1joc96sa56cPZNsbTVp
s4WVsEedVvpO2jWz7gQuywhPSWMd3PfcZ8bPlC0XiHgIYWVFIv2MsagSXGw28MXRCvDlcLBrd9G3
2WGV5aTWSSwJod8/AXx+QwgNAwVagT1HfD5fKjeX7XwcJFMARu+2d7ogVDnvwTwMFVJFwXV8FFcE
NQMW2jSjQbbti4ljkvHASzEY9BDe1t+sHgF3Zn2L2JtvVVpGz0k684ba2ifrSqFyz10rbvnQx4be
L2cOh4UJF96gH2R+BShh0SCOGTKQVEZPk7HTUkE2L7aTurkm1k3mWHSZZ+Qnu8kcQ3+l2tKvfJln
r1SMWrfzpJj7u2UwkLARDkokUV95fP5wtoLiura/CsD6z5b98cuPNN2hP/kngUi0VRr5tEZabqBi
VP6uzFzubzaX7MO5lc3taAjtyJ0542KjethHEG25odCdk6ncNtlRAZo+69D5LhWwzdv+KvVRwXT2
kXbBA1To6V9WN5eKo0bnBfSTeJRg3QQYNtJ6siV61Sh7RsvsN1OsdcihXYXqfV9c4HR08joF+YNM
WRqxtMoooctLTyS1QMyoE23sfkutdXcBP8rzP6IFdrPWUNMVivr45oC5jyPS+zJo79JVb5EFdpde
iOpm8xWRVxCW2o1tTWrnQfGIV1hT55rcYgmucKDdVXTgCw1MRnr5n85prq3xIlvVxqic/TNAovA4
heFE+AOI6zMdlpgWSkygjnoX3IHwRAS5IZvezkjhz5p3uAmRpPTQ3WON/Me0IuNMoEjoI0ByShKu
F3r3Q2/sIcq1gdZzzSnrGFx+9BkmW7lJQnxOwU1oaMGrmb51v501CwnHk1huDijwtGxS0TmvQv4V
YYqaE2Enr+2RE4/SWVuiTOoxg6HhLsjBXY2L+tNn1It0/ciupWnfKE6wkIUiHinyGX+LFch1K2LH
+kl7kkpf8WXH4T86EKiaDiGCt0zmBafRI8+f9p6xZ3/ypguBQF745vDk6CmVotSZzlGqH3Qptfy6
M4i1kHUn3igvq0oiSdkcgybsronmGVMhKelWRMhy9un+6Vs0tIC1nW1jLUBEofSLM6Gt5+GrFC7N
ir+s66DRQV3lHzdaXCDhtbBFKWapePP4B1+jpGyRGpC1NVB4Ywey6BRJ3eH9Db8H7x1QYs1U9sdi
FfYAt6J8vZPN5gDyOmNhaGMW/W+d48Mh653HK46AQbh4KchYtSVTuQlZYP9Do9VRlSUJwSLma/cF
sKHjpSMR2PgA612FNvU7QDwiqRsX0vwbQbg2GUqXnOVzcvPokRP90LMfj5WOjxA01dkvOFCLqvkd
KNkNz7d47U1gWCguGpj8ftF0dIA1aKYEZfgBISa7Ct7gagqb7qogAfbhjNpyIl6oxzTEMbWznZJF
RKWPFu4FDobnsUg6HWboiR9Pt8yTZSkvt0ou1lblgWAzaLblxTaUg9cs9AYUuAdPnhScjgmGoIZH
f8SwAJudw4Yjs1tGd+D3FdqM4gFHxcHUq/MIawqopNaFDinHo2K+VY5eqe/lLPQOhPagBmIvMf6u
26irWDYHu3cG7zeQi8eOEzBHgdPkRbknC7alCDSbQiexuns10a2AYj/Wan1ehWkago5853xWv+3c
2eZwI0k69nghIv3EHWUboVbn7ZF5nz3BxPs/1kP+Y7oKpkqILnVeFiDOaQzy0n9HVwLIgLvCHVQn
tGb7csiTqOSTQdSeGXhi68x6PwagedNou+XQYvKMUZZtxxN2S4XGYYLXavAfPsUJKJb2aPiQlbpG
9xB5lgSeSqNT7wyjGRFxXAxBNvwiVsisl7fp9zvXto7Sb50d9Q081MXCN0vbiZMEH8d8ZvCBH7sM
QB0l5ze59jkWDZNNYlAw6mTFsJ8YNfl2uNv2vjicxW8BqBE7H4nhbSG0UKYJnNxNQP9j+S6oFpL4
TRQeNxlEeIdWkCuIhLe1NJEzZWk22RepTxcN1owu0ZseqsV+9Euwnu/nuSYP8bxWujsml8FT4WwI
/617DlstLYlX9rvzI7P0PXc7PFckYTw8tfJ9L8/nyWWRQPm/hCUHxvVmKLXRWzg+v/0ZUNLKSI7D
FQJriiyu5JjWqvtcl1egPGrIag05RVPFqzCUeg3Hkg35HulxKgydkcaCxS+Bh46XcgS2SLqtAmFF
jp3+krZbbQT315CSUpBnBYE1YmLj2p8BzN10xWmplA0iuERYW5xrrPfMckEdBCRFMEVwgkauzya9
jFx2hxtLaM/bSFM0aWFkn2wuN5V+bGjIzeV4T0SbR714PI2nlbllDROYz64zWYig38Tu1coFpGt1
pyqqk6kkVKFi22XXZ9+z53DjX7eNhW5WrjZo3Bc8DOBTt+OZBQV7ruRs3qiTTbVsIHwFIpfRKNTX
8hqaWnYHf/IMriDkvr1nLSi0ev6kRZfb7+IMqm+0fLI9b85dd0Y8R1j8W8r/RPquZRfN37PI5gN5
b/DcGavbP3SqL1NzkBhWtItg2AbnIdSeWxO0dW1+WZGZt3a5pNFVwN6ZoEblX0x8ZFE/YgXyuLtN
pytWhPV/hAVR74KBe8+5mPVU+LkEYJCjYO1PHN/M6IgZHSkdhTjJmF1NbfRmGQsQ1kxkHQHRaM7V
m6UgAZPMuJb0mPP/icK6E8erlucsvdXyMjveFLcbPsA6WvwQ7w70IBVh8NPIv2N73BiJBCWfCV8D
RUBZVAwpds5a/GYmNhQ2TDbNdOWilDnL90yRsqr26GRRpE9PT3IFBdzBdjPcEQ/GSTE+iTWgy9Mh
8YReZCPy6zfkCGyydRKGdcBi3SGTj4IFoh1Uig0p9OYEBaLoWSo73MFFpNZSmzrB+tNz1MDb5vxR
9ndO7elKv/7ffTGwuwY2fWcvbeNsnlQ6XR5AAJ77XFZIyKtRXRdvacYx8ARAZIOy8BvEnTN7MVNQ
DsJSqu7R+EqeXznNXCN88qfrnepUd294zNOTdTCjeCFN3eBqE575lh8Ds/nUPSAp8jzyIekpXwQC
S6HLbpzCXjLazEOBqMdR8LStD4FzpbQmxlcJjBBDD83BYeZpmKX3lQ1eEOjiRaYJ17c7wBq/NjGp
FDeVxMAvJcZgrFQSYzRKbtZZjvIpoxVKcSwoJpFFnkKUtZWv6ifL4k9l/d/utJDyzXKMFlAJMBgu
pYEpygBzJFxBkVQe4fUV+4txcfJAsun94PqSx4tYrsADH6HKdllMhpV3TE3yzZ18TU7mORFaGKqg
wtCGRqsfmKiLB1uWSxvGX/8YZOZrL8WIA4LLUIyGn9v0QPbL1UgdLYS+OU6LrHLIE6QsWEmRAuCW
KYxP3sYGcyuwhjmUCkysQURfwSzXWmsNx9nLGnbrtD7XB8irMNMOFDRV/uEXdqr4HJNiD2OZndfd
tgzUsC4sGODFUgO8TJP1+aPzHwfnNPDnoUMBgtsY5FxFW5qUJJQLCPxyIVFKK+LaDmv2zh0cdhOw
rDkH6Mt6loElXX2Xe4p8rndG6HwMVemr7aLgpXn/VrbvR9gCibeeXl3X9OlkEgb1qAApfla9W44A
TGuHNzCrKhJJr6e934c/rIag1Yau26JhejAnchdWXF9hqnFqPFDp94/etDw95R4pytsgr4VXopd0
5T7Q44MyWBSL6AdqD8Ghv+W1OL3XWl8Jq8m4AQaIu07MtW2g1WmVc2z2cNAL8NSx5WGnIpMtPPDA
wM/NxLS/+EZWWpcEo5+lPebatoCvakgRcJefgJRpFBEpyuoi4AKo0drpUu0d0D80w/a5m7y7Bw0p
btpuOoGl2K+WqVIDpgJ95pvQJxvoHC9B9yxz3L2oFMfgdmT5Rdl1w7UAPW2H3/J5Tleqiy9/mweD
taPJlrl4huLy2ibAKvXTyhbrS86Yv+3kYGh89cu/kCChjZ8VpTlsxkDynGN6i03xzV+UPSgtiONE
a0tkp0fdsEq7Hfm0gJpY8w39KaUXrDIKZ8b9vyuyTMNltk3ldydYZUMiFMYz4Hv3/IGSrwMq+ZI+
Cnv8bULXoYUkGRo1j29A48WAJJb2JU9fCj9QEtLYbBTXQsZH69pA99WLwbOAvkBGF2sKOS2t4oUX
/JK2PeIo7xlBM0L6aFJdXSfSWzQICwVrrvb8busxvdQmefsvmYAzuF/lbly7/wWxhmU2gtEY9991
vWVeXYImwA9ZGzqMJcN+sjj+U4z5DVPFl8zmHfvGLxDFjCrbOramNOCPlCdKsg+svFO1nBU8CB2P
/8b4GRKpaG0wDghKjLnmr4DCztmguqBg0rGWqYkQthuXhOr58aWJhn19k5D7m0YFLry3soW4QUVQ
yQ+dYNaDHVzGC9TBG6vPuWh2N9/r5pDf44taAd5Ufakix3ouhE0Bw97qnbMA26+tIpxz5eQznSHl
4P6N6ex0tRCJSshL/1G+CBBWoSvqNrzIrnO1SrVk/aOPuRsnJavlzVIdWIeSTYkuav1vC6adypQ9
49MgJrFVFianK1uQK1/YBEXjrwfSIe7tK2sBMr2EoWUDBaenseqZ8dFuDbQqvuPyZz1QEIMKZtRs
w8cQX6b55deU0wc1/EiLjMHsoIEBBJtyylxZwi8PIGxDFEXKRpxQZ/7FE4+52iekHoCtSlasrPXM
WPvSml1qIJrRtMuonW2tJlN+EADQI9drul3Q87HlL/AMYaCG+yzYMJvKyxjb4HmojBtrk/kRX2WJ
MLa9RkcZZ61iQUjpLu88OxfE3moRPRt6ioMrnlHF4tMfFdffs5KBk4/y8Ef0Vcll38plZbWCYSqw
1SAVgKdu3S4/RKp/2e+omG3retMDe6l82NbVF4J+tvcFOWyIPWqnw4nniRsvArsbu2CoFnMILG/X
prtwgdfUdEBTsfZu6+2VPdRefNFVTA86LGQm1FR1eyP+kWBVkzLB/eQtlIfUn/lNt4FfLCGR8Wo4
HJ60KrtC1BhoDuwBZdarVMfpTcWIJCCLTtUrTz6Sw2mc+3ouG+6aZ385CaO8sV36zi6jhh9/QrjN
vG/xluFUS/opzkf6pySzKNwBzgZDePF3Ylq2qWxq2iilTccuO+NHKyPLj7WmSCFYT0hrs0GRMJu+
QRE2V6EtmK1VjtlawAJPzhpkR0atTfxbvPqTSfHs5kO0D7uJ21lpw3ANj6xLcsfsrkNL82QwRiTk
fZWQzPliq11DDZGgmNn/utv92hS5Nd5BeTvkkfvf+iYjfcmtkvO6BavKfr6Bytpe0Dfce+V3FsJS
3JQVmekfsUI7C6l0Zdd2HgzNJysY+/rmk4HZl+s6TV9Kibs5gDfoW2a7TIcfk26w/e/nKp9g9r7o
EyMy+oTD+cekbHhaTNB3OlRLaKfxMKNUBixGOG4/gMjGG/0v4JzG2z/1sStr/Hu4JjUIcESQjiUY
a7YfTnhO+m3ADCwuYSTi4Vxaue7vNkQP4h7IwPBH1h+jHsXVydnE+S/gCZHNw25FXXhjnRdduhMI
39fdJPUOvTe5fStceEjt+U7RhjH52uqITHtyFHOfCxAJNWmO138gq9YflBVy+g1SO1GdqyD5fBwl
LlIxkmeQiHDw3rXhN3w3IjYRDInZC3zChEb5Db1iy8puJNAMhebFTpnbzSLc6z9mWn3CecZ5wYeT
w7YTKyx7pKoM92d9ADNcgKQTa3S4s8vFlIh97e2EoM2vi2jh7++CcnykeUf9uFbz9+vI+s75aUxX
Jq9MfkSvtl7wkA/+DRojy2FemDU0pI7bKH1i5RNaVR7Eu3A6FyiahIJj+L6pRqcViXNjpMnMrhS9
+IVFIr8XlZ3i4zEK8pkaUlmam7Ec4svLiIbbMS+Xb5fvN1SNEWk/rI0CO9NYb7j/mnsVu9zMNbDM
ECMhjx+vKn7vZdjMG9TVUEkxeg7GF+29X54DQqJ4k+lZQodrVzGHUD7wyB/coKIZQguBUN6/DTF0
2lEad2qPLfiNqOVDSvKHY8ERZ3Cfv2mEk3Sc36t2aeO8bf60x0EIcvyrKp7NBtUoNT8C7PddVL0v
yPtltJpRtweQjEP6dpjnkLUFRj6M7cLq2G0I7zU0yvQpvuU4gCzElCFA/m9tzD0zuHW34wM7eXSU
njhsuijjp3gCK5moCnQcdiR98aAnRDAla1hOWjc7Y4Ni6P1MMTXS8zpHoIaXiBsM9O/uYxNwbms8
fGz14GT/KSRRjA1lU0tWhriUToZDTAlWAgIfzZmUDPWkY46wtCwziXoNPCA6daRrNjl4r2WstxHp
Eoki5xNhLSHoQUhoK8icpZjxoRq+2DuqZbgwJmExWzHY9R/bsxV+MnQ1RaDogCLJHsFCRYzDk9FT
pqwByvQRL2eL9SvVsWs+PrExlRqDyT/auw9XFCHkS/koYvWkK5mQCQNgNcFKPGR1ZZuwdjPovUET
LexKEnsxzq98zEM/DKO3PeeJztQ66FGy3JqWyAbOfpyfZSfx5xOnRo4vPkf8LzY6+A7jczfRJvwJ
xrdCE5hPxBYw8cGIVCV7LgV0BUrhFT6g5pky3SaElvOyx59OjqnjErjYNrCjc53AyaGfKzjUreqL
NovMTA2dSBHgi5+go5QVQMgfTNs/Rnsd96OfUFYUlqYI2S+SD2kt0Dftpsn2FjiJw3ZjaIdyM0HU
rC/SqGAC0LBq07Ycz1Dj7MgjGY61zcnCV4c7NACrZm3Cfy0PWnsTXYmPDAWVrGLy+apt0HJOLLo3
V3kJ+6I5KPAhii0CkRPNjGUBeoVtNJm1pAqR0zKjXDoQk4RReOt1eLEnucHIrU9xv9QaVwFcqVwH
s/LKpQBAV/m7gZ4UNcwxBdqRIAlrRqeARyRM7HfnTppHTg85Zn6ihN1pDvHbmNFp5jaag1gKjxDo
38QIfWx77yD4vDWniwBsx2AU4vMHkfNkcUHKI+gG5vYryOwim7jlkKwAUC87vlCL/PwwkGHYEWup
LrBUvDWjGPcdrWsLMrPxuYeYDXHzKWdIIGzOloKVGMIx6SGRfTa9cd28RrvXteyrN5auyPwm1eDH
mlIjm3DfnFXV/4b6HujyB3gtvcJ/AGI1wDZ/iF/XhuR3Ytq/G5NMNPEhZKwQw/gw//KMN+27P2lo
LwCUZwsUWDKCjdsELe8/V7ff95vQskLbB9brwp1cI2bL1UKYCviEAOetGyNIYYSLdTlIfVYnFLFv
AX/hawA4qT5Hb96rU5QjePyb5+PoC4FNTihi0N3izE3R6ub3h7pDRAav8+oDY0zMXlveUqgk9G9a
uIGJGSBtmNPGMQWwZniBT/5fO8VVJw29AG/j9KXGiS3FFmOiS5JBYMp3lzrbnU2uRbnGAloN8R/T
9QHs2ZpQNkRh7TPL8Lmnc9x+RJMqg16JxLXPvz/hC2G4rJPzZPksvgE6W5VHZ8o87AYgtsEczqLq
1DhQvHe4NphV+NP9++s0aKkhtJBj5Mt8n5jkUnFT6x0mxGBTqUbocRENXQWB5AIN6SW+mhg1WSZy
BRCQ/TXCrfnn1OUE8kNaug5/4tnZKV6gBJGcdSR+KI2tea3MIQgjK4U4alDhXGf4oixlr/bdap7u
Gn8TiS64N8SCvbuP3AXrVvO1D/B8SaxYrdDJ9gRiC/JKBpCi6Hfrj1T4DHX8uZ3S+kGIRMvrp5uD
4Ts1FODVSBJ6DGxRG8Mk/dYM8ADz4JbuiGJdhiEvOIiVcVp7PG57aTuEALfHgg5q4H/XBBbDyi8b
QBtRuM9VprHTiT6G5RUucdhwltk7tJxcGG75DlIrCr9lMCSq19dAjWED3fSNgy9y3E41Wd7wwycN
ciAReP5K08/D0tUM6oSluIWINqSA+Fl7VS0HDBnjfxmPzLIyByhvMLDCiNyeKa5e4tLaLS1celCR
HeE3p38Vc8xFvLPZqrGH5bd17tODLCe28i5gB+n5unVFV+x+iJD5NXPk/XZz1dECNiEADiy47h/K
AzDPNdbphff3wynCL2urJQf3DbLlrYWGVa5q/GYf7HaxWJ0pycjPLIqovXCIe9Qgv+hUsfSmQg+g
Mo0W8XB6PMq7nuBwlJx7NwGhQ7vLLx+qjxXe0n1+mjmVB2/TFkhsDIeLwaSva81W4Oz0d/X3b4Oq
ucwrCUE4aBWo4DrDW89psB7eoN3bmKbx64mfGWX2tjhSanRN/hl7VcVT8nC5U16Dxb6ciRZHwZWY
RWiyTtwDcPw4bFn12ExhD15a0qMJx9RkSGdbhQH1SVEhPqMP0lp5rtSF16RxAfI+pP5KZX/HNAU6
bRmw+B8gMqFW6KlU0pJLhr+oTPr/twp1T+cF0IiQJJodqcupcEqju6N42H8NNy1KJ/hh7WqmAmjI
7/1ygFBCPNrXwf9OjVy5eLH/ILtkN1XRZMXFGxcSk+7onq7XYxVSQdLjMG1wuZfC2DiCixrlFzdc
cJags9skmTu8qaJu6OOW68/3e7749wvkBc6G04gvF11aKYLpr36eOxG2+7h/vOQ713EUffKpKqle
JXIIYpDYaCzrOA0H1aLJAjwyGdV+C5mac62JBfiqBHy7MyVm4phhOn1xozv0Ox7ebvw6Y2InjgY+
+kuGNP68Es0WYZErS+kx+fay6OJSAAuruNz2mjaCH1WyOyKUUxCD+0fCmUid3bh7lA4xpMbxkIlK
nAzj42T5JW/y0KVEMnDwucZ2zPYHQiMaAOkuq1GHua+5pynB/NL9dFjfwK2YIoLsZqBWCTYq2a17
ttkQowsmS51V4Sjc1mZ7NdlmXPxTIKaDH3ZW8LZAH1ke+HKBolf3iP3kzHaO4HQ8B8DBHguK9J2X
5DPNp1x5ejun8aE8X+yds4EHMGvZ57/w8Rtf1m9D+Rl8zwQTJBbZTNZJmKZCFMI63/sVru/Kl4Jv
Ehpw8oacHvEU9CHZvolcOasV0jU3Lqi35mN9FPiNvNaywMCZfqDuY0zbHqF+7SMWmBRHz37WziqM
shT/KTCEHa2FjMLh+Xi2Hupp8gh0AR8APWvezmVNg1zQR14n9QLajvW97Fi/lTuuSTZ7MwfDDXLw
K1mLT6nQGPMX37Mu5hxiNj90oFJkla9/IYEbQ+RcoHAfxuldkprOqKm/Ew9xJ59EgkyV9cgP4Ci3
plRdAdhj4GU6ezfs5YR+LwVM3ZGKCewooEP2tEO+4bcvd/rIufFrkIccIT/Og89g33yFjAO/fMb5
Sp1tLgGYC5ZkdigbhN2PWSIzv0LDLgnpofmQUsCqINWO5XGino4XAugEb4RhC4TrOBQy07wQchSi
obPnVKqtqSpWF51bt/uXpdEX9RJnAfI74gyeEbS0RKadbi1RRC5L6AUFSx4YywbxrV9+uefSkigK
+XrZJQekwSK+DkWzMJXcAicLEwySlOO0sqIvxOPp2Pod2Hy3UHPxZ5ShjHENAhyLRXH7/K5hJqxq
1gh5HY6co3XKtHha9z44JT8iA8mwcezspycPvcTO6HeZ3eglMrnrcHT2T/4pCbnSSdgajWrWbF65
mOHpKggUUZ3FoAmko13qLvTIe/7DiLUvN+SaAYVJSV88e1+3rAmKzkMJ8sMd6julyrwgSQjh9qWT
MpMNMpKajuCVIGToqsyvBj/p7u0Q37NnWSE+7jMAtDjuP1RIlgge8sIFsWHO5zCQM5M4b/JkcWET
2JD6njyFJ77ZVwZJ0MCjbiiMPqjj8ez/A8aYblEOKM9rKFrnKf4bRSwGmW0b9LprZO8DDyWVYAzm
hUbbLh+5mif+Z68L68UX9Z9SNdTNfqq2GsKSE90/nKMJAjHhLcOcsm2aHANM4TG8aNmdMEQBh6/3
u/FUqLqj4Lzd6dbVCT8I89bugKddyiJOi6xTK6PNUgHpqFoCC5IWrMLPWtt5bu4IJJJyJVsdWHL+
gd/aPhoZ75RaDWoYpOEUF3M0SGOaY+v4vqE8aR4jqRG+kpb1AyRs6s5KWLEyIBrlFR7RaTegnKf+
43xL4aZtCBb+9lCT6m9y4MUdHH/wmP3rsYvcsRpjUDgUsshwLPMgDjJ6VEzp1Ps1v16k46zWnMTc
+L5jATgS5js9SmSz4ouKykWUYImr+6aWofJcHyd6XCye46byAmPs27dcIC5RhEVVxp637r8sQdXG
onxnBXKZFezd8B0IUyaU5272lnbLXJjAbGUd39XRSf8/d9OuVZM1p6IWhZkgMIPhQZfx3i5GeK0L
yr6S2ywJE3IkWUqe6NVMB6Penw8niOyUQxgWRRoMx+vCo3EsJ4M9ODb/Yb39GrHil6rtjHIivbnJ
E90Pvrg6ia6SnKpKXafzzG92S5GG3GPVRinRzUw3YxyCxiPos5L4UARXFD7L6BlyVuGRQVlMHIYL
bHnZse18Kntt80Cd2UPn6zq2HM9vu464+s/Pbs6Ye8KAjgtMnP9YP6T4EFI7kaiTDqtEg9Ua4C13
AFkufSI06XGz68+8a8tu4HurJuOg+QBcxMlHAg+3dddA7UkpgzDet4qux3g0cu4a6VLbyMeQv7vy
nPyQcxLWdrdL8hKPTWzw3wv1fGh31alVaT3cNa2Tk6eSfORrWqaoslLUNtbwyoAAejFmfaT4Kbcn
Di5SCqqSuGzboLBfQtsIt87AxAS7QSjCbGiE/htFOZ3TtM7OAEM4DSnjoC2ya3BgV4AiYixwxpcv
GaraW7k38IGabIAwsoCDFMPC9qUtAylovg5hi358nRf9R8FtDHY3SMBn/0k89XBk+VBnsD79zmvr
k3Tduzf74ln6vR4qMLulf9RpzkplFKSakfxr9q8X1BnD0pJ0zT4fV/dkdGxp+CDPi+FCFnspQutc
VdUdTp6i4vOHXuzd4THHlGIh4Nksn19CBM9ngzgM1t5kTj38yWSxnfVEghPB/LmM4DHoxSwRHFpj
H2XzKD2C2bbRScQsV35NOa/qXrvDp2xlHDuqQ64BuiTBNTTsmW2//j4+2imk0pDdstOIJ/8hwjTv
YGKfNe9e3ZGQ13MWvUYsD96CT+wBYrkOMr6FrSbmhq6/8ysmy+k9PjLvhI1fmSxkXR8qpzPuIbuC
Ac2fuKcn30og7mcWHntjF0OBdfmTMvMBujXp1+3yjJSTIEqLEg4Gpe20Krc2Fsz39/kXA77xcHzy
YM2d4U6CfAuc/++IWoZNOE8RnNlRFJ8gPmSkhrlN3B5qyJMQS/NMfS3cDC0T+FOPGBaP0GjxiMRz
9Dcaz8FWS7V82lTYM/KPeCVVKRr93+5+dXO8ZCzpSPEqgqjUsE/qpXJ96thIuBwyv4WLKBPfoAqU
4f7XgkaGdHqwY+iecotiqN2dTLWURo7KbC9CzyTqRFVJ+roRh0KmhJw4MTTxMYcbwkdDZnnCLxjB
Yjc0lhesztqRpgZTdLbOAFULHSRP0EfJ5ZrUQ/xzOB778NfaZDLTuWUQIdXk+oAo5Gi9BUp9Tbqv
8MMnDokHmAcP/fknkcz9WbLwuCxDGySay4Ceet3H16wot2R7uMCChfFzyJixyUNDbiqZtauU6H3c
CbpMRbTMycz/8q7u8uJ0/5g1Oj41L1l6q1oPYAqSaBt9UuFt0SqH82P+tROQYNidHnwHaBbhkcTG
JtovkYV2pFLFNHp3hxUagtg7h2QIeqZFSosqSHheW4OERyjHNMMLA7SqEmRgMRfJghchG1DDSZKf
JUkm163p4OE7nqLCpz4tg3NDOLYVW1AMla/LgWl3zjGcz6s5O/rpMSK2bDnY/xlhZ/TWO5N5RGvI
kS4mnT5EpO+S/Z8TSILRUEayWfphpNK5XRc3aXmUrD9/xmfvVExZAc1ap/TAnqof/pdLZCPz+GfD
ohzXt+emPUyiCAB7K8zeFL6EXuVfUafZGKQx8V/zCQ4QxB/Qf9Gs7s4LMTWmP+aKPCOT2bduUCrE
XwvkdQ+ZIMkWeG1TXRWuwrhheOGgI1F1Pl4/EbYgEfh3Hlm/dA5NLgbPd3iYyksxgZi5oNV2VDKN
MkumoUM0LNoci3q3H7eXGcBssHTh1anqJwr+TC50KHQcd2g9zeLb7NvrUNy0iOEsytyW0OaJTgUl
9yT8NfatBA+yhigGsWHwjaA5zfANegmTbfYCyqIuXapTPh7IypQjSLFU58uN1MRvRnCp2kQ2W4nk
rExW9zy5vmQNuxgwMGAVyGkEVddJqVj+Q4eS3OvrID1YPdS/X9D0ucno10jIN/dtThFR2FDJlJwv
1nWBZDE8Nz0mD9Gp4qg3CinwS4lhBbeU2kCwzo1Kbeh1k+7QGhr4CTjXBe48zDkLqcP4KEGJ1KUD
NVeQgxE/vKrpK0wnXjil904VOOl00jcF/lQklD2maJtfr8SN90wDmWBVOOtbbLB17Kh8MENqlmq7
FRAL50qgEjoP/nsZHPpdsQC2NZE4D522FCOV6t94kidpAENTl0rVBQkC2a6gDOQEDVo1Csxk34b6
THA36z8H2vVBbTIg2Lc9PCeldj2LgOQJMtqSbkZHu8BnytTAK/O1Luz6ptFCCmojbR5PL80V/I1L
eS1ihQeRmkuSebX+y1HdyqMz+xybTHd9SGRVeQC0HGkAqf73WyJ1Sd/c2Aaobyk51he/nS7Ihk+K
0vMj7uh9wZsLc/Be5e3sFBZa5SpNkxdAvyBffZsO4WgPIfYNIuyzx/7MJgPmuGTYKciGUAgh8VVs
wjiLWz1LKCUgVirie14TgDZFVGQYYPSa4qChsZ0+UuwFACdlaqqCtRnZaupNDe53HtrkgNpcxcrz
H4leIykfzHLXZgHQQKEQXFsJ+pOPzukPCgZqYlFpC1mQQJjV/SZ0Q6kfj+uHPqPYtJ2efuUSC+r3
JPHaLgdYtAhS4B/Q+9PTWCuzKE6EGRxJIdajiKsa9OzV6vJI0G++zuGdLPxSuzbEGOwxJspRSSHC
cIG4k1tf5TT2aMpjy0ernlTJtswuVh2Ou6T/GmqlTJAVyOc6vWYtCz9XhQKqXLnxTu453JLetccL
5dx/XYXItvzjJ4C87Pwqfu9XnyYcO7Fq50k81MYvPINlLK92h5H2WjEk01wc5rzgMOFVPvEwFsaJ
z7lGwchXoKAH+JY6Qjjdt4Fct073pI6Ym9rADnOlAaTFmfbdvuD6242DaoxzOGNGrPyXKs43B9sD
eDjUM2j8F5AuUf9+sSIhy1qzvmZoD5f3xyvf1UpZqk/nUX4UYXhwCQhEKK03zXP6TYVLx2DaGzZt
UuATsG9AoRWewfz93Rc31eXWODnYZRpwg4D9Jt22+c0snjhabTN0Me++b+mCBxs6mFsHHilPlnOC
PO+AOHJ/FivrXx+1SxKDe9fmF3yi/qQPYURbdtVNbl+EsczKz7Qn4i8bv98KI5a+6TP3BYyTs7aU
b+VL3XZvwGHHb264NfF8q+XPV5gLrUR6gNH3NtW2WmDyjor3jEs/5ZynmDJLpglB1+twC0CnK5Ha
aY0BRGhC0OnVT9cXyJypqbULaqWyHMhf7OPa6Sc2UErNB16jJgG8ks6Ed1EzIIcHn1FNc9CUxOw+
2Y1xBAPEXhWN34FEKuDC1r7BnahgcqX7pbjjfhKGRq57KRgFAV4LWa0waAplCFXtzNr7dmpdaRxB
mQT/ye05V7fN6pzAIM4wlewliApCD3WZW+vCiugUbtDYsqFmcq7wyIioWpCigRCQOqH3qZ92Vpe6
pBn6Sqab1TACdRrQOraA8TIpev3TLaolOMgI49ykhnxFPDMdWvsLkDlfzsGbC7048O2mRsb0Wpaw
sLWq0V34zA744bClwJPQhbwDpNl+AXzcDsbitYCqrTgZZiHtqbkzIaf+4caIEanBLmMOjPw9kQWz
2PcYuCHVDqhh+SUrYrwckMN0rj0gl7q9RBFfz0GZpG6WeozI44iiJJnNOo35MtgaqbR/1/FkdMCP
1XgfLQ24jdshEm9GP46PM6lhIkY5PPzvuUO+ddILNPdydaZd2GrG2BYYsagd4w7oyNmnKjSk8Ljk
IXjciQfBtedm5NGSC0TeQbwtVnA3X9IZulcVGDs5mXFlsDmyDp9qeLWO5Cc5+yBEANhcMmQvdL13
iFrLC1wETW/br62f4/LdkKGaMwNPSRufzsLnXf2DjKmCK+8sLO+v9JidtUZQ8VC6JZKuv7BY+6kR
rQyQt75UzGG6OJ7vG0e0/OCaTonRUlmD7TQnO7PEzFibIC59hgAasGVwHnvP7OovP/5aVfu58KsA
L6ivqIkdjw0BkQ2HG0eia1JCG5F090GfF4liU68QbQkaqYWzoRHqJ0QHRzH9Q7OhaCaPgQOWhSNH
ftyE3DnMzsD70Mh5KjJs0/4jrruoUopw2IbEVYKY3PnfYXjQwC4+8IiVLL08a84lqa8XleE0ue7C
ZrYlMWj6c6u9+RMaMxlMD1cQ+ZDNccjV5AfOZXJ30rtDQ3pUQWdcBaxkLocXQoeNHStFVNIoTiAo
3hftav89RNyuCT05DIlym1Wi1Q4IHL1ABizMI69a/SYlUsvS5+ZgjQQUwvByVo+tYes2Gk7ZbfjP
kLHoxefJlxwfbEI6yuQ2MUmG2KcmmnV6U0r+N5ZSohEfR5e/WQr6XbhDCpSOYS+rDM8XYADomZV5
2N1Ssy7EYBN8Ma1XufZVFDkptuIukJZt551fyr/qdgI3YG5uwPiDZ3C1j5QGWj5QFxEuzU0ycOfO
75rFqiCeelVaElUcTLBD7ARbLrpLZKageoXSMo9PWhDWCp2bxSLseu0VgPAuCFan72IU4DxiJRki
jrJTUp7AZUXhaKO36RwU1i9VI3AmwPt/9LnFwsQRd9ykWQkvt5qESVAyOo0rsN4krxVyQLGlejGQ
ytw7zzrw+dtBTxkwqZUgFm29U/up/XENu7d0eFjBIlVnftewPcD1ctdOXlu5/ntg6XakM6MBFSwU
mmNpfJ2c5AgsCUXR4fuECfIvOFLpn3cfjJuLeO5zaAvVyk5OuVR+B23saxxA9l5ndRkCpysYdvm4
wy8eJaKHLz2YYImXutGYzl2aOrunzJs7WpQf1HEvTapwB505eeuvGtmcuHvWbDVSQGpOWa6xAHb/
jAsUlS3O2q7QXcSgygX1UvIQPUAAwYuxXUsYMbJJ5T+GX7DZ0+kQYn22HId6BkMoCQPNne7Wt6Rm
yMYbDQjjrnQlpLqelOh6JGBddjzMZNMZwM3ubo64rpAAboecfaXK/ud5N2AqPxiWVam2B4lEgaHY
5sciktAtKAvNV15Q1jq4yMvhD1Xlo2SWhFRRR1WidyW2jth8NAVCCc13P7raJxZnUSWTslP8jrwG
WHn/kxjcrrHUiBJnq+DiTFT76Y1UUVxZDM/pnjB/AE5XErSxB64C2Agx7fD5sygx/zXnyYRCp40O
Qe6A2CwWOYaDOLZHSc2KxCm9IMB7jA98pVIFARa//te97EUITIG+nzWls0PldZERf6iEr/3ursh9
oTCC6RrznJVchitdAIiQx1evy0rLr6rj+gvhF693IjCI9HcGhrpc7/1xcEs6yJNse/MTFtca5L2A
KYfXRezmH9flOMAAbzlF7b4f33SJ9KPdzC448AJAayYMf7l5gLmWmUdxPPUzVy0HIoK4YPxlkMWt
5/hFojBg/79FYsBwmyULoL5HyKVx3R0aFBirLrH8hpWhPre34bPKYpeb3QseR6+KrXt8GwGexGNI
yYi2X1HzX9MOD3tFDbCWxGkp/ichBgLdbDFj2l3P5G5ziKCYo8mic4hOrCDoO8rm4ogq/WYknlxx
UbUEcoa4ravoTUUhKT6kcxV/+5ggIRScN8L7mM199JdSUVPPghBvgyxxiD+AMsH2xzm3qsK+P54j
PQU0jM1fkRNgIy2bBuM7z7xgryKsrUKD3t/e1218h6ldRpXm4VoJ32S4b6N3wPSFbVX/dBqyLDLO
Lvug0/FGIhmwTBgqdUxh7HaI3Q1RpNTQf3+h7b7zUwWvddV4veqjMzUnWD6BjoJH1t12GNdvNku5
b7PFRhRnYkxZua5amot0sGEzdPv/Ta9mUfpAd/CUa6vWudgvUuWQ0yKVCWmAN0krgFIc2GdsV4oK
wZPin00Vk0eYAIFSXyn+T0CZibeZ49fiSOgjQE7v2V2z1QH4O03x8RmOSz2gQGnCTkN8g/2NheqT
MAnVprYK3dH1kawQL4QTNM3KrGl4eOoeYKBlaVMVQNsFOtMcP1j43S5LLNFx72Rwf/0l/BHcj9EB
VhV6g/zIBNCEn3qtV/v6veH1lrGQ7nHH+nMheKcGq8lEWYJxTK4k/M4OasQaUJmKDqEygVKzwCFV
Py9Oox15qB+sZifxaxgfTSB45lQzesNM8zVbJJHa0LDN4bF+SCeOw4h73ES5bRSE0PCOxZrYaQW/
mP4G1CVKyLXj9mw+TQYhbABuuQx8n1hHrwa2rBTobwZrsqirppiaE4iA8HF8dSaJ2I9+itDbaxWp
7l7qeWt6XGXSNSeKIIFtBnwzdm8HrAvUu8wV+H7cOiT8lF0VAjJfixH4ZwiQCFg5EZ1HB749M8hH
JSpTVs15/Ic8a+eHFF6UI+i6HZZP4lK+cl7LIYQKoX9jDqlPgFAhiWQm/vNA0OpsbRv70P8Z4ZYE
r3EKP1oO3zoiPUb53CNC5VrqKIfB298qCpCaD1kijoIyI9WXQwg6NnuztpzTIhwkYOIGc75vJRvp
pwuRju62PuL5EoGq9QoU7tUo2uLH4mqtvIKwFUi68WH4CshQgVHxYu2h0fO7pT7YtpJt7RWglHNy
YjlH7+TSNngciWxTDeDuj1CTyE9kMMrIp+F/zRkUq/efSjT+fcTELv+xCnUV2u0IQidln/eppRia
MXjUgRueogcIkNaf4tSFOwPx76vdq5FEA94JiiB+EnHtNfhMNstc5LWS1+TVICplLuBcWWtK8Pis
nQgaqkbW2Ql/e0yO5/FY6C8GmgLdmvahz0fmWs7Xf79xUaKGggv8FRzYO/uFfoku771peCGe3WpM
JAj20Nx6tldQU/BggDimvHPWxaMcXYI9KmIGJVgMapI0H6bWmtDUUn6z5dzgR6LJxcvhXTygOa8l
g76G9Gu9Nj0mReyhHha0Ac2vsQdIosGk/rAtaSFUU3jC3KqK4ovcu2nyeUieyTY7M5eqae4Tuv5V
H7A9Z9RRHeqkLsSAeZF++aacggSHvBQ8ZsaniIQDTMIrNKXXRYiB9gIZAVUDl6lbEAbgwU+G10Df
CFrkxJLdqcdRTgUbbb3agGuMC05VZ4grFC6TaK9YCYSHiel4OTENIp/Hl1u1nx3FUWfzhiU0TfPm
PyL5xNEYPnj5MZ5Z9a7fOUNzpBI9Q3er30vs1w57QUWVknN4nBQr5ULWavYFMsNJj1/LZnH1SIVq
0OYxDhMsZsrGl3H//IYj7j+x06LzZU8cEz4+woD5Gcws/GYd73VKbcN1fcu2RAGkWdmTIAZPuOuJ
jaefwnTHKvqdcyBWIHcgzYZM7YdvN08n5yvZZYvEWdxw0+0Xt4QpwwCeQnXRIKImILnowzoXbdZX
foAWiuH9DnDF0i01B/pgDq/GbgIKGHqQ0YIC4vqZtpqMyiq3lgBagYiXlG664Pra/nlUo//vCrir
6xyUWmdo9far2ri6jBzXtpXszq3UhlEUQ72JuhlMFj8S3OMuE5cP9+rtytBAxsKRzO1a+9GVDYHV
7aYmdATIVOKIFwQcDYO5/SnAGjkRNCAin/ohOFJpoqL3TGcga5a08JdoIXboXm0g/7CPA/ISyWVc
/CdFh8VvHndnNMbHRWRY0kKzlFUU2/9BAOJZcwLq3bCj/FECvlzrd5jwxDTmmtohYwBAd8l6kTSf
pHyba/N+KqXLATD29qYYsvUbC58NgMB727AwCBF346lEczv2+t1vEHsBU2bk9eZ35oeT02OJzXZA
6zw02oee/CekwhB154y3x8fm2BcKkXF+AEyW2v1MkPT8AAB91dpZbe6DZY/9iboO4Up0hepkGUu9
OA0j0f4yFkzaOHdgBZyW0vkc+fxje8j7tnJFZTg8nrQeMzTuKmBcdZOJ45pYw5qaNEHu0J9l6Yw2
EbzPgijKgA/29VDkfK8i7f1n6cBOskNoHiwvU6k1NQqNY5yJAqmgcNNvI1raw+EjWFEy/zkcXIWq
UO9G3p2JUansyTVfdhRSIGee8ohQtrcRHwow9lcqQrKqzxuru76E1zN8U4T84F+0GQQFhqVcGlxX
qHgdz23NxVta287guBWYHwx5Dd/vFeB6MSDvKc5LMyirrAV/tkEPN0ZR4b6WNZCrcEet2jQnn7LB
R8y0A6UmHx5jIYmev7QvEXEEYEdbRm7rfjwm5tHBJVC1bqL2RKtsEyo2wymR6i8OgpuJ82lv8Yrx
YDgWD/via9LVpV6TbQvVtXG7x7Wo8SrSHcAMOVfgFiKrS9CKCRWROljOEsWO465Fvq7KoRz97/dF
s2ajiBs/ToL8cjacvvoynjPQb3kVf/oeFfi5dVOXULLun+FhMV2FpYkzGpM+0PxCDQLXuRO71uuA
hJEGxrMH+6RvxymtPbWXrFNGnOLuQG4tvtfe/+K9xT4jfJwNYuNhTs6rOWz9M/im/iykzyjmVtJR
r8Aau9feHXhgz3UrsjZLbGj1POlib6lRFupWk/hda/mhM071CuGtOLwfg1Ocv4wXZ8Jec21eBz9n
Rv3J7C5Vup7zn5t+0p3if7uSuUB4LTdMIBhh5gdQGya7LFUky8AF7cN6diIaEpqk/sdheSyBpDAt
OfFOvw4ivT0NNP0h8wQ+Tgo7xZlo4VVkrxVIkpD18GqngTLmtfx/qoxsBM/Gy2mx5AUXrZGXE36G
pJX6LBhOp4i+9zC286GH+wE5zjvQvzLzSNWWMINcHizacFdLQ+p5Xntu2W7hZyg7Vpg2P5eNc6WZ
riYUpcVAaBNIfxO2kKjQZO+Lom/GjZohS0ZqN9gmPWwrKqyEqpu++24PopkprwmGAMIOC4F1RXRN
OUzcjNE/x1ka2NH+bq/ViDlcsY7OmEsX4BDENd4xbL4KzhCp9KCqELTN7BJZWofSrnZ0u+G6BFox
ah7Exwi3son1Fzyx4XKOkTtlFIHQ78lhKg7Ap50RhFptQRbk8vriHmyF5wDZBmBeGwwI+PpZmQ7H
UYJZBDo7F19BWZQ+IHVx1DWaWBANH0s9Y+3fj618H/Bcn5Gofm61iq08v8bhfxbURuzen8j39bsK
smrpEZ7YV2mBAH6J5n26IfWrJEj+a1ECtnv5dN4c5iDYif+Eud2r1uRn7ugtJcLdjDBM3mD/yfoV
YmIqKEdotcnHhsNBVGIkEwUfg8TVqo85zB7IueXfDf2Vfjq50pd/REK+ZpZ9W+lbSyJJz6AGpjvR
Xs2f318E1plhIL/cPOz0bgw/09K0aG06j9ZJl+OF171r4F4H88OowvLQWzHjnBGVsaY0SY2zeAST
na1/ZH81TOyIkmAmDm9afNaB5L3FtEiPgWNmZGHjqsS6Ubb643imnq/HP54bl6DbYgbv6/azpyj9
chW2KjMbHyDWMGUEwbXPgji9pwLzqjdHPTgBNMMXq5tw47w1Pw4/CfTw35zkykbNbf2eJl1Oky+x
tMz6UgYD+CasEHRD0KTE14TiYB5Mhd8rolk4J+7CRbygiVsYjaRsqIQoTIwsRM8ifuDOHf0MaT+E
o4VkUbdOj8AoBVaHZHWLrSpJr8IBuxbEKydEfjvj6cTiqhYzNdevIlvOoFcZmyF5AvesUDbmHKlP
eFK+FjBi17ooDcsr0fvpP5Bk01PyoXZNuvaZ7nXJGnZlpqu62zmX6Gy3/gXB68wlTaDS04FpVLyz
f7JhxyNLHgO/TLTmlj0pe45OBTW7rExIbLRMovzijt7uGj15poAAK3IJgJfOBVXlcVEUGZ2FSLOZ
8eCZug4PGIqpeC34QmrU1M1z3OPZnjChk17yyrigc3bs3lDjLDJxciOBMwtk+qwhnYQuixm+G+IU
3Dxj4LOs3qN99dMKZaAPyrrsMLh+pP3dgrIaZH52h5qj46RhshYQaAMxOa0RUD8QUUHEthMoKkjV
/CX+s8lRBK4YNouCwIUfeTUZ+48Vu/ktPO4VqFLqiebawPKIgN2wgCFquo8ob2VEyChY9BIHC9/a
xQKwXkGCBZenOu+2MqXUaeP0r/2l0Yg9vvD9Qw/GnjPB2JDCYXa9yA+88PYzgxzjOOjt0jpWsLdg
bFJxdI4f8Pib0QPQGmpNP29C68u5vVRa7bsqsa/YTVjkgaP9Pe7woIMsqHIcBkgqOKTkp0ZsaJYm
F3lmUQGg7I5ErUxmzYheVQ42h1qunWKmaPvbpn0a6vV6m5b5KTufYHlGIkHkYNDXJT2+4CuFG8A1
uXVgz5DHxnz9KX3SLOWuQNZ7nHy426If25xRWtl7Ntnj+9xaXg1PQ9X5gpHD+sKzRf4a4Rertth8
jDgWCQlMf6FDyFwEstYczT2gyHc96wE+5D/exBYgSbudVLhHZcrP5p9l4qaaW6quq+bk5bDYFzRi
eC88n92bgTTA+X7F8U2bYys9U+HNXiuh2n/DE1t2SwaqfrhVKa9y5qK4HCSa3H14yhuCWSSSZ3tC
Os8Qbqd+5NGtlIrrj/wmmqbkOfH0fOHdwoAxGgofmIiKBYPggv8jCQkIi/h7xk+3Bits3G6gfzlv
9uPjlRqFKOdCOB9GhSwCMubq9sYXbAYeMDkIrYyUZepG8JYCIUrYZPGhM08WC3ItgSvGqie6S5e5
WHYv4uCzrKKattcXAr2Goddfk+sAVEqgzDgQnoth9n4Y6ozxOKQRT8KwHonTXZBCCErKq6FqNd1x
Aoz/teWpwaYl39NK68Nij948Sc9R2FGjQ1AZVQ0gtVzUr8cBxGSbETJpA2kLWTVDujzyHQ2DF1OZ
/Z4ssDIcMu4gJANefFtgO6yx1cyXReEUReEdx+Xb2fcl8T1YhkVJUWm53IwHyyLvWj8n5dag8DIR
4BdRXGOcQt8hxs+i5GI26WFUG2JgZNBLTMXuN4LMNDcWcoETtxboYqWkRlEkEQ5CBrHJ69vNAAd9
aXi6qmEJNVm3XoL8OdBddXIYvTelA+4MQF8G/m51yS0DBsNTW41g9VWAIRVkD4iJ+K9tsminW9eL
M++ZDY0pd5kYHnvE0GcGMqTv0g/RAe0jpIFJyRdEdfj4NyQXmTKhinEn+E9+CbX4BLJWWSHm5qAW
CWh2xlFRLGx4Amcvl9MWiJqVj4/orw/4/G1tcjZfrnS7MlRG4j+BW2YBu+dbXUlxH0kaVlYTwC/J
GtRq0LsrqYv6SOJ1AHdSG7Cz6qOPBzk8+MJ7phLu27rwQ159trOd0SSB3TqJeO7Ulzkhzzi1NorA
Tnxigy3wJaQziOO1+Z9CZvIb9Ykw3TnXV6id7EJZ09GQCvra+NlwJP8NZ5Ggkoe1/VzCCoI17cAx
kIw7OVrleU6UFK8zkYtrxSTSaU8N9PWdmXIiZjVqvVAvmHK/hkj2UPp5h8YWQdcXwr273YTjZBYA
ZnZk8nZH7gQv/cTOX4vDD6ek3YjtyyVpeXB9304kL/z1fyhy+69ojCTbg5UAoVHOAWF49h6Ns1BV
3EiGGo1uC35nzTmBaYbttnFLcdmx6zouftLWbCkytMawCnfUe+wXHAGaSo+NU6b4xcPZP6PPxsH1
Woi2GWMMtlhyhVaIuC/Gn8kdyMc/LGqhl0B9mscrO7bKy5kmV47aGrqqRnZIqIiF+i4ZMl6XuFof
USYwtJsUavY7hAAPy6j2QB1l35BMAFLqsKLIm7W3lmzCjBlrRn9EEIERnhFZji5CCfTCbZ5lYlzK
u1Ge32qPAtLYGU912Os5G3e8FAZXMYnuFKjRptsZxEHnv5HzmXXhpkq44XnJJBtre3QXZVA43ZZb
owii3MBEiWtlESXgjzKgqI7jDXopR4NbEk+KMGudghEifbYvt5HdHa71vSXGhZUqSsQAopFI1i5p
njwe2ek4PWlJs7FYpH0YcWxs1tqgAfSYjya5QBnSvnV+q0y9wYwB0T4KAnQm7dTiaz4kj5npTWef
Y9mzUjmE8No09TUc9KmwEMfs2oAhXAP/Txg2if8vvSyKF3QWpu0TlBJOcy8hMUdkZ4K0J1+0toQK
4hTQxT7GBrq3tVrmVF/R2oUuo6ZapOjP2jsinTKUMdbazs44iJ46UbnnYSoB+FUQS8bqaERYXAmI
gBvqr1DjVVhEnHbpj3liA1RWzgozZk0REwlf6Z2vklRCadUGyB6y1x+OYGetUc2dH+C/wST4mXk4
38JB4jrgzEvdYI6HApV6yaWYtPwOKWAyeb8Y5PXT/2+vSomZHQq243x60ECQaR2SsGCKyR45d7Uy
IBrVngBgyEPlt4WTgCSOCv2hTq2uyPJGK6jMh6DeGZ1Ogda+ajJVxiXQcBxi6DEuZxCZTZScn+J/
4E7tzful0ryfZ5JFKj8yMIxpgK0stGqqZfGsQlIEHaPCKDeq6X+Gdx2BrTWMS7tsdcdT4g+KTR3w
m+OEqs5Cw2mwJI2iTykGFPpblQxtQSVHvKtCDevzwDoCJ/ENIIkmU1wMZzkxnobZnCpBaY/XlYnW
8JhNQW2CFNR52271S0cLLrGwEkPX/lNOHj4YMJft7yjR5HMU3Vg71dBYPCv1ALT9WsT7oWGMrZgj
JXCdEchtyuvslP/ks9Kdw3XBlgsFTrrU4F3N3fD7vHKNeDlDy8KAYHYYGDMIIENeMawb7HLJqTFN
z4OAAKlaLbbKlG7QE9/AKTsPa0i25XJLP7jbBkZhACIbuAhdjHDJtYrp8hxiqUjpx6VNeoLSnt9c
JeQgLY+EXd/O530sKocLpqgz6eUVJfe/nrPucrLWbvtWa7a4PVznJpgk4YE/EihKncj/rQjc49yg
Vbp/C5M5DweMQr30jVK+08xhYwuR5sBhNSi0cio+6cYj5W0/+OedzsxnzQf8fD03EGmlez7EfAlk
OyUIQ210XwkVaEx9ME1Ws2nbQ/FY7Jp3AYf2aJBna3SMAtR+Z3oQYOboqanYcM/nO2INNvEhg3Bz
9VnSADhYqykQgg+YFRxVhWy7j5YJtdivy7bv2LbigbiA9oavl6NIXvQ7SaBNB6aqoESb8VdBuDOS
vLdW1t0sZaYqgiiapiaBJMysRnvfCl+7UsOzWe03tlAtAaYtAxHOUjGrtGA+f/+YYquLkEZqBYBg
aq2mJMofc9woadXBBmr3EdXwinurKu7IWbI5NZFkDXK4iQfqrplT3+Z8HQkhcOrFTDdg6UnLAzAM
JiVb1fqfWKsmYnHH3mT9Q42Riw49hD02Y7i9j27eJwRI8YRWW90WKhO4gcuqZEG+emeJUcA+1xtx
jbhF/p4XyZlQUJFmBMk0mvZfc6nPVZ3446EEx4PUnUytBSbAQek/6xSA3lV9VOGFmaXji4073zVX
1gY1fEK/nH8AgbWEIV09uUylrHry1qhabPXQy1qmmpfQW1U6CASathLp0VUXasKvs1Pv9JqC8eqO
GjiXRFAlo6IzPm2d4RhxL8R9uaAN0Ouhkc3Aaa4o2J4uxXwui3Wa4X6EhATV4co6uRjrrZrZi76x
XB35WElXfuw/wXgH1HEaHPVQvpluIxs427w+IvIwiaPSi/e/zl195+Ov0/46+wgWsnADz6mXlGRI
ji1hFLGZZYSHxpdMbMgb+GUfVSc+qpo2NSA0enWo2+dNIZgZhmtemmmb+cFANHD/5atUANDcIL5p
LluPApgO3/u9qkU3+clwI5u2l4+WviT033Ws6qhieuHkhTNWayzXzZVy/EbrSxWxCK4hnqvHzQDB
ZywwSMgdNJqObFQBboZiEemOFJ7rvyqwuuD9CmVBTyJRLK8oWoMNUy6ZlR92Tvi+fK7wjhKXV6GA
t0Dw26H55JsOce010yUXi8TAn+0/6/1Hy78oNYAbcn8A9EY4OeAMzWQxRCsw+UFvKQEnhv9kYoFx
XSOu7wNcHD+59DH3UzgWL+QPFG3bfBq5yYqiZxjaKzOtEisHmly/XU52lYDIT/oRa3J9JkCtjJwm
KcJ83CMFqahsPA7N8HNSrRpO7ERrrR5Uq2StHiC3HmO7WK933/Vi1fk8h6fakIcxjIZXtA5RwPlZ
9Udd5WT2+MoGtHvyy76QZqimlga6J7urPPzd8x4KYgcG0fUy/SMpxmQ/bJo+TvElEoeLW7RhhqsN
LVFNav2dORGfrEzGwEwZ9f+/blM0U68LUL6yVJ5uJhJUlnFf61hAT2gf1Qa/hdPIENCQRpR0XFxq
srZUJ/W3j5DIdghzr5+GKKYLmjwd8CaeTqK6V/IUD6kLynj48coIZv19ePT2ZPI3FjWK7W3/pOTp
RIThEbRQgggxvgrpisdTs+Mc1MJaFjzpx9ApAkq1fHKgZq5IsBRr+Ch01drMqrBybe41849H9h4D
ZqSpsffQK2TQJDrvPYV4jrpzq+F5fu97fanhXP2S18461jphHuppwST7lIJAW7qfPHLBXRbDmELN
ed2OB8WNtTJS76mCkJn+jRkA95XTGgEd4bIesPtwq4wvT9NwvbXj6tjX7YXI4k/EGds6YuprARv2
QUxsSYAm6ZJYF0JphPhBD7WJSSvKf0xnMFLmj8igalbcMSS3HzyeeAiCHZ+L6YQ9p/BSD6fsLFRk
Q5y0GrBWkxbZ2bfcaDpq/p7Fhk+zp2xponxFohH32R9DU8hknN635GM59kO5lJHNCQ440g2e4Q0C
iLBnylgdiUzDP9u59UTfjVDxuD0n/SvgQWGpn3ttriKirLpLROqt+L4P0h8BO4rqhaI8TA5UE3UB
Tu+d41Co9DPSi7K2gwcwNuIp9gHLGWLbs9n82/PjxXsZBkHoCdIU6X+xhLPRsLMFaKLRYqaf/Img
7iHX8Jd1zIwlmEIzXtFkEPAyJMzjsWrByHnDxXKBNTH3zw7rnDkiLcfIeJrnQhOJvOWwvLS/A5uS
R7yM/IMshfdAjW7sV2xR/m85s/6z4ZGuDuIyu+3uYC0BL9oFEty43YrwLW7eEzDlh/REr3CCkGmz
lPj7yY/xugZtBl/cUGlb0d0pg+2RziZJBkM3X6kHYnY5/MRR9xPnDRhToZmHpjLddRnTqc5tcNtv
vMt1dq1d8iQlaMOAhVYwxfkmuznSU6jO+cvOgDyKaBQ+ho5XGvNW9IeRk/wv4Nen24Dk+zdViE+R
3JlDfD+ZdHFIrI98hqufrORszxh1TA4hMOyicAadGmHW1C0UF/qTsKO6fTJQHi4F/EAOCYLc0c77
Dg8FIcz7Pv4QgxsDpHii/LCciv3eJMW/jzEaIKTYKebyKC8NmsZvuJEHuYQsS+wwfdvZOZY0IUHN
gBIJdhY5XoOSZr1UATrds5uus3hgseFLqP93NM8gnL9Z+93LthEvm01vC2yyDd6T9jR8Onc0xVTa
gt7xkctOPERJjjBtPJRGDKlQyJJipw7/LbU1i3ge3Woj4rRk36gULvBygpcsHDhGr/a0JC6xtDib
JFDC82DHOvt468xHhthejAGP8GOWjXHZKANac2MpDCqnfWK3OQNzKXGw3lPfUKNV+RgenM5yLwPg
4K1hOCKLnt5wZ/8+ESzsDaOawQW84B/3JjzGhaUDbo5jYZQUIX+hdFZomDsFBKdk5h7h7HUbH8Tb
Xd1ZRx1sPolgChW3v5IWWhj9FhHDnSVElDPJDLTdZ68j6lZGa0XNTvIOX+e7i4xB15ryT0/qG+JC
gQ6F5JTGZhiZkjo2LJnOzf1AwysQ4DQ9D9iXj2AhHHsL5XeSpiFRE7lx+kRJ/hMfqSx5Al57Jv+d
KuscyoxG3wjlCF8CBvnklpbjQoAfZ/LAwlCKUxgWeGRcL6o7BmlAv0GMr/pbAw3W3V2G/S+TBOgK
Lsdsl4J9kURRAl+l3e8/hmw5puhOuSRD+1UqBJN7dly42mZe/o6Ksny2Ue1YlReq7eNsEex9IXyE
A4z9QM+kN9Lvda3IHFNM6dKfkd1P9JLl/lH5IsgMTlPuI04lsbD7qz/0r6pfOOCKCczYXWTe4dHz
GebGqb1WorTX/vjHJ8Ery5mHydP+HEZfbMWl/rr0jTXTUN6rTwFS7Bmy1olU4Ts/RsDH63wweBZs
UW6Pheu+URKPiUzcEzhTXf1YIz2woI0rz18hJzC9TfNNhkmrHSYTl8FBrpF1fwk+J8WEMvelFRzn
O/2Sey25h5wLgpul2n0+kTX7TsLjNRZAfB+jqGpg31O7GYKAxh1G0sS/UDK5DLorqMMDa8ucuxzA
aKA9ED7d1JNtrl2UUtD7zJUZxjiSCndXe8CFcT7c2Hd5F+8I36L4OBU1oPSyBnkLPTgV21/4AKs/
VxLC9ceVQmXVeGjhb0QgKNkyI8XalLBOgn8DBbwKVMYv09raXXhx/yqtHXE5+BCrSn8hsP4v6Y/I
vmrMwzItQuzARbsVP9+D2vUsZjteIm3FPQmrU/mTVVBDwBGc8+/NX3PFwaNoTTpMsKyUNzA6hjOR
UFaeEYvHYNTkU998RTlCIat20NYkyqL/lMwDTKgeY9orGSyP6tFRBBMgSzYGCSbKzNjLYYxbsbLm
VQ9IvLMgSItceiLZG3/4kWJ+Bp+ns7czSfuqxrvABhNlund6s1b9GLQZ0EZ2Tafp8w8GoEorZqX3
S6RdQaaOr0YdgPHksqsCUFwixS5Tu6JAu1Ny6nq+tqm+ZwcJc93RlnuYnyc6RCphEX6slnTIHydt
qnPdCeklnF4yLfj9FJhXaHvrnnTPFNYMdHYPfW8sPrilF4qpMDMqeCAHhwwKpgYX/Q2DiJ4u4Brt
+utgj6iCO0AWyrgQ1sH7tn0P3nhSVgQWjnmQMjzEw986DoYDB7D52bVt83BAuhkmcdNIxzljXVz+
KWgmdXQgXA7HL6lyiuXBKXsoAk3Kbt0LZ/NXknAtW8ysfV8dtA/wOZODJyiAopmVb/9y4XGVBw6B
nE8WEK+8/JfJHVOY/BKQ3RsYrE90HOHy/2zdYaGLhB4xZ36VBnksDYfwwXSy//FY+TI2W64QsSNE
VkyHuVLeTQH0PTg2DHQq4AvLvk0LTcNvS/4BYIBjmSL7wf+V822AJW/qPkcAyMTmqoafA+wdWs06
ey4onFbz3Rn/0KxSkxmd/Y51VKoHQvGXzvOgXV5w7LNiK8xDpT2HEMz1LzcaVPBdc5nPcRnstdLa
IObbnDFGcl3GmaEMIsN7AasQvtk9aWTHmXNIb00XICCE3WyD+c/+sn9DZglhdEYiiIJC0cUgNwRX
mnfO8agt+aHeXDmJKKQk8wZRNsCZzEQjx64TKlp/nV4AXZzVYAwRJocucVVL4n/9Z6P8nXtC4rw/
Kn51ZJEJ4FeJ2D6rnTre3gUNF93ik9oiVGYfE+lkyNMFBClfU23wSxEvFUC1iNEfI1ENc8tKQiKI
TVpjAhQgl+R363/KXVhC9whIVHlSrJKuqJlyntpbl+lblopzWWTMIem+gU5uKsV44wFiiCXWzhHd
YiSjKmSDabfJW9na6j3PzUkNJYP3ISDwqkrXi9Vhz9WMt+3WGcmp/Ar9LU3Txp8OY9xChoJkGOcb
PQDmAdDKN4yBIe8KGBc7rgOsKiFjmgcVtladjjREXcSKAuiJDoRXkr5AgsVJD7ibkV8GQy/ZMnfj
SdauQlSx5Wu3IUzT70Jc3djpOKVRvdxdXX7qdMwMG9iSxNruq7GUcL/ptDkL4YaOiExDdADd4MvH
NOTt6W3J1TUHtQez4C5NT6X5h9LBu9j0jAXVP7cHLzQE55OGb+OMuQYMMml4c1OsR9VGKvOwBZS3
siRKv4QgWj6QSI9tDAtFNUADwHRdol8d21dSZ/VqJ8YdRX16gY2KCrP0kLS8+WTyYHJQZqA1YOUy
ek9VMKnAyDItlUlQG+Zp7Ye1xVZnbnhxqYKpGy5evWGVTKOuAbdnOMymGP7Z0rsE/zURAGwhSelU
G/FoSdEc4ucRfs5h5Qcc11LeN9yT6m9dVCZJ9D8G24I3DVmHld5RYWdl8IWCAoQ8VdEM5stpgqu0
H6KOP4F32Rebt/YGLfEueEiVbBRlBOY9TwvQvJTwd32jucl42GRqi6DbWcZSYtmkw+fLt4AleOhb
5MrpvR22qCp5jwkzmiXEi0mmfzA9i8P4WZtroIWr9wFz2WRn6k8GQHJjPeID/6YHZa8jZ28VjFK8
NZGWHIg+Tpi6FfCliJEb3GSL9uz2aFXK+V824T0plHezrVLKlZJBf7BGbZrnIKoqoHj+8ERhnwmE
Ntd2Ii/MOaP7rw5Y5Y9XW/NBfyGgdRTspw2ic98RNm7a26hcHoWQEUg8vn/c1MikkdxF4MdB4c/X
eKg9wq7kumMJWk6PwDQDVlldFWwDxrBy1PsS5qkLFqax/NEOapz+RFdLLsuDmSLg1DxAUNCJRDRE
49c+xvuv7shNPq9vdfnP9/20dA8goxUGq8xt9xTsx+isxPh4M8iiWRc8fQPWG0CNMy2fBqRimoi1
2LGubpKGe2Ew5hOfiITng7WDPkf2IaltMc1Pq8D91Gn8BFt4MgN849mB/KNywQnZxiYdXKzbPvsm
zr3SSbpDfNfxxe0LGL51ae7H/Ef6pqztwCKK80M0IPJRp5O9ZQ+bq8/rwSyJ3uFGT1CzVnCa4z2b
36OLdQvc1ynwCtY+lGE9aKbMUksLJ0jyfVtps9u8+Srxu5xtZ8saGKto8py8BBbGuRcxS5S55gwK
a0nRb0kgbemzzD3+WykILAXi5+dYiyn+/C8RS4x8XA8lMYgb/LkOEAtTXY8arHHhooY/lPBqiwnm
hiAnMpCGlbI6sVnOnW4B5gKsEcRN7vKQUf6umV+9Hzt/Tyc8z0RKfJZfuCT32jNqP9LrFCSkg3dL
lAK4bHVZH2hNT7QLbHMjrLe2CFddBEjtidu59XWfkWtgo6hG66cZyRFdiT6ffIW4rAkRmFwxrdG5
n+nfvYpbvwgwe1g/S3d+uXcTQ/YsQPpe4yXy2MzYxpXt6OE6UBoORfMF4c9d3OAWAYuA/5Ev662Y
pSFjPtJNlvzkiqiWs36fbwyUkrxNTMg16LMqcDpd+6DnOvUKvftAuKWdtowSO+EwvvWyGS1WjInS
SW20A/EfXnemxx1fGWQZ4E3V8lO8v78kBJLXGK5P0/1kqWDc5oDNoq4eQvs+fsXWB8v2WdT63t7B
nkQvSuw9Qh0ECglK7WP3e36t5R+xUM3p5GCYe72+zT1HwDfhtjUbZ26i5aDx6xtrQ2yJQ2pFNw/v
iGCsYxUZ1Khz5HGXmm0R/14KYLloyVEc4rFZhe1NQtUu4hgBimI8zxqVO8V0exUiMPhtfxbO0Vfy
CMvIGFPnnucouYDjyWf3uxnFKnjDS9/pF1LugCEU2m3sVxwJvbM4/eVcQXDr76Y5vuanx8MbiTrb
NT/VYGHTpi6ZcCqI8fGsJ+ADDcmhzwlD/SmfVRI9aXik4CgzRTMwScB0KL0bMksxQpg42VDNHaUP
6P70LRZB9rMP3ArQMppGzisjCAd/QLUn5Foldxh9UyL+LcLoHqgyoxUFl/XCVH2HiknY7Z6bXkGq
64UO/pOlbSrix7+aIijC0Y9SX36nkYwzTD37uu+g3F6hdKGUsJZGQtxFSPW6zx1XhLHpcPUdWHot
HUGlLWc49azJX+T75nc4uTERXQL/1/W3+h/EIz9P/DXBsYfr3Xag1yFmxVhKVw1VuLysK/dN3tsu
HMxiR38kupKrkDQfW8aYrFmIocdhJEovsrH+UpzQjJkNOH4k4Mh9GvyKuRyhOvJ5dtOMSnBdKUNZ
znFg+m3W9+n0QZsn9+SX43ezP6NEJAY37NfxdPe/faQsCyfga9Tcfbi2hkDjKTa9fadtRID205DC
MB8wSIACgZWHoMbOiehgSgRRl66AISX01vpshxXSYHuJnWqW29EyjBe9nLLvlfjluxrkYQc1UobA
6UR/J6oaNY3QRuHSd7CidhJWDP8YPlgo+mWv4DALDsFuiUHtfzmgFnQLjkL5RFtVHQI7o7HmPPdh
REpwsjgiaeNiiyfZDRZ7tLzd3lRRP6mDcDcaKUVNNz68BPdtv4cNDUlu1tnaW1VXcC3oASsbTl7o
2b6+vWveiVtnLPp3Eb7yFE1AsKoP0Q5cznQODx9E8qM9bBWmhMYL/cSa0rNkQtXqGVaYG1rpJh7z
lxsaGG3aYMCDs8t+BQglAOfu8CMcPPyI0kIzWov01NtFoEqYq7wF8rf+kaNwdqhZi+BjN5qhK+nE
dj+utdxq8y1YIxqUlrJD+JRM8+4R0q0ckDE+79Oe67Bnjv177hiZo8p9kshTUOWYEB96sDX1XWaE
k/ZUUZYIcYBH3DyEhCNSfqc58Z3/Ol8acowhtuFIUxRxtIXiS0iujqpJ9BtM92Qbn686QVCB1CfQ
N+ULd69Wh4v9qzeDlqqkeMcutxOyceY1wCwq/rsNZc278UN8p0q13j8mk6gk1D43Lng8WmJCm/kU
ed0/1vCi9oDAY4jLBGhBk7Eq6VrLAj1X5k7oM7A7ynrC9bqEn8ULDS28NEkwFDxoow9il8bc7aMl
NNEeHQTGycWwU6TCOjYgvYf11/1g4aeGml3uHiXNLz+ZwWesY3tjR3j9J+unVWWJb/7jWML+U2tw
W1ymzrzOxSXkKGdCXgJPzyS0PfF41oKAU6L60Ff/o/bVgGzpUGeMWcODAQLWG1W7YMxu3usBtigc
/c9uw5tCVu8FO4aotGC638CgCqeYIC0HS0e4fMeGvwIsImXniMy5n+3ZcJQC28WjbtomK26mhGkO
lDiiXp38G+ltugIpgm4/gcNZ2/9SWe+Vt4tNFCgCDUWhOBpi5Q3hy1+RS80d2BjeFhoMEXGv3UBB
cqeiPXPjVPYkRPhjGSixJIQNLEumIOlOQsKew7mMZgGaBcLuB+qCHJoIWo5CGT/YegAY+WqfRNaX
+zV1WRenRkPkaeYCH7V9armrvF4fGBeQpPVWUNMyOqM8EVEvg2Yl2UG6MuV1Agi/0oHn0HtxTMzK
1pUkNJ0kT/DobMDqjah4adpm+SLVVV/sYRWWXqpxceKrZgQ+jaasRm1OBNcIWIW3LRwnpU3YU6kn
gT2EyxnyhYurpPoyShkgUf7ABmhZ8VnB9/DkeKnFcXFZHWbeaBeyTq0wjAiolQPrbrKzj4SjlOvT
aclUd9kIOcJR5w1Al2M6m1zFFm5Nuv1R2E0yb7HPiADlyfZJIGsRe0CvBqdxtTq+NAuNxsXEA6qt
3LcRBzXsY1R3x5gLCU/WzFuJ44PKTwuUCccG+rL41iJ49i2oAzhQuPTVuU/EJyVGdyf5HNTihsc2
Vju+06RkHDnbFeYJXjUns1DUuvT+jIpaMOmByNoFbJ6BJSNzy2jOiBnPaNabF2Z3ivh1Q5Juxtkm
gV7jBFuWMRNK0z/j2gZwST+u4ClT2JbVYwiOaq3lR4b4PLh+PST7ykVOQQHJzYK4DSTKW7XFLgE3
5Kjl+ngIOKTfjGnmlSvwtHPFYsdG4P9i/LnzMZJ2l0Vzl2ELBDUkWaLUpGOBbIUqwlZM+lTcuUPV
KL4ze6wTvwekPoEgEDeQs/I07T69MBSFEUq2QToLvH4O3BySV4ivL29voXc4yAgY6P/+ZiTZmwIv
QfiNnbL5TIIy1tZLyursUPUosWGp/RtQt5HFTcpo6IVjydOutWLhlgZa4DJALq8WvrytvxOwJTLG
+SP6ZsQ9thsD3eIROe/xN3fm8FPwBj6QYcmhTmsEkHGGVM7zH9VhzXbXR/G92rmhmNf9b+mFmqq+
jcqZLuYZ3rP2s6ikYQSI2L1HAELjNLAANFwqNi7ej6QxNysp4xaTjFMTYFjGvxQQupQHldgvrEGM
wRuKwQEGCVO9g+b7z4MLpGYONwuc0cGm8nZTJfDwoPIEt2cTYK9BJDxZFuShXXfDoIB+IhX8XWuS
FFDPM84zRUAJBcLngJN+RpB6suU84lDTakCiTie940Vn3qbKqiLbvAzoMp6oxf7iGd5QKZeHQ/9M
5gEiG86L8/UDZ6QLiBn8V3d1BMXG13qiUU3jxTThzCn6C9d/boFf9fy1F1RKILF90acLJ24cQ87O
3eCR6EWprTpfmLxp8tB8DPjsrVsezRCTicqyYOiZJYxzYWsoceCRpr/2ifNjaCsq7ovtqyzlNEJq
qN5lUz4YS9U/RQqcj8YSQas/gFihFpenV7BPsBVV7QOGvcvf6EtQwIyfHZTSWev/wqgcMAnyQ5N0
mi/Af2Zc1/afK9CAy9IW1K8CxydiRyJdI3PxajJnAdXTrTTNuYci0pbVXfI+UYrimk1FtKUtaPGZ
HGsTRwP3awlt3AUvbWx2rRx5cuYLCrRhznsND7jSQyWbWhiUaNtJqYEJhuKuoa4sP0SpxNG/8Gro
k/1eILhXpP671/Un56vKA6HyVAcX9zIuHmrJbDvVPfREN7MXBgyAyChZlG5Jiw/a5xyZRyymI69l
DrwDh5hWOCsX6jAeHQ3EbWSzZQy2oTd2FtMbAqguUuSqYpr812HT/lvjXNxcHuPE54R7l3Me3EaH
ofRCYw/H2TdgETlVPasGFii0JqxCpo6Gx8X0z455Sv6PBDPgnSN4m1ySjPckArtWfRWItucrFfsB
sN/5RvdssbKCyGXQT55p7mDh5vl0Ribg8vwfRm7tWKkW6uGk5J2Qyxb+mWLbo1Fmtju7/6LKr914
FgRB27r9uKJWFoasFQUf83FxTLpL/5lyxExc1YK1gPvZtzuApeRcUXAe7IB/TADnJn1xyqfUljPP
GfIYXwsR7RByPIrI8kDXolMnZzP3AsCM96R0+x3Z/MaxOcqSklmp+HHWXk//orwACOgW6xQ5Qs84
Vlsb2PQQdYqoAD1S55VEmBZ7EPjcK556QzenG2rN5EUhU27TvU2cXu5NfquGUui4Z+T6lPitqzxr
cc35LciK6gnuymolVlY/Qj48Weh0Me+tsVMA53DPuzibxCbPdIW7twV1rEW0jtu6QXYMCjDLpd1I
GHxNIOqdh2h78kiK9zCEmQnB6t2WEW99beiHYkEq5bjIJ9raxC83Ykw4vnB/plu4p7+JmF3p/FuK
CEmTQafwLARKgMBalfza9zEpzgyaLHvM6XqxhT9j3uWp8h20rEudJYdw8m0JKJfIV1zixhM9mpcC
04Sv48oMamCjHY+UkGMxNqIhfbICq7mbI05a7zoT5CXzKfHY0eBSYaRHti3tUVNQhBk63diDRDDo
jsx88wZ4okbeT+Ad7+AFl1RqRU1MbME2zXXep4zozaqgM/vcYdglslgPjd8KN4vJC3BZXIpNwjr4
y5+GDD/dw0iFyWSN7O8MsVN3VztjJAtu1dYpESMICz82r6foNVAT9qkrCGg3CFM8Lw0HuV9BROi1
CQ9o25r6daWoUEvbA/cEM1C1zBy5BuODZMbPwLCS7PHsdboT7k3L3IcY6yCi7FSj6zHKBjawx6qf
K67HGGPPcZZGHvLHYhPMzGaKIjojmlApThMNPgJotW7samN5qJbWvG9C/fPjMJZ8pJ7tKSJHH/OE
CF61A5sZ4NPZ6RuCpq8WI8X/JTlBrUPbt9i/zPWdT7wIIQvScYivlMIDbbLKlSn3uamqn8CXN6Zb
ILhK1USrAhjt6yBsGsDLcgWaHmHAmHJzOY2VcEKP+hsxCiO2H8qnZWJ3G0mUo2ZMW6LQWbXU3ya1
+JdECDonDHkzTSBpKMotc6h4cbwx+5+bKaijx3gMt4O648wGkV6dPNlr07YodbDB3dwwTyLOsfE4
cPNdhliv8ya4a/WNj92eWHxgSCq6gklCdWIiNF+bBEQDjbs+Y32yTuchcPAVch1cu+5eNW7FS3e0
cQfYm+6eCvBHucKO4V5EpCwyM+c/1vUlLuBQxak2T16auIxHQDfoZEYPEf53t6YtvQmI9mdbBJhc
NZt0YtnIOUbpHoNPWfZKdsk+CkE9MgZARsPFsEK921w7dUmtx6O5DRriwz0OQadBLbTneMzIppYB
87z+lVfm7/HW13noufPS2I8iotv7SrNOJgwwNc/lPeQVvMETD7Cosj+C1DEMkgPGhDTwa2GpRaxg
YoU5jyYGCML023XnIteDz6KSaDS6yQ61i8gh47pJYOkDQn5eqzoQU+zoI8azlmWMAz3v4c0wCtYt
GcciG2LrPJKKP0tnLewxs0XbLKj78JNYJdefP2DjPS+Y5JGFyJZ9yB6DrvnSbeGtWiC0E5qdDf79
CsyrDHS0z+oNRqxauDWbDCWqX6R3jgFNOJcoYIamSTj4cZ2hM+RpoHUfjBjQ7geIAVdP0nKso+3+
qBSg4QKEGbVO6fIZwbeBVe0rOIaRCVJcAcYO2MkExNq9mpUld8yYs2Cg6dSiwAg/2wtCvcuzZrhQ
M5+pZ+ydyJvABjj9vkQupPgez5xHaXerX5IC1GuigduT3+dpfb+6q705qBl9EV0cDyW455irIP+w
Ys7eCdrjm2OAsCGCw9Dcw9b5S/GecReZwElU9isfSTSdXx3fbPL6XJT5kYiibcPxmM02e8k7YUF/
At1hHRjwbOGvmpKlKrOI8ZmC+ivU8aFlQp+23W9s+9S0+nBDUahsqaVWxjFJlGDEOWcrGTA3rzrw
6VAwBsQIDLeAUXFel7dDwwSpOQLF+j/l9Yr84YfNRKMlKg57cT4/Vtr3B8z+Wxvexl8ywGclKESj
35SAJzmRjTNLzARNHMi9O+C68d+o9uW847Zup+mg/7uFPHxp/1Hp1bGdpQdnPZbaof7gsCvaD7eX
SgFndYOc1OOOUuTjC1vyw45XagaC+coIJxJx2o5rSMb5I9X/GKlPi0WLcbbljWTtHQqkExMfQMxF
d2hBSP1bUYFR6qC7Z0Qrb5IbZFQ1g8vEbq2SQC51v4LIZmkhbwaLUPBA2Rq6hcF/SrRT2GvpJ8Oo
V3cJk1TxniYDTk9YAOYWlUzQ2VDv4rVe36BUFuz3NN5Rt9RVYPwbbrg66WU1kUwkNLqob9yy0SFS
GiZPftRHRZIUCNFliXGjRKNW27LpL93wVvumjlNt1GZSBejffzCqUMwBqVB65blveJLmRp8r6Fo9
LgPto1i4+q6/9Lvlg1uMIgVhNJkT2eajeeJI0DqF6m0v+pg0rSUpH0WTEZyWsMdp8hHTEGnyweiT
9bWpz1ZMggFm89WRa1m9VlWH3U3yI72fFfEGy85If6wXGJm2W+3cwFL64tCYZ9SA3y9xkThtbgrY
T0aWYeoHREDVBnzsToV7HaJZ1V4N+hgSfJUqh99VoUKUN9mw0OTuU7ma3tSTal0dyTM6fBoOms4G
SH9lKFIdTuYZfXuHOt+h733KTXgzqO9cvowRDmqjiBnVCqQPvXJkmvQSt3gANrP0vJr0YWtUALNK
AMFZg+w1567B4GcgxvrnqBFhp4pYciRMpQjJaB7OrhCUo/3ECMjJAD98zNS/4HVJdC6sYiSe2Zay
kXJ+2JUkhJzvQnp/5dP7quKKofszl/RhfDruB2Q5lN0VO7w4xLulqKsf8D9uVcaoY7djz9emsl2q
qw4nWcc4BEf0XLKD903L8WSkg1lWRQlDIfJeczgimLjUpaNAXzzddaoMagFtHTluJW1r2Kpn8RN+
SkGFNgBhlBZ4Zvc+FGcW/gn5MK2vurI/M+yrvaquCrUw8i/aw8+oy6GVvcAlAUKkSGcoE+6jkI5e
23Qv7BZcSpC+3WKyfwPSwMu/fuvFl3kucj6msGdLnnCdimwZndq0gqvEZRSuqh70dGBX9eGIziR1
GAcWunoL2IvzZWG0hBgH3+6DPQ/9YtWVRqeFHfvKhli5vxC/7qGrXcUbKODS0uDZtpFVkmnyOWh+
21bxZ770/1s5ph+NTEUhAO4cqbj+teFM6yDkKJENQFXOI3OsRA48qbgF4As5xW59fs07MXYUQywn
8VcG0F0SaBHrvMrcLn7JzbVvHvbsvRmywNlLTZbnm2Y35s4LvNccigfG6f3OZDT++kXROloMr6vS
o9SM9+C3MmrsTU1/Fe9J9evK6IndW2ddpqcu6PisUd4kCjEsbsj7YkfdB9kVzqhLJa57z5JVtpnl
v3ambZmYp+bGoApIXuRxLyZfxEsufM6uLpYeneeUc9Y3fa0NAxmprO4qr0ROhTFbGqpDGCwkdCtY
YOAb7HJA/C6meIQ0vF7V6N18t5OmOPdlabUlXPZ2MIG0PZwmcfma6n8/BaRDPBKeLilxttren+ix
/7YdFF/C8QXQG7CqizKOwpP19z+fIs160wGAWZh/B+hZ/CMSSTHUvNbyKSH0hvfQ1lQAjNP9E73A
LtsUHJcFwhAqMOwqHXU4OjyIB+dVIgfkuevwAp3gpXdzmjvpvqVoN7iSsvDGPRnPrlhQWkBBVU1U
ciCuwIuCdJPkGVJPcxfc1GWhcU7b/LTGcDJzRTQvuZi/VmsoMk6cuOszG0PSa0BHCOJzhbJIiGQw
M/4BJLdmzI0gMpzqwEVTL//J6CX4fO8W9ZXuQwzlRcWP4j1itYeSvaXhLgcf3pOONw4awxj9NnLd
GqFw+tibkNo3xUREHJqibY3rnSMNE3f7s1h8Xeqv/R5MVU3HAnNgY3KZrgLxq2k3vyLQYFuON/mr
ua8FQ6MEGEqslyyHtJUU4uedFSEOgiIPf2oa9KVVk6CFtrlVdqr6NMmt9bWrMp4bg8qUGRys0co5
QAPopluhw/U+j56ohJoa+kfyKyWT3VCpwcA5vAk6ZkoPwlntr+QmFQp7Z9zFSJAbWJoPZYgPWiMv
LGdzhHiziAR4gtQhetoPp9UjIfdYMYLvKB7vqEo9RUnUUivSCzVyYFSnSbe3QuzFiDYgYeEq5J3C
TaiePnfimmmgeSLXvTQ4NBzSY7aRLQ9cJPChDP+7XcUGJGNdlI8dnfkE/IEAO1KdcP0eg2pwg867
IqY6cWDiu/1pVfvH3VZcJ8TOrxr0He0jCIIPTCHe6WXGVaWB7Fap5LC5He9N6EmCk3K4tnkNSWQT
d9FObyrwtyw2OLyqmZIqti5SSfGTVkZRPafVSyb6WJ0FKT1flWgwnN9dj373Sq5jQJ0duQDUSqVr
8e3i8mZ/FHH5sN6yKb4gycD8DblUvCOnQrly96rLUiXmrBydYvQ2Ht6jx9S4D2D5abSKhypwx//g
v8KmqE155PRd69Rlob8iNm5X0p8PAtUPMi/d0tQzO3yCVkGksX/2+D/fxVicdZuth/QxzFSe6Xyx
LRj9o1B8E/cWXS1I/3QI13WIDdVbiZjyBoQ9LZQGCHCHA8oEtKzL8a3teH04jxdJgiYanVDZl5K+
nP2vX8zsv6u+SpgkI8HU4Ys7ECSjXrAmG9iBQUyZn+H2sOI80N6H4PP83kk9uKOGUrbJU5dkdnNI
c+fF70spdSj23RocgI/LWxSDj0ErwDtz+OKjY3DQrEMTnMp01uU3IfjaGbDd5LTou+vDdyWtTSO9
oS0xWML7SZhL4dPBh/KnJ/nVYxJrudd5E6hGvWgjQxMCjvMU2sZD/ZYy3jRuvpob4OpEIBbfrhM3
Fru0RWNhV+VsWCcZ8jSRWQKFYTtxjiHod6sst/Oc1i9tqScOwcQAcrU5AdsP3NYPjtpKnMkTJGeG
+WrIIYhaoMjU84OQuTL9u2beNE3LGuV1VD/LEbk9z5aIeTUrbqkwxY/A/yzRrp+IT38u49BkNwNU
Gir5slF2+sCNcvhguXLEirlPVRO2JNwsT7/+cvvKe647SkEcwb1d3LaoOeHXEsY9yyFcCD3Ty+PD
C+hTz/taf64Q1Umkt+0HgMORFmb5T08SkwLwE8C5ih/HQNzYXv481VhN11mk7TqOLvrTzn2Z6ExL
cCLaw4svQeEG2r66LRA+RLXOegBQyXYI+y1j9Vw0RZXRt03NNxSfVtmE/G95ygt3yXgeVO4XUffH
nK6JUuoZEKEcvsori2Ov4h87zTvUUPLs4sSddepgvMG+Nw2fFSLLedrD8iMv+eixC0ybKKOxTpiA
Avjee7P2f+FsqIaLjxsjvIj6B/eqSeNXCs0iSHS5H/UwAWGp3e0viFL265BRgrvnpN/2du9GULM0
x6+y290abo5ZVnR77a61l0uLZsF8TEgEluoObkWzSgUUVHZw8pEGdJDEac8wgoQtI//lchpQv74R
toHVeTFdiU0Mxl6Ei/P/9O4A75jlMLhy2v1cFMlr5DGJS2nB46iu4XXiUThSmnrAotTZqZiZnHvU
qBYyXIWqw6bznmEECqoPrfrzDJbgY/i6z0V6WNAjxPud6hAnngcPuyYVvhe13cOy3yH7WWdhymEo
UBiKir53npwI0UBx0/UqNLoPetY7cPdF3Tic/pkCXnQKfAZurNRwjuiNZoZxYwPg1Zu9gxhoaJ3G
NS09ETixPm0ypG7Ud2b1RY2NqmJW7bwg9SafWTqwDk6FIAC7POeeeWK5oGGAk2NhfuuSRfkaDCnR
dFm71/QqQtEcIP4eFpyiE0yxa+j7KiQGEgoEFHMszbD5n7jrKt0U7VIIevVKWKDDN0D5t41CY1Dc
t3Cb16a04TjH5MCzxxp8zgqqGABWEQV7k10wMsHNCrWFJpnzlpc41OG56QN5uDazjju7A3/iLzIp
PhumHF00mB8R8eZV/HhPWbnnXXFWXbkKe150wyuJCTqPEcRNOyXVd2e1LYkUJCppS5W/Uj/yi+S8
eTrPOsTUk2N90/5UpmTKhNcoSH9005nPhzYX+MVd4qBzHsHsDCtIy6YX1GCQ29kf/Q0lFZHNxquB
DyhZF3qhnWDZIQLzJtvx+8i0eozdKjdvsEK9NGhKJBiNAdDGe0dF9FVHUrKDmcrmvhIAI0rw3vR7
lOKSWqATtjwUguVN9GMEeM+gkcVPENKXbBWx7vVzZqq4lsOsMCpeihgdcUm425N5rbXyBdN9rW/t
nqzaUBadFf1emA4UXWPpfQ+mqma945m77y4TBv9AmAdlCBAwh6TF0hkcRlareVh8AgL/DI5iEYzj
reeYa1HHqM7xoeT/oxQCqSmRrV+u8dosYdCcoadoMpERg500/mXpAbzDaWJtgS+vxFUcNPZJzBDk
HlawJA9CEM7BDqvbyXE8t+UoVhXwxY0hIeTh3R6n1TfnN6aQrI4oBV8k/GfnJW9r2O+CbUBrYXif
rxtUy6qp5KQS7gWjOQuk2Af61nHCtC1Bozh03/UqV8XWV90/dwhfPWVe0nbFqXsJ8CmFv4m/UGUL
RAvKcHr8rPx9K86BZfPrMFgpx4nwnG0dUsnCvvSadW0V7OUB0LQDM7MNTXMmqYLtDWiNfpPA0Fc1
6/LpcWw9grWAmvg8kKc58O3svGToM5r+TTdSePb7IgQxiXFyLkkwEoDnilR1N1mXhc7kKJf78Iz+
cUngGoQYVSG1kM3p9CJB8zHn/ylKVUyi68vNc7iMmo5TenKdSDxCpcf4nPOjyjkpo74t/rFMtuvV
fxLzWHE/S8TevMLX6EnWzUug99laPVYKChBZNev83pTaV+dNchxDMMmugV/Znkf7/nieuNDiEq9F
ZYNoG2SUHTsP9hDxyJbeBFH5i7Cgca3a69qitlYAK8xjOZcJWu/GQndilzI2zRjOMn+KIWtllv//
qQTihWhgbjYXwWMqUdJS44v/jiArDpe9cNxXTUaZaq1zeDkzBq7LDSYN9LI1zAiETWcLidtBifQd
XaUHkLk0KTQHrpSfKwo9g5gjwjstyq6/qo6ciXi7EW3W6VbbtClvNZ5IRbocyIYV9Zon2xzOm444
rgse/DFeSEcuGCDQBvvVeGIQfiU4eVFjS7eeHhjQVoXuKHi5GAYvoPzuhLHkaDeGxeqwn51ae9CH
ivuWxcJw6xQmI8FREss3Yo6RcO+eU3n4nrXejtSsiVLTIipvrd7diTnuomqrOfVE3k5IfMgmuKse
AbBsoJi/QrDrkhrTO2jCi2l2uKvQaaUkk7H2ZZ/5Tt2VCFQExz43r6NzzhAOoOZZGKHnEFgv4ZJd
JfwXCqzqE0/0KvimW5F+9i5923nnh9Q3KG+pnAUi9MhK+4R44vFAbpp2YN518DpRZsnHX4hGPj1t
GsQVNryTgvWpHfh3R/k+yAAisxp7CP7gyLfL5DLHDcvfAOMkT97eWJKxoKgrg+naVhG3MJEz+7g2
+NZK8D7rOPYyy9Hp/IPgy2Kc63xsOFs2c7fNgfBQrNS84sQZU3gtMVddEFQSJtgZKN79ZSa7MGJW
fB7J1/pS/BAEImxvOKvRcZfZ5OgW1TAEUmmSnrkDxe4nXsQws2m72408PijsE4rQunTpeuzkKNyN
glRbFon6fFWoZRHSBz+Z71nkgNiCLsAE1HC44zHGRSio6svHNl6bC+dx3jv26NBIy8UYWrzG2I7/
oTQIzmJ/cSbXuRLqkga89hZzm7j1H9lGwuHC3JfGpI7k3yrwOMUh8A2Carh6P4pcY06zqUfohkL1
WAp3+bCNXomWD44uo7yshhI2mLkBHUl2iFlBfr66QgHktlQIrgm227CxJhe/EjVsPWvPF+6o9M8a
ir6VDHCJFAoX0WcuVC28iUX6OWJnt5k6SpNRnrm2Z0WvgpkqqYxOmVKBbA9Fcj7vIFbJnnmIw0dI
N1KykKz5XSrMLRpWj+W1b/dl67dqYA8HPH0LIP+EchtfnOUOU2ra6uK2vK0CvpR3A6PQABEj1nGl
7v2PKmtO8tq5lpIdYz/Yr1/fCVRf+NzJwMgEhOSpS5RYbdH0zhW1UNk6+DCtPhRJ3ZIt6T4z7dg0
yZw5YWcWfSTTXCOMQ9vrhnXyUomT8VkD5B2GRum9DKYR1ySvdMCGIDmXok9v+lnrwx5to+CHeoUK
AYUzqEK+wyzE3NzixeyvTnJvfYKd+mU43fB/ek2iIx/APaSah2emmLTEeUJUjwrSPoXGz12JyZfW
1UKAjOEYXLgzirO7XRCSQuCVuiUWjjLTxiFwEJCAQdUfYAfyEm0oV2uEb4WdKvzCzTPdL6hHo7ZW
8Y/dhaRRM/TZyCmE7bVgvtiDJlWV6RY5XT1M+/e++BnK+CfaHdXj/MQVUn+GGhIMiXnoxfwH6oRJ
HRAPMwBMvJBFCDMu/2+JMkBPjIP+DcAjp2khQu6vH/DF20zw+Xu20WBIUATE7eEsMCo23JYq3KHS
2pGpxu/sckM8zCcO8/dXZEPFpJqkSkH3HCxY1TpFZiqhzRd3DAlbSfZ0fHHGG2UVMuLYDr71ZDcY
4zHLeoXsMdUXJ+W6lVPjk6X1plN4PP+9vnmevf5s/a4DSfbhAoit2oh86zSWCSvA6qAomNV5vEmZ
4bWeDafTaiagQMxf54r1m90lrCFS5Y0iaU4t8P7IK/YnKfTmZUxnCzUGyW/AFUI/q3lyD3c6ixpP
/j2N8yXyDWb+n3a1z9aNVjK1iCD8l19IHRgcyVVrLGCEeoNY1vY0hc1X4zsYnP5ei1guNPtRC7K+
tFvPSD5Af7D9589M9NnruPxDMftT44ZUMBYOHKX5V5MuXMc7beEtlk/E6KykDPOzSsbTpnFdI+fR
+vferO1+pME9O4Sy9psklWX+YaDzkutQRVuBtjETv7AQ6IYp/mGklQZZHYAAWEgD/vWjAtGONY2k
Dvfv/weEhPSkB5I2VSZ4ZN0Aqu4JOWo1bkWYt72seYB800aaEoWqi9BJuxuSH2/8a9fm8Z6j1qxO
4GuD0aR8jX8IOdClYf6dzIvzg4YPW6jHJ6uqY6bkfvHQSbNgkS6h5lm7Np8nmdwWTsniDeEyT8In
0FiYmd6V445jYL1vCpxP6yCofj+pM1CO6MUfH9lrs0+OPFn/+qc13SqBjPVKDQxLsH9S4vC5Mse1
6VAsiLDukL2vY9KWvdQpyVACLaXeHX4uk2M2zmFY982KY516thru/JTdgtPERLcOWkFL4lLaBZDG
Dz59vdk4ILFzLKJyJko/zwi1PXN/+mZLh3/jRv/d7xAiZhXK5cdwkDO4LIcRYCaB7uhxdMTZV3kD
Wrh8e6a+kho3oacrXqihZrR+ZOeVm/1mkmobNkqk5uhcvBoeXV0dSNVOcj8yFsE7S00jxTx0jckC
IlnghBTKgcoDDG62ufrfi2ihqxQ0HVaa5ZY38kg8zDGsz/FlFul1p5qQgoFza1xOFyeaXTPIqbnR
nIoa+tXxnIKsLoXT/phGVNj02JdczqMnQysP15UgYTKa3Bemn9O0uQR0C1xgOzvzn6i8fj1g7rEn
Z8PVRevhhVPPH4Nc5FIYUULZ7HoWmSRcLvJ9iz07JWBdGxgaDDnJZmvtY0KVkNZP8f1BIjvMLl3C
1eR1M22ixwNOtOfJN7SDOeLXoq1fcBKLMSeb5A0am0ZJjUrB1jX7nqdeBH1d5B+hdADqaJDj3ZjR
t2uaZS3589bL+Tl0bpshhoPUtazoH494vbqWrddGEFZfnMbb9QickiiH3Ml9AybtPBozmLVdII2k
UrchaI6xu9rFhv7aVYmjh6ZJFhoCUUDxdtWub6xrfNsxHnGO4RI/W6lqR27OLeeBe7B/AL5Al9HH
L8NXyTiPUuLcdB0f+gh3fufGAGoo9wFodec78JCpjpxZosO8pMFmfw38XHuozen984gVUY2upuT5
blnXISg3JXFv5gakxjpMGtT379ljLP9ySMbnnCYfnnS3jdAGGBdN+QILkGWiARoRTHYsK3NbSY7Y
gltHYwvxxH71ZMT+Tg9E4e2NpsYsQhlrcHTwHSertpwSb5JOuDmXb7ClBbdKZcCMDUDrQhoj5RGc
AhiuHw2pU1C71/pSOpXudT4THApDlqQNDo4b/QI2qL7oBTbueXJu7lN2FVGj5qYITX9ZNJyFcRlY
ffEmxWNdIMnFlCugy8yQS0/wdgXkjj9ALzAC9xCGtW60YN58DEvwphd7O/O+W1HKeblIVbcW63nR
qSbdyz83rLcjc7UzuHVLNHL6E6U855i8hsuEdLez4Cv+XiC+UjvQo+FeUg+2pw7LjLcIaicFUewJ
QBYLlvzQUmcNilRRCiuA88i76h0f7mOx26GK9szLWE/HOacMuUL2p9bBkqkHb86G+bi5SC1HX1we
06VF3wmdTVZYkj47Eft4TgzBfqc1bMdHOcmd7CC1ZyIvf3E3CozXWv3RJ2qBB1Od/j6l/cT+HsFK
RoKUC+9PAnqsKUpeYER/kRsNBa4nO0bVNgeBTuxnktgjGDfjh4ub1SxBS941TUN+vUsFv7+FoTjX
DtOmZZ0njS3lNBj97y5A8lDj6Ds4aAQuNivZw1gE/Gq5nVxBGD7/5a3c7JzHMoviFhyOUmnykVgF
zf9CeYXjHevKDRJuxdYULtBseNlCRLn8wv91tmIPslJgvEsFwC6UFIWDOCgcOVSmagpaUlS8jYDr
ioGMuHh8Sqen+1EIaZLO7GbF91CH+GerKE6smpCs6SrjYl0Z7jxb5U67o081UuF2FXsBl0ZjNZbO
O912Us1fZZoWX2nD9QDdZise+/Mza3ZQuF75sKK033aqGhwoOosoWi4P9hJWu1PD0YPRed+oZu8m
37vRhPIGAZUBXRkpQo+uqundLBfUUAfm9Calhesc2luG2EQFJWGxHEq11eLgOAJ0hIzdn0GnuNSh
rJVgfOVxO+jozVLtHE3TS9C9vKCaavhjG9N+6sDsflGqKE57oK7veSHfblHVuM8S/1vVFbQczu+D
Pr0+/hKCbd/S/xBAOKCiuo08/08kyUWXQ3W9hMbOHqqU8ivT5KgE88oTMkwIV4ArJFTFYrTl2b22
GtOrYva5dmg+Q6OEDCjd+3yuYwQnR+e66s6VIwbTVigRJ3ZY88XiFm/yHtDQd6qL9YuhxmpPQr40
O9sSOhNHDt6EEwO6aTs7tIOyUE9VhkWhrjzQekns3EUV3KeG1ZocunCftTZzUUO1SQabKw/Ol43P
hsz7oknzf4ZY3532+Zy8WjM/H4Z4gR2vxRvSAaIm8FgQAnvbMjZgT/1pUs6Z4cy1/OTtVgJdF06t
xeE/cRA24z8K69u9ooCaS/SriQezVN3jtk/ls+Ud+OBxTZ48pZG+Hgq+e9wVeMcj6AizBZNvjCid
DAcyajc8dPduFobEEthIIM116a8KY7UQXFvLUerMLms76umyN7+TCjNL+ERQpyPzzwJth10oY+cg
Bk8l/quqqobwmUS59MPUqS9xYb7BMYWLsNwWiLQHDA+nRGkgGMXeU+GOwZPPdLJIquZ8EeXeh07+
PTDhOVuU0+x+cJmKpIWBZPw4/mb/IeSnbvL9KmEK40jogThrGZu1GcphLfRqKoHRA9QHxkGUA6Fk
gYL13E2Mo3FnSXyhRTr8F0i/hkdqUt+E881esPbFZR7EgeIU4fLJJxT4U1JDfl4+gkKAAyexZrwm
UcoDiSQvjFWGQtqjLXaSc13KkWyUptCR1pkH34vS5FZevk4rNw4bsp4cuZHbisFJg8pUD4q4u1LR
c5aWx1irIB+KO+IDCcgqky35H8peKGQfuJ/djsgTiHBQ28/AwZXPR33iG0S/bozG7E5XwzImUkyk
gNhiZtHptd+NsKjhAnSBwe6qi+wufZ3VWk9McCFVoc/qVzfqWQeFN6r5aqHfPwxwjmpLw8dNeW/q
J+qrADrTeYvqdwuyh/6HVYvYajOkvtznB2p2Hgr3AXKRA3xbuD9MK/UfhYUckA5bz8oJoqa6h4B5
w02atF2jap+b7MLrc1ZxsgAFQR5nODXEx+6sFwKbp+qwLYsdaNkTB+2phUmqF2RtH2z9qkPvGPY4
kJX6+4VD3TOsfpLq8i8SgapFNjhyQvgpY31OepkXotOauy75U4ITrMR1dfSf1jc5oBdzxEMUxrLR
m0ea5hMThBO9tCk6UGkxqp4zAAtHVOFA9TpZOgUKIpLlYUR5kyFnZtAxKBMwDq2RHudXjvPoO0cT
u+ftA12jpCOjJfn4m1307FQ8nEDm/s+vw7M1JXxUX+4GAX9SgZUX6ivHeTCYTLAx4FtdrqnOXHYd
DeyVfadQbPaKuMCNPWDN1FftBClvG2imkC1Pk1cuSDJK4FDs1WxhVdA9+psLFJ7xrXRtLhqQAWr/
VDk6kbtdtkxwwuc/Z33bmJ+LMdlDDCQgfSonOVgcWvBl7qul1yPa4uAhebGBnqnkMxbWF3A/lcIX
Vomwc+TKBbIgDLIVk0jGxJqR6pgOLP23oRumN+cGZJYMwy00qBPJaciqhBW2lFQd4s/DVaXcU/aY
sN+/rhVo0W1oWdz16RGT9JMLsMAnrMiJgKmfPQMCekbO2Lp0OatD4KkLIjh6NCDEXoOMhR2ayBQE
WXtD5Ci5M3JNRQ1VcoiyfribnQXpS2zogQagQMZDxQodPMRVgFzwCVEzGpl6IDA5BCr97hOb1BlY
lAUXtIDAURWWKKw7qtGas4sqWo6Ritfc7ftFwQGuiTRrjok3DYUoKNh5VS7e2vwVWIKksTC1UxwY
dOre9N2lQ8Jk4XBIaNQIpSnOLaOW+Maj0BO2gTMKMVJ2FTe+Gfg03BSQag9kTimxnx7SrT7srzH7
MYPCFVWX8+bLQw7VwJ9mHGtUDbs+pJdIa6ujHH3/o9qvkWaNjzw5WA1Uc9MKIq1Wt+7jDkFM1vR6
34i4jHunpEF81qM32Yz+RnoQ+7nOXLZNeC5m9hkaYmwxL1kPvm0j5bEePMZFHohBZFx7mKFl8Pue
2p6BUYVF6nY8ycMFiX6c49fQC9HViqlXjRxO7O3OOXXyJzypwsdugHg6uLM/aZbodkySkNwUuwfZ
f1OBFM3RVHIkxcS2CL+KeY3CGSeSuiLxpjRK2ggoYiYGfQMb3SwXfH0IeEG0Z982ApcKbflGp81W
EQyp1eWyMhTZE+/Hk6s0bZWkrbfQt1HduLmnLVZ9SjYIziTRg8cMGLi3WQf3Y4OupcK+TzQI3P1z
/SzyJPydT0lkbH2IzrkQdawhOlJcv0O3PcQtxpySdsa36iEPXkw/VZKktSGw1uVlErmHpSlKoX2w
fU7BtOWOBs2lwn+YAsgSQLyRB8cTUVmg8RvY1hg93QvVvFts20rzYXEKfCkt2QhD+k5viwb87iHd
vzFXTARAHI4jud8bcMLnRhdLed7nwfoGEnUN7R9W4AaDg2cg+262iGXpcXOYdAYbJl9vDNbJR0vY
oocwElBsjIj3lJCHp2TMzkJyQfoOaVmABYkZWBsRaN2RBBbmiMzzhTPkyFH61700dfe5Z4vPwLq8
I+bsnRm6uX6MJ+ssPJzhxw6xTsrrNrXvmgjxFoBMpyC5AKLWLUumOx//3y60eeoWCekZo3Rfv+9I
FcqZTjuKaDbW53Z15tKHrgt8/qC+9TVM9lXd9BfCDEugeLumpLKGHBEnF1aw5CYC1Ew7K+pM5iO6
JQ3d33c56+fIJBoFIHVQcXWKv6+mqvJCxxBIg2NuHyEwhwO4bfA1aqBfgyZc1Oy3qa05E5itDk10
Fw0X06GyRQV6d7mXYHHi8MW/VNl3Cx1BIPAhX9k48jUnrIfuMr22D+jljxXQ7MOFuVwYAq9zb4HK
7nACubUJSOiMEY/9nhWtxF0l+KDUaomNumTVwF0JL1DsvU9Uwu2efeqe5CiAC2aaWKPmR66rDbyp
azIAwfFOeIDUyQ3AYavvnI4TGrV1vc2hwT+ikXSE6IjSXfxoLIFBP6MAnTqj/nhKesjL7Lb5mDqq
ovwtMDwHInxXQ2zJgWRRxr+XvQPqyHV58SaQHloLOqI95kJbsHyCqW/7mDvIXOWT0/ZbSiiMB4S1
vKZbNXLcTMd7fYRaoeC+DBGOEqeMHXY9p0vO1GfcyPu7EoA8WwI8o88N4K0gHOz7SP39UeKXJQR9
RfrTCNLSZRNao0v3SPjwt1p699pZJuJ8HpRJuNwN5or0B/O7j3sEUG7G+jKilPb1xwawfbD/Vk61
hE1luPch9R9GfbyGMrBKvNYbhRpDYLb3iKeMUX/HYlgwFuvBp2jp9JSIh0ongFl0SRAM+qIBYjVi
6YLNdMOCt7iroG0ZvXDL9pYi5xV24q9/SKKeX3QMvFgu0J2dSEX+xsDTkVXrzq78hms79ayungHT
dK2X8ZWItnefiYljWXDq6uvL6eQkG22/U5lCsceqkED/Ig7ZHCZQFkgeEVV6VBNouWp2sGeL5zCd
GEAykOBLW1HvA2NeGdbGtFBpUvrDy/AAM7A8Ld8igX/1+YMeTeQ0g+ID/fC3ym1t/XreS3/TwgI0
mR+mx/lISm579Tjw1atxDcnYq6BRak5EoDg1OiV9lRxIxD1saPT0b2GJr+OD6RW05y68n2SM/YT/
SQsRKjBxIhRoSy9QCaFaK5QsJiHb4CO6fehYeirJIzCGEP+L59/BAlhOTMsw6wHqrOBswN4iQBMM
B0atUwzRwsjmqzWBx5VtfgnttGIXCj5vl1v8PRA/Gf0FDxVtWCBK445+bm0OkwpZ1TkzhHweRS/C
HxX6Dn3iv5OpNyHOWKj8nXCejcO2Kl0bPdBA15q6BakeqeNV832BURaZxgmgR+UwAdlG41KSl2ep
SaYeeq7LBfJ8hUlQznEWhQgtNrWYCnX3cJzS1JQq7Cqmgs1iVEuxyjFHmjfe4w9O3MKP5EloKsIb
QGnzysNtPi5vUHKGWR3XTAsK7ArGeJGACUHv+D3G/LxS0eY5JVfxHTEZ03koggtxEvPVKYnhu5Mi
7J2zHB1zJ18OaBcZdW+RFNt9TBQ3sGk1DFZVI5vMRyNKEh7fWf5tmDjGqQC/oA7D2r0+DxzxZAJr
er1gUfQraHe3prkfPC8q4zRNFLFPG/5vlCze06lHmAp01WAk1eWc3q0/U15QKWw7H6ZrrWj5JMq0
dKeXVej3LXIB0iCmBU2ZcRwEuRLavgcs0hnrwzB1A4Iwx6OuN2IGbEdBoIXncsjCCicAB56v1LZ8
Bd6f+6PKUQHMf8AgQxaQ7zZ96m/a62bjyKyEp053gHKMdjR4jKfRLAQT+Kw4TM1pcza6Jar+damV
YI52cN938S8wHQMk6md8IAxs5Lip1KQ7E7F+8Xr8CU/3LSGaWwTm0U7s0xUJWmpem6zJs2MnGeHH
4UMQgOV+dUTe3eQhK8YrnC7V38WmGc0t8ecPJihA0EauHXTiSPugwBhPtxoXX0Js4b+H9WfgA9Xx
/J11O4lf41pWo56YCqq9Zx2OFZl3dRQ6vLeqA36qbcfkX0OZSQiAp69xPVeEdXUKSOwxBPv6PDs9
/Lb3pnKSo37PTOh2D7d+RSVCZmtMIYXXzrZvgAauv/+buNKpUdqaP5jcUumVzR2zaXV9xw/UijF3
6Q9DCIOCIesa2e6q4b7Fy/EtSLDWhb8Bugi2r93tZZtiuvm7ejxVICVw65oHQ4qEkcfWyzj7KxK1
YIOUKMgkrqZUe9NDo2GUaLwhYYmjdxfaBV5kSp7tukmGDfFUF27TXU0Y3y4Uza800Ht6amjYtM3j
efr6TwwoozhELjL6YegXXjyItBRJ7Hp8qzQt6EhQCd1Yw/0cZdq9dGhLObfCzql91/UwJ8SH20SF
eCXLmAp+qKTcb5H9YHkUZlOGFH7djjuCMlKfDiNzol7EYeRkQpl5pG1MIZvhIPsHWejMIVjX6Zd+
YV7QrlX0A3uFDcyfepjx4Cd3nN4vAYMczvXZg9s3RPh83lIAY++Ga0LQZfR/KEbGZrphiYnGMCVt
xjrtC0pAh4Nnzbe44SmfHcHhHec4ubuDPb+oV+wqCjeO0BJRbaR3R6YcLnsXD2bXNI2jJjCm56nx
b5d79A84rt/4utiZkyDYza385Ks9q+n2P9hWCErTJpnbtrDGkWgC3VgcjPSoNDXPW+A2Pl5UII6e
dvrDMOxOWcxabtz7G3syBJt782XwIAES/WJgRYW8CXngAd2iwZjtToVtx5IBx0jJrruupIaUmcQo
raP7WqRMm1XQFWiARMwQ/fYm2f++jTomGj050a6kXQzCvgJdENh7NNhz5mrxuVxAMVWJ5jzpcUj1
lCgHCWIaEHNehv5UlH69o9tbhLbWnYuDo/qOpx0Nz0+w3feWN1PwLHkIKg0IL0uQ+owsmUdCve1G
GOvJ940TotH5EuOTy9NIqTZq88/D3NxauMevXVdPRFyhRVL1zkm5gd+zKBxsSSKeF1FNrlJ9TGSh
kYiUWxwMsnLG4BpudJpA4bO+71B/gR4iJT/yz71trkUzI12UDk9p9GtxagWzJ4BF82eBc+YCiXzJ
YhSeFdLbzLgogpWvTx6RF5ThfbRH3vH2n70NockiBbLNA5QPue3c6hhsNvlfQ42hfX3k5QMGgleR
hthVhg7yT3Mz78KLAaeImowN2uVsQXTONjt3aAHz2z3zH74xW7Iil0eDSJ393M290H33ckU/lYFy
S+p8SjlXRc4LjG0hp9T57GkUeBUp75GmGi7GAZmyJ+U9H//SkDnN64bXIiDYy4cEaCAYiF/UXT/k
4ZCFIKCASak4cYxwFbozPbXnh17fBh+zaVwnlrubquZy5KPaofNeDObzdXRoFwWsaScTGjHdXJ4/
82YizfAvaNW86RR9ntkBFDtFG/jWkthFiEOfUxvsoQDNwl9mhEFoWHmA0Dnq7lLxaM/44IZ2w21Z
U21RVOklEjfiZ7cQlQbeGXrVt4PgHBCinaGVpytTgVZugEqaayPI4nmbVbXgi3/DMu3xx7kMMFJS
nzbuWu49tyMfh1Esmc7Ni3YLuLF/YzF8zdy98o55DgKK8WG0J7uHjgXFJuAcqCvuOrtzWn6B2BLg
WUYYYAM+0WwWCNdBLujQ7CHxe4qizqOgFMdkFSZVM8f4GLXMAxKCmzaZfdJbefoiTanloKiu3znR
0UeiaNOzPpVLPQxJI8OOqz4+6i31emGGDn5Uc047I2CCdMUg5ps+YrIVWCzGJFV8jFPpYvDjiJi8
DzNEdXdh8/1MKHSF6sOyIaYZwHpyj4sXHjgEziKfXdMpXLfcfu0POEHmOPl/WmJpLHeJj+CFI1f0
8Nd24keyORVoN/I2520K9gPLyuHn0gdYRluDbR1smyQvCFOe07G4NpIhvBwVLQHy6ay+EPVSWG6C
GLi3QFjLB3Un6b+7kCsJ9akOjPW0BdLduQM1a3sYcrcme/avAEOCBFtvwq5ORg91U4E/RCbUkEHl
aVLZmp5y6LlIG/P3cLVYEQn6EYhHRRiJlPnXQevy3kj/n0d4y36AMR3SCGWWnfCdF3qqEhtV+YWW
i73NIWzI6HY5FC77erA5vUEJFsfaHFZZypucgC9N1QiLlCSsKEnVpotwQDDvzyfqnUtuTQ58Xdhb
9ulVkXymGF7soSNWlWQjJQAfw1y3D+NhWqH039vtMjPtRPQtfJg2D28n0NIz9dx5+q08U49FCzFG
qsLWxr5arLw2RYQsR4sCbU+r8I4qbuqFu9VNLqP9W6HkVGDroEv1RolxxGsYTfhiTSCKsSGYPof/
m8FHK9+zbpt0haRjJTUTj0a206Wb1FdSDZvZnHBgf0HoX2IF/340IZbdutE6U8GqaGNDodOr4Uyx
bAq8SokmU1VCBdhrlVqYWjVpYzsN3qSjSctkvqxCusf1QulCFf4J5hFXCGCMMLjV0XOwPEziXOpJ
u72bS2YzYY+s5i9YG3z9ud1hrrXJQcl2G2rFsyRPeIsnVFyF1I0dSZPwxzwom1Ym0i8KiTzoyPl8
Jcz7NY2ZrLUZFPAOdzPVyWZZndCWGP+ak93RqfN9u1PpNERRKlMsrHdgSwOhSvIe7sKgI2oiPAh6
r7GZ/iiILzP97nAPLkesZN1b806sqsGqHzEP6+jYzJsVhKveSaYgFp7xnBWJKhqs91X6RJWEkvS1
vJ1/m/rTBamsrmdXPsJLYWA2iQ6KZB21+Qa6+DtXhx2/Nb0tcgdOQo3IXjqy8nitPDHc91BYRVIv
thA6Q8DSNC0QZ0q8fC/5XAw9G6zqznfkheW8sz/yT9GiWIIY5OHoPJuGn8EuTVCEM7OdJAu1tjo5
G7aAslW0SXdezL35Pf4lZA3G6w1/UbkvHUovqPYxBPzOmsc9yUJuBqNe6IfJieA/xrc90XsF5wO/
L6UuNUVP3RDKr5jEIcJ0OBRp0cYCkv2RdpojHLFGP3v2Vjq4ww9ZZ8yHViDqsCvsg+vUqC2xnCs2
lMNQUWLjsfcOixClurTawwC+nT6WBnmsjPDz6cNPPDCG/0i9wyIjB5GhVySN1GT6buUM/inEYbQL
5iM+AgKkA2UFFWKhQRH3+AiFd9i+Z2CpRCsKDsw7TXbgZ+vrjOH5tOrp7d9jctkgI2lv5uf9eIHt
C2CurgQslg0Rv/Yp3Z87zwhKbGpHrc7axHxLY9jZHaA2S3W0SgEnBLaWukFQrSTFLgUz6xZK7ciR
8jsYQuwuzWcG3prBdlV1X2B8fiKIrjwdDahBEjLc6SEr9Ch7OgVw8y4B18Sye6MZCu+TF38rDuVS
3tzwGkXkX9GR9uLJRePK8NyFaFRZvSLIP7ppng23u5MLWjFVnpa2pCYH+3T4vagy8NmpKLdIZa0k
gcTjTmhwI5Jkwn/9B7aWrkJJE4enl1pfl8I+bmU0ZNJPC3IJuvWXO6+mT5L6Fx/4IbYrug1E5zKy
KmDEUch4VxF5qx03l5y7RwGMy5FCNkrWckVrR5I4C36EoJcptMIRSDU2R4pcZV5KKW8kkI94T9gX
dRIGmNxcbngxx5xYYjog88yYFbNwwCMsUY39dMaH+jvK+fUA9miQQOiGH4rwbH/tzRS2A3+5QmtH
BcvzrBYmKF9ujwHgrW4inLqhwvj9UyuOsDuyBGSLYwebH0G8C3MFrIGRd/tO1pfUBufff/W/U/HA
NFrtEMmZ3ymJhxXVJmFozwteB8zdu5ShpgbGPVWs1QI7L4+Xt9zKT2+OgduvUYxAef3ZSVpyzgGa
xs9id+WbHnUYNvqXc5qIk/UvH2W5JZTVdpOCwrhXmmgp8sci5l5vnf9IlP36NHEDnl0eU5FEQQB5
GSTxqDQcFagfP4U3ToQ6NVFw99E7NvMtr9cZyowjeFuTFVxXokNlgDnKJVFrXDVsr+ROYx7ra1l3
c/db64cJbjOvRnHIFrwQ9D5EwJuaSJLPy5WucLxenFm9FbYtiz4G8e+rg6JapZt5gPE+rT+4r8s8
v9JcQYWzCSXT/7+jV0AKYz4QXq0XRY9R9xdx+Fv2I8DVdP/enx8whtN2u281IJts8ZMydofGFWRO
RtfP+u/J72arXBHIymHq8+Ix74BqZxyN6AI9/aFDdDk6kkXKje/Tn18Dh2ZRwW3yXL06uIOBASaR
7DXGfJhhGCTiAtsIRb0yG3yANWTjfeiSpt2MSL8G9tIMxRGWceNMqicMXyj08YbbEoWmPTDTGZ2L
roeolS07cXgwK3WQbvbcEmNGA9KnCvQMZYJHtS3flZh8CeEIIL4SJp73RBQ5aiVPLaQV5x0MHkdk
ZexUDnefdznRk53HGvEzH7wdoIli8pp6uyrInJKLxoWWLS+qTzEA9bMNZi3KfREz7wYs52AUFFgT
5Z2/12C4WucQv0K9Ya8NhNcEvhsFT9qFwDwzYH1C0qnUvWtyaxZ1EfUAuLZqLtdAel4a/rs1Dt7K
GBt7XL5QPExezoG/IRo1OjtfElp+LQlTPJwOI5jioR8xEo6A7AWUFbzw7NoGAlsnE3WeBro4xlk7
dyHv2UJA2zLzslbkGZnWWpCLP+opjIpW7K6yo0gdEOe4qkJWV2Oi73viu3spLwFBhCRokFeFbJYd
FWLa8suUHR8Q3bakMwE2Xl1aw4Db+e2Za51FQusnIqiJ23zDeL1GLT+XRyvKaj4hfStfRZfXeDSF
dZhfpXMChzIhteKVJH3wrWuWUlxfQY7xDDIWj338vnHCgLLDR8enZDZ0SdcgTGsL5ll+Sva98l6y
/OVTZ0SJh4lFXBbpSw21JVA7So/Ws0M/xZa7W2Guj4krpFSymKPQdc4iHQwmO69tGmtzZbBSmzZm
f1tANYyd6wSG6ffI1nwOv3L4W2jxsJdlTMtrHg+99gMxasW/GPjpq+zyiKGYzpUf2fXFevFu99N6
h7DcuLSD9YMOW5XLbP74q5eiKABr+2r0iltgdF7KeQ0ZQUJrd+klGpGsTdyWUS6tFeW4mdKRwQQs
gXInH50Ud+r5/rAeHyHRE13PoGCPfaxoSKRgDiztAFeaetd9TYOIkWtpqqgFuEghpiSs1yWBTYJE
egkNpMDsM7yW6TTAidLJMZgaygwevKwMqHnI/Fy9Vd4NsW9XGecixtfLOCyAccKJhf7DStoWPe+7
tfo6Jvm1NdFPWNQMX0vvjoAdtW6sJh9guwm/BOgBamjUvgx5C6wkukDpLi+aV+0xpNiWf609cUow
hOU6fyS890XJvbB4YeEmpqTptK78O7p22o65Mn09m97I4r75ETzukCGEhIamXrh/2R8+uUIBsg6G
J/dH1sZTH7Dgx43OKh/2IrQEf6c6eykKCI8n9Wy0iPnHuuLCo1hCcWPWdb9ZH9CLyb+cd6vGovRO
lilMPJaI605jlMIsvWeQ9UssWNFS1ucP+UhnFk4pulFBt1uSLhgtDZfdtkewcugYiXDGGcGgYi73
fnypyvj0aAg1buOFDk2ntDnThrspbL6m5qrpMbBmjxg0dm7tZIormZ5iNxhC+77FnwG99XJE7IbM
kKD9xCoNwG2MT5PJPoX78fv4TEcYIJSiDDbcNyDC3/oFg5wCKaQYIm/wkoNBNAU3IvP3Dt8jxYK7
/syRKBWHSgFXiRXPi2d2nABiq8WFYHGSIYLq9IAgDfNV6HhCLKfoQ+ZtvAFrp6rzjdFTN11tresx
Ta9TplZxPS0LE4leL8HhdIpI+A8nVByRVB1MnlPZZLJn3MmxsT3PLgSPuMoRDZXkEQQQpbBwmMYD
w83ME8Q3Htgh5SBezt1O8+0+TyDRWPPFc0+iMniTvwb3KDrlfkZ4lxC1bLEt0xSO2MnF2pt6GP4s
AaKliTtGmK16Ib3B2K8JwAoLBxNPrsvfkaZobE85GfAzo3kGcZObijjhU2JjD7+eYCtSfVJh5DWf
jfA/YBWzGoabTHt8UmSnMuyltwg+ejSPXv1nxHhRidfC00VnKb6E95TGM3iaYga9jxf+BUiEdcvZ
4Qxe9owrui4xl1EzETZr9togDv8UqOkPjWthWBh/Hy35Fl69zgQJWhjMZIcZG6yxeS4PV4CR7EvZ
Ss9yWluFZbiSNbyCmMf+N9QM18GyOdY/Sozen47ZnihVAv3gRImtC2xyWy77o131azGC6TzTwxQW
xJ7h5epe67bskdy4g/7eRnLITe3lNzpSL5KEmLP8Kw2xa/x+olyBWSWkUZZSU/DVkQqhMsLGjjsx
nzPx2uW9XxDpfCuLiGh55R0gF/B68kegBzZO9oHQeQ3CKmGxkwGQm45E74NzcJHvWp2GeWgr6atD
0nxGYJAJzUaHka+Pwwze14esI53MGhg1tdeLbTKefZb0avxKNbpmlxabAy5hXfX9m+QyPMOzNZGc
4aVDBUSJdoJ0+j4EnvW6b0ekkd9Hd7kr30vzvQI/iAK7adnQu5aA/XArLcNGAZK0oieYrXsBT405
akJ5HboIq1zPXQfSxDoIKoiaBdpLLFjkmLOByyONVOAJdDDfuJr2/f0PgmQ4lZjfdAEUDQ0YncjK
r6m6nSvHfo2bBIXECGjHuyCh7EAj1cWseRfb9Zszm04N6Y0UWecol4ac5IEvjfB4pcj6uCYQ99Al
pM+z/8EJtjsKhk7/OnZl2oLxbaE/popI+eOhJQZuMdt814eiL9FxwPqP09PpUpdJRClTldiNIisd
wOMxyLOq94krNli2XPvNozWi0WJrTYxoB1ZRwimeYgWlIFvkpQ8TC/5+KLQpYW4KQ28eM2c1cox5
/IyWQaMg+Tu9xevX0EHCwCu9zgP/8GuXYoDLCiaEJK4QpT+7mvIy+pC1vEqlVAGGPjLuFeSf51nQ
LsVrZ6pFXVIuvnUqfC2Qhj+juUfrIGv65Wo90C1OQlVf87WfPz7r1ojPGV4fVwhX8FCyX22oYoeC
lNUhWJBm+iBN/mQdxBj8kX3AsauvSYb0DfhED9HK1CJVjDkbAgCsq71I5Io3czFMsbmJ2gZq0/IO
fa+P0Xn1bj4W+w+2OyN3CbqQrouYTEXiw7yK02U/lh5HsbN7gUOeqqnJ3PaMDOZpMjTyTTH/+hWA
FA/z36xbGGRSFagTQ5sCkh/tEyVdKme9UkZxlWE6SR6Rn0fHKvGEyhIHddNWfAi8y0AFpRRwK+Vx
SVtisRkjbwVcNaM1hGi/n1sFkRHnMl7qGTGU9wprc/ehEcqf/c5Pt9HYxtLnhgekBOEE3UXHjWDr
/Irf+TmOyJ1PbH148rZIxSMc/YeKYETYgXq4SFw9XB1VwyZ2Lhj1HJfHjldhMOOvG7N7sg0kSJqQ
v0Ul7/9NKkhLpnwQm1U6BsLCAm+joRTwd/f7rvJK85eKOiPqsgnlZVyyn74Vcevw/d4Ld1DNGMDF
+fSN/QIM++ALuTKmnmuCFYkitOVWd8iG0jSqp0KTdxUDJm9XfnWFeSs5v4w+JP+cGfp4u7L8kJ99
V9ezbKvLTdyudjG0WBuMKxn69XVx1rQ6QS6ikY8qX9SgA0mfqhQuR0i+lB1Ksdm1F1MlTxEkm30f
W6+kNTTxS6o/H1G3/YmVHAAHRrFCWcpvNa9bFqymveJAbW8l3GvetUp6w1Fm2Rjpaxy5/nzMn4pe
WlYB4NbEeL4M43vqc+hxxw4M/ZZ//ARWSGooSyjbC4dGl92VQ9ERiA6jj960uQN2ZOZBCCAaF50D
CCgSPc5oxy6sgPxMb4bvDCTXg0uOQcBq8RysABor8HeWV9LipOt5cdLO6OssGJotH1OScPnGoXto
aowBubHtEFO0zE7U98nP+W3LsZ5EjtEqCSQftIad5ADwpARTBnNfQjI2jtnFAYS72EyBEiM0hUny
dsD980bjhl2OXkA2bbQnr40/ecjvZHaX0P7pdp9rl3QPpL2ppo7YxgERDFvBozXRMND6Y4JLh52X
QfKKzQ8ICdGnnjjZmWqZ9T35mTZ+j8+IJWmrhpaQ6fcteU6TBkGgIl2VWVKOOCrm5P4DkTmycjl4
+dOychpL1q/3mR69Rf3hEfyFHFCdAD90pETJMVW1w58/a3lsin+z1aXy853yMVqWGTEDiyes/cAt
uEZlVxavZn+gaLqHngNy5m1LW3Itwe5Qbi2t8X334pnl8yDYxCRdrNUh5TlsD9SQyZzO9nfLfGdE
/4bC/JnJ6dRoR13w1wMxpMH/txUGC7OA6YCO3yZFkXCT958OiCh+Cp1a0AZudPf/P0rzdZ5G0sJj
saeXl27jnIR30cLkn3fMoF1eMkgx1kr57xrzkG3ONTjBIinlzyyZVRmsidxTkEreMKPz8AMIrBIA
MnYNUnsLG4Q7kXkgiiNMxAoGRQot6ncURhbuyVeijRYxn2yBtsx2qreATuANm/puvfF7q7VUzfXk
rVdYxW549Gj2fVFtq6QyYtTy8lFVl5AMQ9yl1asy5hztjraOVRh1dwp5brRY9iXgxWAgx5WNKMof
t+CMI7lsOYCW+qXh6y4h+loMEkdOTqLOYY4YDKfsyJVsuvjEo2r3xFJgMI0WZ48LfRGY4MnDFUOy
BSLZXbpcc+0X5ACRZJxE4ATQFdvdWXaZHYBjPf6bjmL35O0gLp/HIqQuPI+ufSY1aV5h66M6OIy2
pwcBBK4OetURpob8rChdjhaQ9wBMZncbfC7R7rVQgqzuBLnTaScB+JefYmyvbz0Yw+mffR+jllzn
7uWS/dxHwT6EjMW5vdCXzexRCAAWMhh8tdvHffuNZVeG1rlsV2uLyzZXAvkP3ePAb/j9k3mKrxDv
oBnVgyFwnjJ6e9nA2CyBi7uZQaZTzEUE1TSxJELFd6nM/rjHZx8VzlnRziJgaHzgxB+Asb4iWFrM
O0m3C0NocYzePVep+3575U/0/8kCCYIMT1CFWuaH9BpsXVoLQ3h7uE3Nbu5ftVMl9nrDTph8mcxi
H9loCkTx5YmhMukPtQx+2RFUwKUIqRJOJgU7iMxsZZODyfg2My6A1/ML7rhSc71h1oHoFS6wEsC6
p73+taprxAfOF9PYP0uzBnZ2c17eVRdcWrPmVBsOuEWwVbZH4lLdZmPTYyOTj6KdyACokN/n5/RS
aeAEqzfK2TmXo/gEo16Aj5tugehQnMgglyERdLy9Wr9HTVtAMiRQ7m/rZUbj0I4Yc4yfGICf8meD
/fvOq6FT1IlJlCOW8s1TUaOQJuvHI/ifvW1llQrSFxyN/ridjbjdu+hIZm16BSTaFgkfOMKsFfoU
Da0fIdEE/bG3cs+QLe4TWpdZOceeGXnaEjwYaKmUERxkBX/XS7njR4Hc+1Vn3YLN+SSOU0zoVvh7
DznTJbv6VGYC0neAXU/ls1gst+9533wijhkC8sqefGRywgZs3Cipiowg92CUacpi98yaDU7AERJr
K6izP9mg/G6/DjayHU0yUmTGNkOHS1dR/J9zAcKP8/HDOjTzBgM8AN6aOu7qB46PoopwBExwxaLu
JYu7W360XKYUYh79cPGKrKFzlAdGATk8go+zG9aoW3Y3fFG4QniRsNs6XocKwuOzGli5tKlGPg/z
7KN+cuRRRlCCsodB5NtSYicwWOs2Z0MnCVzRyaCor+eOYY1+YBF/luWVRNV6CSlrCLk4NGRqekUp
d0cbSbNcQGaqK8GIvkjV2oJ8Qm015PVxdir5iUA888HIglg52VXd2DSNw94dQ91foyOKVAefCD4G
91L5Rm4GGRtNdNiABjWfSfCxg+QwjSfzNQmWHWvDcXUw0f7UgFY+/7iv/scoDqQg4tWfOQS4AdON
qFNQSQcpKlAgsvVgjz0eP4CecSicYG8RNIvezxZWvq57Sev01EJWcctz4xQZ25+nb0Bokj4Rj6aP
4xqqj6NzQDaZV5UFZdfAdEAnCcOOmYDh0H55ui12izIOc42ykEt8QqTSghQG
`protect end_protected
