`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
obXXhxRlTaHjCpJV4uPTkRwgR3GpcvDfot0y8VTPyFxY1NMmmd9nxF2yYzxY4op4aE47wJsPh3ch
Ifk4Z8Oulg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hmzRe/Qr+6nIcxuhkGdjIkYxpmHpO2VQJwayWf2lxaeB8TRqxhanf79tJphTIT7qZJNlaejd5WBb
CQ1aMumla5wg4w9VFCJ3RfIX218tcMJOolbR14I3sidO+tsZwyzxKpPgnD/kd4T877IMOTrRvnIx
6PdsYAvnCf3xQFi7I2w=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
x0fTehxzghnOkOVVaF5ZPRso1LEjaAT4Ij9Za1bH3Oj/tMEqkw6sMVwuBHCx+9OVt2006A4ekCrO
o6bGNZkP9ZTi3rPDQxJqDp8sg5+LnJfN79zDXHa15RdmKwVkjgf3nwhk4ny+EFYVb0Y54aV8MR9O
zAXbiBIex84Cf/eo0y4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ic1yv1cEiezEPDPgDJrMxh9C2VwWquV93tLinJarxYj+AmqpzKzI5K1H2OQZe7dbFN/MWnbwXkU3
VZ4HTFO2LNY6CAQ7agHefFUAhNGwX0QRTr7VGuTBYmzhsAHdeMqszybd5GeRvJKr6TK24gNATQrN
nT2+HjrdVmQVjknT/su1Hfhm/cYUP3DwaHb/YUh3OhjGRMtE/ZGv2ChKMu2k7R9vmk5m/gNYJ2nE
08anLKgzUjVJXgO49+Y0G/wzgXuirkniHC7vyzJoNICrYz2RxJ622p1143uKw66xJyQQhrd2qIBT
Jl/KhVnIuyuaJXAkrqwFPiigy+IHyR/snmCbug==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LFux42eTG7g9Qxp237PDkKB2zzr08ZwHBtwQiK5Ci6HPYEcDQC5ARtEmy5K+FX4t3iGvCUCf7B7w
WkQZxeuQq5Pu6G1UdqUYoZkYnIGvv/FBS58O80A7wz1hDYmIuCFtceYj9Pc2fMtYY1GsiMPo8DHK
SwPJ/nBgoPhAul+T5S2sYyEyPKDBAHo2NS+ueZipFxaUmHpYSWv2JHPg5npmpprgScJtWI7t52dF
UBV3yLc4chOAUHmW60pHDB60diNc3yRD3AWRAYuPmEcz797OhGqtq/0Gf/sQq2aaRuUjcjmv7RjV
F0UQ0AGzw4qc2pK/6BN6qq92U2093f2LWTUUxA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mLsPIi/Ovuty+EZo5FSaXGTuskBHoX/S7M5BlV63QV6xgpHFSsvDZ9Xz7MoE307jvEG7GvmYbswJ
7MgGzFiYjlGDXcPhjku9wDs+Lmtnt1wDk3JEvFz7Qw/y4xrtBAKwKEzSCJWoN1fsuG/a1bHGMBW9
QIANQXT/XtWTLwK/eGYczVjN8LvuNEgutpT0ch7ABudM0jLaNAh74dH36yQSfhAmYUPLYgwDG1YG
+aO/K3xh2vVQGtq+ZMzL4D6TG82lwyl33sG5zqpY5BEVhRG0s6EN4POou3ixu/Cj3dzQaQQh4MGA
wnkI7caqlqGiTD7K0fMqU6D6LxVakb07jRj56Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4784)
`protect data_block
ZSNt4Iv9z7W52E4HVDUrJbeeR7Q0PW2t0Pfo6v3+LQGHCwgYhwzTe4JnjSXGYdxieaZqe91npCPD
PCGvcZkjQRlHKK7g4ch4C4+GTed+K8R1ZHdKSHk+OhXeOBFkDQjUdWgTDZa68CBpHYZY76DH7KgU
8qYtHccaYNEh7/UIFgwfGQ0aFOH5eLdecljwOvUE+F6F39iAw8E3php/NptUT4Tb9vOhKy8qcOsK
vCbBiKEwXQnRJopmciPBQcTAMJvbnoPtXVG/eueYIppoYUl/oP6THRqxyEhOkT0sgtzSc1ZQumUo
Yzz4zSCOMinVrIPRXtuD7nJ6PKiKfaHlGrr5+slvt5sk7aU+1qSnqSZEXKjkUriMkmRi1r4Z+knX
hCTnGND5A+kEmuYfDZMGqteG47dS1+vR2hxMv666pDernJCwf5HsLAwcRcMdBDZXCb8Kxg6teVFd
qMdm7K3z9H2sjtp22HbRvwlauDQcYd1LLR1RwUMIALPentT0khk4D2PlqVjAtEUgoGeNEb5RhWS3
nP1OCkpxulsEDktZycTr1NMuDDiibFjzjFdR5r/cRWRMtMHOh+QuQZlN6a+pycpceVjbnQ0pKd85
mf/wLzlpVKP8VJ6itKiPg5c6oXzdyUm01uCeUbd64QcL7kodY7T2Q2qct44MynQTDHMBhdCMOreH
EvtvmGAPNh3UdvPt+csvgfWv6GHoXJnTASazUNGXUu/E5QnvAdZze4hxdrdugJq5ZVc87bfYplNA
W53S70bu+CItwc2Y2nnZ8uPBUpky4iuwqN8BPjM3wn3lcyRskVoYPb7mBGLsgphtPViRb0hFTzIF
38cEw7+cU1uHUdzsKe3fSPtsK13AGLKiUHg1PPEvnlDgBoFm7mYYBMW2imejgRNkDmvL9+jD895W
m0FlQ9V+rJrx+bdysXPO8qOOcG9jfCuWa2wyZr/CjvLcn5h3b0b1K9zCj4aj6fLsf3VQcVcgYhLk
/FTghPRp5qbFPJi3WDS/31ESiE4tdqZgVizpn5gYnpF5L/ZDlsvsj6v3Jbx3CSfP+3vk/r7uHakm
2cxZNo4H3eKAjce7EmGDa/yL8dv/1JOmiQr9Zj/5zvMq5tDpEcrKnS8iap09k8GtbkaqkKbarhA3
2DI/5ycas0lqD8+af0nmarNxbBzDZK03E2AYC13HFPqIwcrCTmGsGYC/EhO+JeeRlntOovkJD6tO
Hp07A+qDZju0pFDg9Py2gYP+hMo4HQqbRsPzruDvra5SIMkba4J8fdEEpnf24ZHdCmewFSeBeHx0
x9rPxx4gQDRUKA5u+b8Av4dlaM8H3MJ55HfunJaeFf43wUf332Jq7M0CWhDDonRmQsYMuFesuF0O
u2DYdNKq6FSYU4svIrdPqrlFQur5p2k8RrUrXw8R/1EMYo6BGhOmA0pLN3Gq8VywxAcIMZsTFZQp
hGtYdtdEZwTCuKpMt4JHSO8r1LX8t7r3JUwGOWXbl8wM5OaynsfQ8gj7lGVpkeQRpo4WvLLL4Pkf
97fTAwt6K46juscyoqGkx3Is9bRfJ/kMTguHvpM8yue8Hi73e5F52L4pb4Q9KM7Ecu0BAip5XtI6
M92oP85L+WV+/AiFiInKLGIhvx53m6+IhumuCfrh1cZdI6yD6oJnPmisZpH+CH+H7qmZGz9VPYX2
9yyXXD6haz48ntLBzOGzsWS3IzADnNALuZKS+XZ5aoA3uy5SQlEgUDaCSWnV42qygdNQKxkqvPUA
ud2cVbDs6C1kp0m37JVMOShiSx4YGoNZYjEkJXgCRasqFMJmD6/lkWJNqhkRKJBlYKO2jfyN2fLe
UXxUfp6EmNU5iO8JXfbPQ/LMNTDQq5lg3BYUEsTmebKdKd2g6ZYLa1tdb1wcHtUPCaHhZVdnWXk0
cvkM3KUf/xLcTsbSNRbIL2dPOHKOD2nJ6i4bsiQc2kYFMNINc4mJ+4asFGGeh9eMtFQ3i5OW7jdk
ps7tfOK4MJIjoHmorn/rPK/HmFOcEwJaaoL2WfD2zDw33zs6NXzewkLN/9LVmN4W/Z/NXzfKGMrw
bFJimaTU32sHsYkyI+JnArLTDtxtmqpNp2HUNoDdTTgUrD7ysZ4bH7hDFbGw7kyBI/ccnxHJWNE/
gZ/pIwCfXURv8rVPT2p5RwMcxE3q6G6rCl5cKbvk6UpiLlPd8QcZz4Ksuz6EbuZhzlLmxbSCowu4
mGzFliTYuvjbz6GqKHImzWKymh0Z0iWvM7jUkvEGuUSaz1XESacXorGXAU1zmhfGCdHXYblQODvA
X3mjQEpfLQCtOxWDjr4qG/8zwSSXPy709mBJphXa1tuF2Bz9EmGjYbqeJ2jOkXk0GVfamJ3P3zcu
ErbfBi+wBYZLBfAMliprD4WWkQ0zVkZ19s11gNbqZytuoYxnmgGAdKSN2dAN2SGRqT6h5CynjeU7
qE1TRSyH53yHY7IuLytyWSsT+Y/o1PVGpYbneGUSb9iOUR3ZarX4Y256zSz8ysP+uppBW+u7md11
QOSI1QxuXa74VBGc6H4/IpwBLgA8CSZVlgDAqd5Qgb3yt0wcSM++i89xyJte377GJfeGoXZIKe3V
88Z2/RaMc31JkiNYiPCtJx+UspWBzJbPgW93foSeT9vDbMvuniV2mV0ZSSguHSfp+ztuuNhS2QCU
P9ie3SJgwpb2xaXq2cX5I7yzygUGfZjBnMqUGnKkhzZmNCSx+lmcOpJnQeKN8lxIjAK/mEfALu6L
8zxlaoQAn1yYnFJV9BNaeh01c2T7ew8rEK0Du9JFQcOtx39IOTxpKpb1S74E00A9M3H9a9izhtTF
sDxdYJi6j2TE6GY9DZci8yOLD//yCn3V4b44jRoTEERfSk+Ej+gBoDin4KJpxj/3qRFfaC9mVtY2
cNOze20+yLld4s63QG8Ki3XvGca/GuulGycw1ApBVMbb7R7Fo4sPbwYnVex0dU24k1d/GAP9Q6S8
OI9rBQC3O3tm9plj1Y8WS3qoPbKZGVB+k4Jh8vLllY78TwbM0vHFkK2I37ruT1yGslIBBUVo+N+A
ZOhtYTpr+fvStfNWwNhIAHzyBH/RuUour7fdLS9TQ3C+jDfLk675H0FeSgRxXdEoWX9dxoU15IuJ
DiOmq5BgMLPz6KH45G/yQZLYWLKlttFqjXw85JjeDCmynidQktJgvVdiaZp1LX6vnGA/nQ9VWWgm
gn+y6VAwWhMh4w4Flvi8qUcggIvvRxKiISTM4bPN6Vrt7nwO8eHVLTI/5U6uEJpWzTnmmsq6HtOT
RXb2Bfj12bB2aURtQaIIw6wFclwvpkEIGAJeK5Pi+pekmN3a2LTi9Y9AGi7Frf6q6qEEHFs09cid
OWYWO7RcWIbWIM3aZgA1ziW/vodSjqx9w4e7E/tCgbolXu8I21lBVqpjyrrumcZqthlAOJknfmV1
iETVMf2Nw9XauKxMxw7TuHq+UmMvm4nuDrj8lfPR24/ZB4Mjyb2/cdtlqeozybBmSr2YhDyGiK7P
qPpKM5NiJa5kLlwmWGCp9kgREhbl4JBvRCDlKgwjjvaY8OQOOkf+zEM+f74lZ+r3ILkQJJQWF7AB
WJFgZ08lwcmjO/rOzM5QblElqrV8Ugg50F/uGUsasQwon8ZwBD3EUjy0867uzSWKgQ1xJo9KxoLN
TCZwAQaR0IGtQ5ImvwwOJqedWDm6c3DlHVcijeYMMGDexLu8zwZzemeSA97GBjLOfQhh86u07vtg
z8N5cE/j/HQrt7aXT2EWC5K4v4Ei1dvGTeVCxj03PAjm5KmZs7APh3giN740jIOsVxGiVvNWw9tV
zpwa1TBt9nqnD0Nwwlj0X2fp7iLg3kAvuMoBczpEAfcVWe85SDf1NjcfQuD6Alf1Ewo5LhEFZFn5
LxAg6iJT3DTT/S8YdV2Shqxmkgwylmokx8j0FwDyEERwF9jPoH2dLM9hWwu7An7vENaJqjbVrxgE
ua1iPVkf/d0cjvss2+nlNXiO7gb81i80YUMd//zRCdkbT8ddkjaePlQS4t6rMxiitR5DU9oKx7J3
kPOuyIKy1NPQYLXrwnZFQ2lI8Af3IgaXNADjwFb8s/UFJD9AVRw2Gdk9tpsbhZivZRomaDsV4L48
KKh2b3aPrTKNausgYSqLFztQLIP1YywQuEyQNkRjGw/P2JopmZ97hskPuJqtg91Wv7AlVj4xOLu3
Qy2uYBBfNmMsapdk9h+7dz5Rw88EC1x7bcm28rtVlOAc2ry/Qq1WR6cfsdnGjYRNj4m158mz6Jk/
Wp2EuQ7J5uVLvgZdSfOFomBzfFc4Oz/N0zcZmBO9uru6YAn5VRXyMgqEhxTDFpVGniTE9eOXDeCn
RnKzvcf09msWOSeV2i3GOChaCdBlmujyrm5gbFGjzF6Skyuymggffl7YzB+i/lPcVcyuJgLD0WzX
HcnFvOjBC0AKA5scI0XeHGM99CSqPpO/hvwk5FzYN9guSeKmqZdZg8dR+Se/BeQJPj6FlBbaKOvD
wUxVQpp6bwgwKjk6u5rSTnE+zt1tMR4xiCxmX+2Yh0jN9MlQZOd53WFTipFa4meUDgR6Kx75sU9T
PLlYti2aGdxuKrLXvUMOPE30kw6mNoI/ULeZatXwJ6giGrQFmSJ9Hkq8R5v+knddu1dnkiQCneNJ
unMuibIn63RmftcUgZxoSOTMYb9g+sCCvjc/qLtnqlXDYl/8fcQv1pmDlQ+RDrvkaLwfj2JEuJVZ
Qpwf75hA47x3QNxM3j+Czwl8wzg+ZQy+2G8iNTfWF9eqzVFSENGi3ZQ4TffBjZEtwqE/No9cMutY
CiOyHBELMTrzpwAcV7H5XVi+/TBgZm/2qyi9Vc0/ba/Eiq4c4w2Tl9b8TfDvbJvLTQoXu8NqacdF
opT7agzWYfH6cNjnkhbO4EeHRsKHsl0TVN/yq7ckxpfsZX6QAIOJ0pi+wCk0sRrRucPtakZJHKid
oAWyqmc8spww5jJqWuOfDEpKamV5bGPX6Jp0Ff0JwzN+CBl3ORxMV4G4eiOouYmAln/iDsMUURAj
AuXYKT+9ftGLkBxeER5Roop9s4w9Uqjnl0iaOabLSdsfk0uAyaZtfbu/50RqDYyXlKZzNaTKpBJm
Ya7vaztCNgfHX/p7O5hUl0DrDmHoVN50fGmCZ2XyKRyEG/anTmE1+ueqqvOH+1iFFbMreGxDpmkU
EnTm5swWaPyX8qgnhqA+vG7/xxqWqrVqt/k4f1M+ae5mZ5wHZow/VGhyDt3MQjqjGh9qSwRMujIN
1PGFOmkeKCO8B0glqLU1gSV+fdQkbWRLTLUe738AssyW+qEcObL8PBMde2CP2AWkZ/zLV8I+ivWW
dc2FOIrZ+yC9fb27mbsy38LO81/73FUZ56c9uINd93BWl+nuAEAFoEvemAUGNNXISS8SRJL3dSRk
uUOq1xcIpMBuFI+pn5svhj5j7tNM1I+hZ+grSHfFRdSoV2u0apN8FW2jbTHlFnfHIhEdH5ugXDW9
IvKuRlwMmFHH9gE26pxbgJckl9ouDusYgHM1sAE/9JhjRKCl8VuHvbCPdNUGVd3OXiYXiPQ5m3mS
0u7qbNUvE95UHwC7ZLWWEXFx8PUTgUwC7CmNL++SbNWTW8XIO3gFFz5X11IPHmDk881pwbXHW8o8
GPKH4hlVH4sEYX4WgcIpxmjw8M4Iy13KQ3UPHDHbYCPth1DqCCCEO5y6DFb5kdD4HFkfkWfby+5Q
Na+eY8szudw2hO0ii0Te1UEIT6YfQ6vjWnkuYz5dJ97UJDvEaDoqZpdL46Y8LCQ2f4txdNkODqK9
GIH2GStWynYBvwNytQ77vSrrh+jlMmFwukNRLQqpb6g12DPysaPXZc3b7LAk2YTsb4oW+zthTGDs
yvntpwvlw9Ed6JIsRMGthVPeChA677u7VlJ6VaJGFshJnAJgE+P4tvSm2ZmqbAIEB1pl0wolwJ1Z
fgnPIy4mViCc8f1ZLMTNLuRvgU1DBnUOfYysF0xxEfHhGgl27QUHX777ZOc01iBTxqWsxDbA3h/6
+yvs3cTNFUz4x41mZ3UG85+qOvZPvDh/Nb7XxNKQA/HyPRsvn23a+L9migDTxzwaLNGutmH8uqSz
GNp2OGYi2TDh8O5VLtjCkZW7Y121GkXX0gIzDuet5C0fLBc8iUzKNV357G1+GCpZrwjEsIkVVsg9
2QQRcUEN63sjX8MFnuhoSxvYG5puHMDkFblIHlJNKkNp9RKVI2iCuIocRBv0uE9yPGDCm53PPhkj
JRTi1m4KqRsumIQ/QusktK1jutFcH4s92bCHaP6eN91L6BG052u3M63hMVsCRrxD17NTNVuyxxo4
HdC/Ay+tcqt7/SluE8d29MUd4mta7cOsCYK2ng8ODWH0UrlHT3ufN9LrgGxICOisyDhj1C8=
`protect end_protected
