`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
obXXhxRlTaHjCpJV4uPTkRwgR3GpcvDfot0y8VTPyFxY1NMmmd9nxF2yYzxY4op4aE47wJsPh3ch
Ifk4Z8Oulg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hmzRe/Qr+6nIcxuhkGdjIkYxpmHpO2VQJwayWf2lxaeB8TRqxhanf79tJphTIT7qZJNlaejd5WBb
CQ1aMumla5wg4w9VFCJ3RfIX218tcMJOolbR14I3sidO+tsZwyzxKpPgnD/kd4T877IMOTrRvnIx
6PdsYAvnCf3xQFi7I2w=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
x0fTehxzghnOkOVVaF5ZPRso1LEjaAT4Ij9Za1bH3Oj/tMEqkw6sMVwuBHCx+9OVt2006A4ekCrO
o6bGNZkP9ZTi3rPDQxJqDp8sg5+LnJfN79zDXHa15RdmKwVkjgf3nwhk4ny+EFYVb0Y54aV8MR9O
zAXbiBIex84Cf/eo0y4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ic1yv1cEiezEPDPgDJrMxh9C2VwWquV93tLinJarxYj+AmqpzKzI5K1H2OQZe7dbFN/MWnbwXkU3
VZ4HTFO2LNY6CAQ7agHefFUAhNGwX0QRTr7VGuTBYmzhsAHdeMqszybd5GeRvJKr6TK24gNATQrN
nT2+HjrdVmQVjknT/su1Hfhm/cYUP3DwaHb/YUh3OhjGRMtE/ZGv2ChKMu2k7R9vmk5m/gNYJ2nE
08anLKgzUjVJXgO49+Y0G/wzgXuirkniHC7vyzJoNICrYz2RxJ622p1143uKw66xJyQQhrd2qIBT
Jl/KhVnIuyuaJXAkrqwFPiigy+IHyR/snmCbug==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LFux42eTG7g9Qxp237PDkKB2zzr08ZwHBtwQiK5Ci6HPYEcDQC5ARtEmy5K+FX4t3iGvCUCf7B7w
WkQZxeuQq5Pu6G1UdqUYoZkYnIGvv/FBS58O80A7wz1hDYmIuCFtceYj9Pc2fMtYY1GsiMPo8DHK
SwPJ/nBgoPhAul+T5S2sYyEyPKDBAHo2NS+ueZipFxaUmHpYSWv2JHPg5npmpprgScJtWI7t52dF
UBV3yLc4chOAUHmW60pHDB60diNc3yRD3AWRAYuPmEcz797OhGqtq/0Gf/sQq2aaRuUjcjmv7RjV
F0UQ0AGzw4qc2pK/6BN6qq92U2093f2LWTUUxA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mLsPIi/Ovuty+EZo5FSaXGTuskBHoX/S7M5BlV63QV6xgpHFSsvDZ9Xz7MoE307jvEG7GvmYbswJ
7MgGzFiYjlGDXcPhjku9wDs+Lmtnt1wDk3JEvFz7Qw/y4xrtBAKwKEzSCJWoN1fsuG/a1bHGMBW9
QIANQXT/XtWTLwK/eGYczVjN8LvuNEgutpT0ch7ABudM0jLaNAh74dH36yQSfhAmYUPLYgwDG1YG
+aO/K3xh2vVQGtq+ZMzL4D6TG82lwyl33sG5zqpY5BEVhRG0s6EN4POou3ixu/Cj3dzQaQQh4MGA
wnkI7caqlqGiTD7K0fMqU6D6LxVakb07jRj56Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69472)
`protect data_block
ZSNt4Iv9z7W52E4HVDUrJeMgb+XldKDqCetylmR3xDloDszn1RI4cli6QJboyTTugHpb35VwVP8w
RYH0rPbdXvR5vxC4rNO5zZPVkhSMLR36lXUKymwLB/c5AfSmRUe+7c4MSOF2YA8rP3Xp4bJWdpUy
Y8ZsjGHEm26eq+jL4Mj1m3odQxKbjxAt6UsiGwM+BdcW8rPVh2W5Pht/178zi0/V26wdF7NcFcN4
MWR4ahjRRFEPt8GrppqTPLdK0B6VuIZA6djURspniDLn9NK36m7PtNlBNGnlMOe+R/qs6OwJi81V
2Bk1mH5nCyrJjr0Ia94pJIkgtL+Qc9Ch2PUwYGtOP3mJMQ41AIGMiwMz2FfK11stDvGssgdvUdlf
bFuRKf0Hu+rsTESXC5hqBCTo2Xh1uUq1JJURTZbvC1B8xvou5sClL3gqLuKE1938HQ1F6+i/8csS
rzr0CPYIWKr+ojSTtmmtf7sjUVVdacVHkvxtBV3tWU57+B/4ejSSO/p7BCSV5HccE1R0cBKhyvy/
4zna4YQyR31Rw4viAxBzyhd2lQt3DmYlpOZl+a0ZeoZJfT3yZEqt9m+7tVNJvEUV77GIgpX9PHIv
4Im/VixH/P8Y/FrJDPR8xZ4SQouOSX+YX44GuPMpuz7Ll2cgyFSdY6WqqKJy2ra7UB5CIKzeqBI+
ZR0anenXY0nbw8v2RxShKwsIsFIQKC41z6mQnIPjs0a0cJ2B3ILK+JzablJIZKbi29p16uhzqEYj
3sIQ2Fz+L2/e5px8n2LMfrdOtky3q4EgYUivnOCG6MJ+idK9ko//YidDumPmrMUZtPVclY+Iiov9
5um5Qjz3TnR1Vae8pj465wiQtxdjfvj9ZlUm0GtOVFApNdF8oZKABjK1FmGsSNJh08PGdU8j04Cc
ruMvej0DKg2Lj2cFUA10fq/VEUJ8eAkvCbZdqw8PXTZjYGjYATbHfZggIjKXOJyXPePr3L7QIpYC
4ZSz0VFsw8HmZ8E3nCL8obzC+JfOlc7Pqa5Az/hsfWvUYWMfJIGcpu8PCvY1mWJmU3djk4vF403z
bwVjSfg2Ul3YQZ7IcUKeDCHxVqv8+XGOVbPadtvUnkA8YECw8KXfrN47VwIbGoYDlaSsHpSqr9q1
va5vqeghDrmLjDKd1EJ5M7KuuceQwj0JYg7JhN5DJCuWQaNHNSqkKlax9phQobgu8SBPigAWTzh4
TzXEef/ZjnuVpPADvYzKyYvGLmMoqeb/da3sqaoq0Rhld7mkvVxv3rIVn2F4p/MliH4lk1+MCtib
DVs1ZcGpQOxdNubltkMhCqDqWi+h5Ln4r04Y/hd0ApGGAWVb0Cw26IeRD/dkYR9l2J8/zzK0MTkp
OnISles/JqwMLW8kKOGbO6IJZR7aCV6tP/dLGSLHgpXiKoO29vpB+3+voGNKPzcw0CPBW+m+n2dX
/oAQiU5ZDrBkAVZLS7JEAjbVJDsR3BhJwN5buW9ddF3zZ7bN5Q66NBNcF5MPjR5G+e4qLYTAkch6
ER+cpWBRVCs8p4F9eRZoNeDkCK5/pYhTERONOsqzwCZLr+cvZs85vY0mbAmtR0vyQCb/rP7KjM/D
8VWWt/Vk+Dr7VCVKsBpNxaUX/xQbH3V7CSD0Aeb4BDdfsy1FJKaQY6ghksum32N8ZV9u9sOpynlW
dTJLHr16JfZr4F7mr2s568L8I/2/L2kkWODKIPOYc56ai8RVxbkU7kbbRhDkgdQpcz2HLTB0dQCP
QOfLKL0co2os0Rp/r4q8NDTinbscSqp8UD9eWBEgeFrat9mkD08i12pdXrWV1F8sb3gk1//9IaPa
gBwE42bpONlvRgPwpPZfsRepBBdgGtC9lMYOBTbXREEWAUwALrZKeOv4BwQRrBKFaUQyleMjsgjm
hP6c1Hsh3siGohLB7sp6BVKh2nxrGKTIlJhDZCKIJITEA69uXarTanbxobbO/FgqPFXFaqQegnGJ
Wq9CmXqsMEp3njkuKnWMoiMQENTmkUb5kAgquEgZWUEEb7qnS0h0z5ME/2zjIRPoKZrVwCM2vhbe
0FYcwUQQHzka5bcj5Ka579xCFs1S5AJVlWTddWIFcYrF0lyqGBE+svAHmNG7RN0m8UYy4NroHMID
fMfj9pWN/KcGg4kSpKiogyxNdyJWtEppKxhqt1ia658HCiaZTIVlGjF7DRd/RejHLwDjeVGGDv2Y
lv8hW96VpvpLmLLvByOGh2iyLSEF/0iibWroxDGEom5LiBV124sgIF2tA+pOwdSMEqJ7TpqwBF/C
ihz8LZKSiRZKWw8dmyybCHV8yir2vZp3f5nbwbuFCTeXNe9FzHR4WZjdEuRW1OS/Ek3A1NYgSvZ9
ZWqTVtX9lnvwHZgsEtxWsazzssCGgt+GyMvVPr64JuEFdaF0dySRAomgXYRwRre3fGiKpdldzvFb
AbaA+9YIk6TfL2A3q1QddEOkh/oOOm9iqRYERECBq6G/8pFM8VBOllIEK7RrkdIqx2zIPvLRNkB+
xdArUos1rwTexj09QZSF53OuTAkNXAlQf36ys1L7/vTGkzwW40tUOOUNBSq3TYmq/5KnIRuj7V+t
sktCZ1oJsHrrtzV4mDa7tXBpUKqV6V532DL5UjiZePxrS5qWd265ri2zvFQIbQxhUXHK1Yo6DBuK
z+Gdx/w+eoPur6k2XGDZs0jej6y6gLwwYvjsIbQ+1VHs37nbd8e3ZWwad/4qaaD9x/use/86FmSu
J+KhzHeqCudgtRdPAOSUtrACR7Y0YHOYrZ364fthJzwQJhu3//ejevnPEuDyE91GAOLxH+S9i9dG
RYNx1YI7npnBZqM1vrMknHDx3JSOiT0UojvmksZL7DnbLH4wQCeXTxkmPBfw/2xVfPCnZTOsYhmg
pwnZNYHkEM2JonDamCqbVO+l3IWIg0JhJutR2tjN2xmDX5e5Oy/x53Mtm2rHj5Jdd1ib+zTqdUsE
R24W84xZszr0YlB2wZSt/P2XZcGXNEk5D6dubM6YPW1O56jdPqhk0E3VuP0yx3YlaZKpLnm5+ihL
bu9p6h7uBSKZVp5OWxS99DTAsPqv8ct/4VfNFX5aUB/VuecAyWyQO9t2WSB9Qlo/v6OUG5URVX6d
1rjQnLF9BAVWdAhb4IRHQ5InZkm0I86swTY95Bil7y3KOuS65FHlTrJknwYR/qBjrOuq73SiVNfS
NFVYkgZDFIsCzAgk4BB813x0Qso7rV8iLNFKYajj5X8xYET5zCoqoHy0VfLx+ZtLVzfuKXr+EAEk
EulCtVfyaGot71k+O0jslSGOj3nmXGTDB8WNt2iHy+g4/EjQduygK+nxfFIijDm6Eg6hax/ubnM3
nFJHxsB4+35Sce+S5gYx8+BEvYRbNtdFbmNtnxBZinsIAeC3Q2e5LiiZWSCFOn78Sa3KCxIKS9mr
Rsjvm8CIWzRUcdkZLyDcAA6e6k1AzOa4m3pdEheJ+PCbspUVd0egRDAHCPIPV72XTvK+TsolpFYP
LMeFeCix0P4aN+02w89FW/gJT7TPFDo3q+nDKpR25680pQgV1CLtV1zmoGIFRdP1eJz+FQ6lS1W+
tjaAMeU1AmKUPLdKqDEb2Zxpz8MqJaq3jgHB6XNbQE543QSFlQQLLj7pltLhxM2nXYaPaVgGeTpt
oH6MbJFODuLDbM5qrhlYsBlI2hyVLKsmsLeD1K8v0oEX3B6lWksYTMvAr9RALEhN46QSQB1EBZIA
Zl/7Fyuci80VfAbc49iBdytbrIc4x8SkNu50bH1UN+vFcBUC/ruImU4YMuJ9PEPdbUqQsqUIPrUI
8gcIFDK1pb3bc0m+bVe9RwVQpKprJhyZh0dTTRdTh5xKZYfSwvQmWcR6w2AJdrudrgZsfypE1SG/
9SScm/e8XN2Bnepw7r6NXZnDhyPX+3Atom2ShTXVL8Khf1FwVjJQwc5DvjOhOqPS+fMi6ktKmRl9
oAy1gKzuwsNBwMthmJN0OZgnxW+jnKHa61ZPU7H7RJQiKJbaBZmdS+ZUNg0nhTTCjGOpHOKDAmKa
DXxnOf3/7M2X4HI+oDtnOFz5hiRVii4Cotf3icVdvLal/un4phnZfrn2+cGRKXZuJu2XbTTd5a51
bKFXIgCA0zhpNauUX0+FRaDUg0RepSuWgymSJnshOZ4SJG6RoLwpE59CKVXyO3cDdTUga0fraLy6
uvDMcniHXyz1xj9QRpyMrJ+x65vopVLXv+DdFa43m+mTwEZJzAjHCfIfxDSYxxCN9Cz8D9JJAB3l
RLMvlztK2g5kpzhsmDa/YUFOayDSvIz2im2k4lpWpCQESUv40QHZN3JMknL1Y+3YWzcJrMPEIcaV
UhUnD5lTNgti4tmT9YhoWhJvZ5O3uFGE38qFTzpFcAv0QL9bLwlUXAzXVOQRGGz9HyZRiHVrbFXo
dBJ41LSf/yIPx4nwzyETTo+KAmvLx1ruyguIARL/hGaW51emm53lEStA9oI8pbGa4nWq+Q7AyG9k
VYwcLZ6J1bL/fsWcVpju+nvkXVl+zjXmr0AqDOpOcdwp0whXi7jqh/tsEywiS+O3Nhrd4siExfVl
oGvV6jRNUrIWiFwldV5Fs/WyK02p6346nsJgzEpF7JBgOeHdmY3TSzS4SyCqg4PZ/PYhk6Fo3V4l
WENsWL73fh7UMd1aNFg3yPkhBecydkZUGgXHZl+zIRn/jVPkH5ytFoFlTJB7Mj2G3R1dhmmpY9gc
B1Lzgjc8U4dIDug8u0kklx8kdN/Y2FFlrxGLhgIlTqq28tRJyeJKoral50T0Ld77Tk6GnM4oNZiF
19IX5Ga4P8BzeTEhE0E+uagvUf1b4Lci21QEnEMltkaMQDYv49Hra8kWVFQq4frXvnP3/efY6adR
CMspH4qkdvBE+22+vwQVMGYgjesxvCGWSALXKqUtZnLBz4wqx4usm6DbquH4d2Z1uCDhqmbQHBts
0k4mMqllxG0+FmPOJt/DhXmrHMhfeN7KKEkGqi+zptBPIOLSA3bip22dRJUvBWR9vKS4bYK/85KF
nkC/n3iA3Z8hPV3BguvW2/QSug7KXm1GNzi3+dpGRFIQfzm61Ih23Tq2uVfQ3NIiuac/iK7QOpWM
RbnXqi7uCIfUxiN4J4SjpNlkWicvM5MUNY2bCQVwJxD5XNLyeo1dZw8mFSWBkr26MKKEA9OCdR6Y
RrTDAfJdbXNfAPO9dCvbTjYWz7av8eWHfcG4iIgF8qwYdtBDz7/gvJuzDKDo8siZ98bPwjzubjlR
T++JHrypCLScGZCkIjJxJlHO029LvWhduungMqIltpDqkyzX3u0ypdeFVhzdtFplEa8iiijNRUov
aHTIWdxLy3DtfYXIGZNLFuQLu6mNrwv+wypWLAKNDQAF7Yrqv9V418cp1WXW9UCF4VUofwYVA7SH
n5nGP5NDag7EwzcST1k6fp679gAqR7i0myy1wBP9FD93bAFupjifZzlwxAG80svTpIP9ej45NfRK
RWnqkXjhUO3AH3yMmIdK4uGJY80r2VVMyF/5jfbko8Nse+/uOExd8wIvBk8zkry3S1zNRx8r5w8V
JBYPoxgIf2wwh1qkIZT3ITOVOZEuyTJNvlTgHWeZIfoMKhK7bArk2qpPM1a2WpowCc+gV+Ste6iN
5lxu1GUZCsyUzzijESnVeQfMFtGDMcj5WfYKTcfvaqnHrke6N4EIzharfeeHzoazIAssfn+1XUio
Pf2ref5QThqaqJBWCjFnXhX8Cd2nu9Fs3akYT0nhvq1e4m9Qouy1DRXQNnncP2XMiRSSQSHKh+Vq
ca7GtrozpafnD1m4y9auRgtF6LEOQq/amOoUD836VFcPMHBZrEHoZ+nR2kqJJpERdHhZYQN3toCD
ACSA+qfqLCY9kz4H4IXGAt759ndLlJzJ8cbz7w3MAulscDotge2NVXAlRct1Z26YlyKqeTWu7Byw
RktIlt7Yrd8JbB11+T+H6Tqw83aZx37KqoJJsuOZKfDMZD6vca7VLmgYlGb5xEvi1RG6w7NX/00A
P2QQ0w54j5WjbMDyyLFTcqFoT77BUytmZV5PhU5UUl2m61V6hYr1U4GlcxE7tGHs+m6GyblHLUbO
U/1kiJXtVQSQWjY1Qx96gM6+gCdj5pqMtEtinUMEcomwO7Tw+KVGkXulLKOmnb4MaNlnJLGpcQK8
uBHBMh9Dvb2EwIHyJZkYskSN+3823N0Re3YtxIuRI9wmSS8FQaEHkDXbCvnEpGJpeVNjgAGIYTlb
s68TqlKpCBlfcSKwAnnRSO09jK0Eku5gnQ/+QnTKajblljD686zTAk5/RegIJ4qJ+VoLm10bxPX3
dokvlhV9ViH+5Iaq+9/C3GAlPNy0sUGY7gRNRTk2IDUIR68hUvh9pr4ueyTGR/jwBUSipZrZ8qFe
C3CydNiduH1r9P2zaUkTlIViwtURCCe9pNmr81bjDn6KXC5aMaO9j0kKBrE7MEEU6vCihKpUzy/T
lxgQzhGE+rzAdIWihhrObyfQWeUNGSLQK5Aaugds3l8xPJdY/Yrld3DIrezuRGN6DdbOmX/Zz4Ju
NDfxB6WMy+SZy0O8T1Q3SSfJu/RGlKdlMGR2Jl+PDiFCMIxLZw2HQhQwm07OC5IbOPyWD9Z1yB63
RDPqT/m5DGTGIImhko0qqNCfLcl92RQscBO9LS6QnQXe16RdOU0nULP3VStOrtq/3p7oJRoE0h1A
v18kbUup1UKPQp9nrpKJfZNVqK4kPKsliqu1J/2oXNHAOOoD+lrlcbW6pwLNw4yUA++zZ1GyuZRw
DT0lcSv3qjUraWcU4BEI0KuvCA6ma9rDhS7Em930ZAtHjN3J9RVvGEeLJ323nK4Yb8L1mtMFEvrH
wz3oP9mugqxQbC0uBXLiOSxc0WJLwzywux3Nz8u4CZAxLLaa9hcw/UyzORTHAmCGXkCRomDG/Zq/
e0+ziEnmN4DoVpMeCHUu4OLcq3J1injLHBaB51Nza8M+XGZSReF2ffT+3XKvR0H2k0iOaB1uJ8VI
k5As7h8zfTnQfrz7ivTOURj5p5KFHHLjg9eWEvZUOs2MWOtR6HZKGyunwD1IxvmSQSpQqwPPIgKs
/LJcLpHRBWXlQrEr4vwwkZZ2FGFjU5KTnZoHdxVlGj/Ixq/CnjE2HhbfpxfON8TQ5WeRJ37a6n9O
rCCNPqRaEt0RsRloLyjf81HRZW5RB244cEYVKHpcdrfzFP6HuKUHdvmL91zAP1rKIQ4uHFw71DKK
Nvxr30sHfJnYsyhJG4BizJElAh0z9Ubfp+uxrEST1q+CzvREwXqgycut4ck6z8kImVIWZWghCQXs
RDap+vo2tmPoqnK4Hqezti2vARLJ0LJQhywN5Bp8slzydIqxu2z8C+2UIPEnmkAzYjlB820ha75M
KiMX8aMEJ0iGKrzarOF2l4h4+4K6FkKgd/u9ojasHba3KwwJAJ0xMDyIr9slf6P2PD0BXZ1Xa6f2
NcL7/s4FcqflJw0Pg3jBky6gzQQZEIY04G5L7g1VgtMtVPaArdf4qCMDppqge1Bav/jt93y5zJqM
wMwf1PyUrf0s9lrVi3d1o5JThomn3LIjHOsBMxXNhlM89jT+p+RNA1Ytsar6gminu41HtX0/wsG6
Pv8DXuPCLAk/4p/kxmpRwEM9+lUm1hPeoCSIpJaKUQKxQEMNEw1qjwBTR4D0Dc4muj1+R7nWcG26
Q6WO1D3U20EjUMyXTp9Io5qjI9ZfIJU2cblZxTmj/TDpmxZaIwBqdtUvbBU7s2APvdoj87NOLJEO
Iiae9CpQEoHIF56q0btozbua28S5HO/0W7xJ1mG5G8YXgCjwfAvlDOdJB4Q0t4G3+W14YhLa58li
xNO6uJ/FeqiTCy0agEQ0u2iQI1Y2N3lKdqchGuF4diK+etZiL0dH0hOBKLY0d2n4yoC3ZE5l3atN
P8OZ9xL17Su5JiwqIHNov0d2/p0vZpCHaNNRXdQh5jFU6eG8L24sHhYTLizTR99Bc88Q2DFvR1tx
7xd3ysIZSoHjJQ5bGFzkMVKpq5f7zua6MZNCmoeXOMFUQxzdhalv7ltP2OCL4duOjXJtrmPSWOBh
OpZm9NNJK8f/UU/dirdkdwMe0Hx3RVVRZ7flswpJAsVHlTDYVjATjn4cfQB5hXjwKwL4fJSJCqhF
Y+KA/ER2izgIDHRPC4E1GZZPsxsECwt3y/va7uZ6Enc4LPm6p/VspGhIyAW9OZofNyfuNYVt6E2B
SG6F3F2oTqUZl8i4e+E/m64PVLKs9IFtLBPbbEVteyAhmLVM2kc/9+KcmzDzsX0cYM/SM748Gc5X
3Vp/712B2oazTlCIgBOqFTps43HsqLbTmsBXWCHQ5VBOWJl9zK1LwIAW64rbb9c4opyDtQcQ8Nk/
yxHTD8KhBDaum53FPj76fvFGMOdQ84oFlSFxM3cQ14BhfypkXDaad4YrKc1N2iDTZrhCrJxCk3Uo
c3q8RMZffuO4moMR2jrqgNVdwHoUNc/GSzV2LH3DoVYmATYVV0n4UZSfCIFkjPzAcyUr1T3PdI7s
7oOmnOhJEC5EuL0lkg3NsO9xP/GlIDt7T8ihCgOnYWME3beAO4RyBqtiZUDg8e0sWN8Ke9Ln7lFp
O8He1nujAkTvAUxucyRFIkxylEF4OM05fXFlckcbN4buwDb1OKl++QRrqT+ks8ePi8CVZL/XgyCM
XhPrbkCUfwpzoFFYhXiLX6NRJmRgS2DH8vuhXW3vGJdEZhUx+s3JkPGP1LFwCPdR9EjXeVfq+0mr
Sz4zIQHfgkLQLPs9YPAcT0ywfsPgZHnbSjRDovkRDMAEfJ4+2wsLidjg3cKwGhj2Wu5uD6Ll7HxO
fZ5KJwGa9Xng5+33xZn+1Cd4gdAh19K3EkWTWCcccI/VdRa+SKfK0lwB89CjISoDKvxzqiFZSPqD
tYd8aWX7YIGfTQhevWgSQpR083Ba52VFaIEGc9avM0QJhqgbwf5qzLmnX1PbJsY4kl3FejEuux1b
unDIOINyIIaiETt3pZ8zHUHzpDpJ+p0yXKp49fkpoO0D2+oioI+TGNtmta7+CXhkqCm3mKrC+GC+
eFNOj4ZTQQiv+n7ZByFpXS6wcsnxC6qeS2g0KyWZDWTJPZsVNl7puK5m86FqxsueTUF6h1KHY/yi
s4XHe/qpleJrS8Ef5aT5qTgiB+GmYPympXd0C99/8o+5x99d032LR7kp/aIvRbTQrcEnAib/28qP
4Gjv7HexbUvWgtwEPRv/r4hAG1ZQmOSFGPQ6ZIFfYt6OrUkthsz0d0xtOSy3iaBbmqGnU7lEvc3j
ADawzy2Tj4QH1LZl3jAxCykE1kWvlGao3FVjGqFM8p8zY4jb9brHyRw8HM03mqZiFifgZRa+Va88
AxIttY4c5WYIUSjEcwvGl6OL3ZmBB2HJTPxIZ2W/mA5dTzGx3adK1d8B1Qy5NqRPrdRLSxg2ENS6
JwzKAjcQzN0ACns3OcK+1SqkeKwKXnsU/LWEF9BXGEiR8gmXzPbv6T/L97OnYRE6UQWKs64hZl4c
5waBycek7tMZIEEeSzfz28DUUKGmOt2ZBSA9MNQCaw9zFfiGTWs++SNmVjOesll/cFUezP2TSPd/
7t0kdAXP3Uz5ohZn2N1rAoIX5ClNEkn0zLs88N1TaKsNp5jIXxQEtF7zYfJI2gps4AnMf6IKDUGN
V6ODC3mxWoFSo36GenmgOO//Z40nfeSyD/oi8v/vEnYntnUHdU18vImPUmSwO85W+GJzxznGmw6u
jE5KgnEh3+dZ87xN7uRrRd/8bsh9oyYJ8KLauQ9x93mxBl6e+7kFZcHka1IOtyKWui/we1DcEU2C
Bd2ch2+LO8cJFGUD7zMKys2Bzkb8VAqW7iIVi/aS+ceVzsLXFY1nlSqJ4qoSAqW+qeTcq8V4mRhV
ZtH4UvwD9PLkPsC1CTrUfF+y2frx/duh9jVt4EZQWjoxbeSOhzKZctTg/mwel09Z2b1VRN0aP+Cd
WNBf/0X705AkiLFidDjHUhRPMsyslT7ndEix2S5SwpAoUAhA7ww45JiM659yMfiHhpbbV1kPJn9w
L65ZbRtMoA/6/61gGed3ZMCk65zoMdL8muMbco4bM6f0d6iKpfbhjnm+RIXOIxV7s9rhN5JUery/
uwUXMwqK9W1GRwkehd5a6f9XeZ5lK/wVt+VNNcc/Nee133jrghpz2vaUdkwHI7Pac/aR36islOYL
GsomKPqIRrBuenKh2jOMmdHmue6Ux/PWNeV9mbPqDeUp6dcyRJ22/Lci8gAMfEIUrIMyw4iDIAb4
t2cxtoCzR7LcjfEoD8a5+Il6SRTp1FuYFmEIpEfO4uhH3HFf7qpkg4J1xAU16pbkvYdgS4C3BreB
QIndFBqrns/+BvzskJSIwamPK6rKKEWChyd/6EEXWGvPMferMTnC4lPSDZRxOgWN6e5Qmn0Pzn9N
JFiooz2QhD4qHiPxNDbF5uEDdd6z4FNGtcWd/i2p1l1vYeqab1p9mth0PFs4HTcHohgZGn9JOEfY
+tD7RO9TpqCxwE1zQpBlmkHtwdI0KtX0DUWIVaT40TjXS0RX3SuY7lp8kPrrgjLMi5hci1GZr/fT
MtWYQUo7VNHfL0NUVBc+Bm5h6pnaKsSt4RZ3txje7UoUeNW/Oo1pKjsPG4pLoB1iVtwU9Tf97q9E
RQ5XuCjCbifZC9k/4NdFYQMhg3RUXns/FkUMXHQOe+QFqEcpHmUIl121bfRefn87SLUV/i++ZX+8
QJcWLKEW1bKxJu8W5jnrsuSC4BKCCLHThWcInuiLjOaY9dJAxTwPwvSQlOwQSHF2xBzfwvJ08dVm
PmcS0tqUOrLGnIkiviNI6k8/Jrl6otlJHRpEqNjX6JiE4GhvtxJUCn0BezYywpKf7nMWgJBNK9/R
TO8LybMiqiYw4t/iDeDGCyI35q427eMKyu5+LzyGuUDLFXPKOoKgI+HJPHkqiV02bx6NHKEe7BW5
SF41966Oxx0kXWINJj47/JRuRhZfhlnaMX+QxA8pRBMubQNJD9wSMSpdkTJdn42H1FMP7yt6iiOm
qvU3ItgnsOePVVw09i6iXOnuX9vK+Qe74Fgbr/eZerv5LbB5mDDuPmhbOTjS7Pmyj1yiHkUi6PMg
TTlRg39klqKpr+Pp4kkQHuYxcitF5KGX+R7U45OKeo620Dv62s0qQ2MvcRuaqOaPTlsu2PvH3Qf9
rKpYFKyP6FJ4p0O9uJSWbNTpcPgZb2jfzOMMtabbuUBOSramQu4RQwqNwoncItcBs6n9/hMmizhG
iXA4UmAv2Vqb/Wh3wewzL1x7K1Kqyge/9WpISRoap9CVUSVJpLsLOCDECOCwi31842gyMf+81hJk
hlxNgeOi6JiKkipFNYDcZgBhiWkW34ZPSXTl2YBJ6wTMNrRtqjEL3rJ3u3v9e4+7X4Tp12rB+ogw
JFHY8PXkkAtjF5mSxhMosVN/F6STsGAYzu7kyrzZpY5JPpGo3Lzc2W/7t4uoJPlOmybr6zZYmOHb
ywlABbhOoTN2OU0X0j/8UAJSilTs6kTpD2EjVUYl2HZXcZXCW+gUJYJYtAE5dM8VK7KYJtnrkvIj
06jZ/8tDdBjfEY2cOtlw9XNrrezVqUFjD+YQ4sL+g+hdqdcPF8s9GqcsEoUd1ThB6Ig/3GwlFRBD
dBumTZ+E2FeNDo6LW2Ps4iGhQEaKtw+kCF7qroQZZxdbQUgWydkVz+5HJJNkuzJk8gXf8Tt3/ckF
FtF7lS8E0gvQ4FxyLptjx/BvQknv/VjDq2kKHDhFeVjQu20wWjJq6hk2Ii2qngZFNKKsOsjTiX5h
OtC8WnQL+0OPqNFejmVKeGZUpbu8rVipWx3V+mZcZ9FYerRJmqtv5GMn0h5xQmexkA+q0/QG3dUA
ceSkMym+w/dJuL8FVMwdR12W6EGteR6LJSf5+RmOipOb6U+IGhFZYKup1weBkNMF/hgmo3aYx7Ua
Ml7qFNdp2EXWJ9mq8XPWmrWOb37q7VbhY1jm2S4WvilqO14t2GZ0/9+0f6kAKuHmTC7SMkKMfunz
Oev8hywSMYdfBfutPsh7LfU2ahzgklAkJXeVk/PHn08KBSETnGHPQUEo6XUEbHzxLMZ5XAPo02kd
OyMYd2s2AoD8nbzIfr+lqoItsgNut4Z23OsEVEE2MasKzccj6Q2X/7ugPtDvPytjLmScxwiObhL7
uoyVUxYX+rikIvLenvYTvmuLDqYr/U+m6j2TbHllZ0hYmCBvFVofWq50mdleTB0wAYXLBLNmV7An
63DZGt+m9pExz3c3EbenTsDSzxSaospKujWaIiJDc47SQ+8VG3knZLZ8BzOgIO5xYWQT8r0axrM7
3RE1omlZrjLcm0pcHDkTZEx0baLoeKYzcqzAno1VwH/QPQloMkODKlHUvl+Iwz4tfkIJxrjOlXVb
S/rKAidvTbG2yi9lHtRz5PeeaT202qZIIRnjI7DkuQUQmtan9lwmN41qmGIN0hU4qqaHMoEEpGPu
aNLoqxC8E5xIEK3qTTW361/jNIpJv/iL044sjWAFfjhjHxSNlVD03R/pU9j0AezNQGo+Ra9ZxKXc
f5nEP9ed2TEm4BnZZQy5/pNbpBT4Y69ZMcT5DZqbhETAcKArRzMRyOF3vTCanwbnCVo/vzHvTvjQ
zcWdHxGr0LZYaBblIKYDXhQZan4z+kFNmB6WYrP8Pl/ydm8ZDrZW3GRXFGVoef73nkMqbt2jCc3e
okd0Y5fBiBpz78dTMRRrpVTNYetciAMpZvmJ+PqQpEjKyds4bsZgtNkaOGkS+71GxVYgwXnUZHEW
o5+QFaNzxtbmEUTaZ3bRxkrQE1xgXvUeEnF6d0k3XoOgSmqD/GE7JjmgXtpnbK5BPEe/WgmO7Dkf
53taI6sC8CScTKo1jJKFFpplPK2MU2Evv7lbZJ8AYDPTu6X28NjO3IviLgJwC2FBqTcVYc4Oju+2
clv8gRSYJEK5BjC1OWRMWxX2SbV5tp9AIlDHtmptUvA58y12wFTrZdiQEG6h9dCAaWh/1Iw3g7Bg
rKZXkxThkBIwdFBcZK/9B1bpQXG4fEMOZx49k6j2ZbaoUYLfe/HVCv5cVdSrNnvny91Sh41v24aG
HWpFFwJbYXbug5CHwoOt8RM1AJtnfXYxmOaLVMmARWTjFiEjzvHMDrPsaqYgn4SoDSjGR4JxGc7D
gjoUQO4PDjLn+/u7V3yQKi5vpNnlV2Nr3wZ7zITFAbxV2V1P+sL9H1orlbP1hJXsV3RVA+afPhH8
E3O8v9od8lCZJCMCvIzUiobUbmBCtwIUvhygPxX8vl0woPaAv6tNANImmlK1wktulM1owxf+d2ho
+nvUcfuVQHwXX4hB5tzYC1jN0yOtI5VEgvUs9irsKcvxPQcypg1QgFqBdHnPqTunRX5sfcOhHQks
qOsp34TM2saFyfOk9naitnDkOn7aHdT7ypTPc8f8mKRzqo+aAtEA+TH59KbZpRKvYv7m0FxQsd1K
bhcQw5I+200jXYsddGJfsHABXkN2pO965O8t12PwSAbQWLTT9lIjUCmA7EoxhHqO4TRG/mqSyRnY
IJJm26Erp+6AEaUOWlNBo7fDCjtVL6VSwD2SGF2F4pCyDjAhp9O4JX7XFl0ygw2yQCivzbzNEeD3
+z6r968vVRpR2IeWr54rx/Oq/9CEuWRMzArgO5kbw/SHaHEgcIjhNANz5zmf0j5ZAjaQRqgFAu1F
z4KS0yh56LkqL4n31TjspZ25gIcQf6ehGgLlbAyKKiPoGUu7WdQViT8o5qKp/ow5aDY8aiSXVqY3
LmN5At726U7XPwKzOqkUlYyhgGImItE9mQDl7mCOTzoSBATuoQo6KSN3uU5p+pEx2JM8AIMKj930
XKmMOvXL4N5q5ZZl4Qc2Qm+hE1+4nxtJIxuVSDxdE+r2EEbVA4hD03D4DYjGrwZvLBmOEBOUHLaC
fWpbsPnwLbyI0Xw84ofZFMpRW3hLB3ziOgY7euVdqKWPIM7yHp4sbzzsQdgz6VlYrQCUhK9adLZt
laSMxeSaMZ3rJqjN+vi89qW4uUGEcpjI8gKEK6OMXWx8ZxBjyt9mbSOCCLXoLL7weN4DLFOYYoI5
jZigVNaa7hf43cJStfub7k0pdQeJpBg5cSrdLu6OSquR/1s+nhARXLbiY3XvDgJzdBB3XZy4LcMM
0bQAOUVEyM/mcT0HeRYc+D6M2/wmMte3adERkMu3eKJxVywXURuySYtozPC/vQ2EaJQkdGkileal
6FRWrJ5g9rcFSsYciZRmAsL3KCFhFFuRttayl92TQ3iPBk/EgMRkjFcWn2wukA2JhyU9y4pJd98K
GO7VT08EixnOO7uu8dWlUfZkVnaiE6eP+ommM47sCUs7V7I2Kn+5GlnCZ039GMHzlKzYaGeOOfcA
W0sGCCldGwRye7snIcA6AfdgtBLknSh7pzeSDwRJpGhv++Bzx/PPLLhXf+ms4YRqe85fooLdUhvz
pNHeNWJXY1Kup795+ji8qVisjwVe3rMHejIdTciLXBYkzdSYN4/uRpa3djzek9Uxcs6Ht8l8UQ63
Cb1PVCyf9Ue3OgQDK9wPNLAkeDtSb5yAXoU5zlRFtseJOR7O5JF8LGU1fE8hAvOFqkCb7Tw4CObv
twwfk4uOJbtGpVq4mrt/KdtHkl3wGOAXhMiUWxOhqIysaGKmVwWgJ2q6RB/78jPAWZ+GPcJGlouJ
K+RDAJUuUKC5TT3Dx9gMUng02M9RMRel4+h/XhmnCsNdJnWS5vmwb0wBXPHuMY0B7kwINGvopYLK
0cspI8bw5JG+L78SQxU68Fogln7GZeIfiK3+2+TTZ5NfoMyNpF9rAjUe6icOj00WJScHC6pvu6Yj
5BysbHDPS/SQ+LE2c2XCXhC/MC0Vp7L8L5yJSwrQGlSls59AIVs+yDsgx9gCD+N3LQTKxsnney5J
bU4DiAb+6jDlx6cpkR8RdkvG7/w/ICBczB5l+UT0TyT3tAZhgDYqfm0NfCILjPa0zq8qoMfQZ7HD
MTTBCOgqJMR0lvrzvyUs+hlLYPrJ9cAC9P1C1xHA9faWOVUqda5Kw+WP2tL8begKg/u5qZHEqd3V
6WRMGrgnzGYC8VOT2DLPAckgwa+5+1uavMQtbLP1iZzgw4/krjk+Pma1Zu5AC98SGm5LbNetHJNq
7kLpOrb5JbOFeBNNdggpMUrNCuM6pzfXIqW1Ww2E2R+25upl6QWI3ciE9PEF1hoC/QVfS/FFAYZp
DF8c0XOHAWQRQrGEMFdMo3eY0+7YdXYkMpf/ivcMncLMNa/U93zRFWPLPs86sZw+wlvy7NqQn3e+
ADznteRwEgJl6oz15Rr+P3EibTE8o8eQUOmj4iUyaEEjBAXOcQt3nvSOyHI+AtQs0YWVoxovdHg7
/AZZsvDGRZeOzCcjuU1MJNqOGayxqC8OCT4XOkrs/GEUHmq0mZQ90X7hUtmFvQNC4toGqRaNJghb
HTbjOPzQ0buoohtTPDothjNVUpQPocsIkSklmiEpza49GsCMEsYHPrXlvHuY0vdshgzgVR2KCQcw
1c+1vLywSYByXdsqy+Hd5zJAC7Ua7Du+sflYAo1Ntnst6OQt1B63RFcbnWG6j4y5+LrtCaXW1GsP
FXmTWIHtEX9iGbwBCHosAzgecOxAsWmxxOp7isWAkHXBhNWcZh0Cw0MLpxvT3JUhHC8SIIoZSob0
v9G3Uuu9WsjgwfHyNHhiyhSizFarOcNUsDjAXUzjYU7X6R9wbK6u/qVYu7Oh0hNHSwpX1G2E2VkL
p0tJFcXZkvKnx4RmIxkUDhGrhDVETDm9r/M3WoWzpbvwA9A652APephp/SbhNT6eRlDUNKLCeGdN
1wUEAwGdX9ERqvB543KHwLktkTHy7douykgyUYg5r2uvaxB9/8GoLYAyNyoJShtBXwRKXYqG6qgH
4gVd7+eYHcDHUvhlh5xQL3Th6rtsTHHtNKPbMuQGzoA3hBkU8SQB562iz9zKHkurfyRBvsSKO2XX
DM9odLmBEz7hwRA3cJRKwT1P4Ifl9e4b2MT8dbqsdUc1FSzXcx9u5jrpVvcZL3f7ptSFS0Yd3sPc
l8bsyB7dcbTpSzcJkQ/ZLRXxNg6/Kr7PMwr7QDiIZA/K6RoES6gvkpsOb58BRxBqJWoGkEVcQa9V
sdLLc/YLoWNr/VzAMzNiU+CRMV47J3ebx9k3ZrYDeP30KawuMtWGlRpDY9rFvfZ/LRoYHo/d5fgO
2yMKhXuJNBgDqJXXVP42Se463Dse8RD8VozUQCg23lwBoZTlEdl8nAb45X5xD2clqFlciUC6Jc4K
CNKqi7xmPo1kmdyWSfutzXmKMcJHbD87wiJPMpsM3aMTM/5UMWnxsBKTenqCXeZvAQzyw6LPyQz8
Vx2X5VaxoILT8ZOQHTyonUBx3pyVFNZneho6PJkKr7fageWHpVmnNRl9tEqVfe3DpJ+SRYt6XF4s
TKKv/FF1Tobv1Z27FuFBQyS4LBC9kIpM9Icb3kGexjw0xdz2d6m0QiYy7dRgfHbIeedIBcmGyi0S
PCnvrls2/GtOUHUa/nlVsQcHWE/bYKkq3wy1VL7shNEIBkvyyNs7eZLvVvJRx07lz1+UadDQf3OU
gde8v/28hQPKKoTb72hI/LyzJrGUMQnCJmJK1x36GZTjI0eFN4i+cH+3mKjAFLyScS2GanpnvRG8
R8gkqnEBM4GE4qDlwPyJKjv8/J5a7Ky+HHKlcOVoImxAFNDEYDb2YecXNP3XvwOqU0eHRFDid8Xr
4/MG5spRKJeDUEk8d0+oGVGygGvvDpZV4bliT7Vh2hZVOZQCsnPcO57G2hCGLHatH1TCd5W2wmdy
QRKbW6LI5oC27P+X/QQWG7ekJmPI+Fvv1TVECqR2s3YZlSd3IgN7MkF01LtvaHA6KG+GmkRRbFdM
bYQBX1AXOvZeV+GiIHUKwCKP0sdCD61FMczx7aJbzYx59SHhXnMfjGHwhLbmmxUmonxBuhb9NgXx
1VI/OawwlFNbcO2yElinmmVlrzK9zmzqQ3hhLztPKYz8OVlBEmEbCc7jdGwoaN9PL46agzwiL2xE
QA6rf7e0z1Dztc0s2zyWdqEFndduPR/FV/npK1Phq5XDzwbYRittxRWfMO9blpFUeIUJEZla/HU1
V3OcQ302G6IzGdima8h3yjO9NmHuC79ULbQ2/TCmsu6Oz6lirOXlbM6OICI9eN4qAyoZunBfZY5C
r35Oj64crZeqrF8Fw85OhR0/MbNnMwNeiGm71HSMIS2tXWDliP56oGSJ7rW5oZKw2eyd9olec4LI
ODT0CTg9I3XlftCX/BwlnjT9hq0J9XA1mbzx+TYNJSP1Sb0pXO1y33zMRwU0ds85jOlWAIgtCJVE
qQrhBWcz7R8seHMDHGepeInsYdT7FkuWOGb09MYZ1/b1WYW1SLcQMZ/JpD0QXNLbKz9jDGChCz4s
LEJeCNNIgoljLGnZsaz2aNZXhmQTo0nTkXj5o2nlzf+a/9//EaOM4O5q649BjxjIqjxePRTt9HSx
cdJ2qR79XDp5xp3S3yB3BoPAne5o6vCH+iyYhsJpFTVacAiWVOYV++OQU/I2hL7hiUVVtgvu99Ke
2Wz8vLGXYXqmj0Uh9EmQ52yS2HhRwN6LGMZ3AEqbn+pfFRSU4PD8jRLnjJOM2XwOm/Lvq9v/bqqd
aq0oWvwkYcITZV2+fotS/Z5U3WvrOJyb+Z4SKB5XJPT9qEYKGTbkVZYEhqPY5XRiFItdbRemkfcC
t8DYFDtyHLS0GB8Qa478wmwumwNxYFz8REJawayKEYi+DbjC+/kvu8YKQLjj6jUXR+7pzES+xoqd
1mWH/YThpnl0kbaPH7bQG/jXKG7u7m23s2wFQrramh6MqZu21r/V5ED8IgcGnS7vRESEgEsEZXR/
Kf+scenaKAJJ0+UogaCcMDsP2mkV1k7fF0iFDZLh2YAiWOGTNFrsRPbqxCp1vGaMwVsTHAoyyLvQ
d0TgVfPdC5SrTC81ASPb7UxnN2LsQ3dOM/YxQDzpz/zkXYrQ7OtAZbwKXNrlM5P1ZVduuRx3jppI
mrKTLoLkopkcBIvMa6skNzpbycHK2nv6YbzzTccOCx3jXdFr9zHm16ec05VSUIi0OzVgBNjmxuo1
GlRa5Ulf9nb/I6PRvHLxMyRARydo9DuGyQHzAt8Yt2gumTAghZWHNcKJ6zgtQECbikieu+iVpHHd
CokOgHLO+B3dEaPE42lBrVhHA5bETyNszIdXQlbVGeob6qqC7XDJTRKc8VyhVnulPwevGitgsBv3
qOqSy3t8Rq/HQu3oUBNsDEHCDoapExOpx2Qukg1i+twsTsdZqtHNu0w/SWrYMUROZvM1K4qhRMk3
oQybKzgElmjk/LG+H5jhbI+D7HWkmlvRltZooM7mQpoVRLS5RGY/cHD3PMrP2xp60jZVEk05i4F+
sATlKAAdU1jtQuSZgx/gcw/VKiC7wHUz7af5cJqTqRG2X0EQaQyMRKhxEeV6+QA3x0GyTwHD3HHt
EFrp2sOoAz/oFJs031cknZC31jNmFmkjxEzVStJKWFKEwFW9H41BWLvJRa3lgmo7nPrxXNoa4wF3
L6QeNtF8E53e7+QOxsCdS23bD9k3Lpfl0n+gemiJoiOaP7BPpivCWZs0/Hk44uKBkK7v/bVYcm31
EmxxM+T1aKzDHA9iVFT4DI0xyEz/fiZYj+tNDWHaqsbyyKDD4Ibi0Pic7SEhd3Dx+P/bMr+YFJrz
S434AmZ8DMLL1/GBv3FmbHo1SdTU9Kc2YKl0HXoSaQV7ANQDKWyfyNkD2dPm3mGpfZ6HXTMiQBiO
PmFAHSXS5W9aoAJ439zDXEzRvtTBneO9Ko+cUZhyXB63EhErAr58yrMhLpSspeyJGU/2V57dF1Z1
b1TVBzi8gP2GhXNKjR20e5h3/Dl34G0c+9mE51YWcPn857Blefld+76RAFUc0Or48mwniI/2fBCN
N5lVVWR2c1IjzVw5Ypxo9vKViimmPTfBd0MXiCazEY9rC7dFjXE7RFosJAWTpgBLYt7zlz1KOzKO
zc6jihnClazOk5uyCny2nkdCQmgrKJmnFsnqByrVFwHCWB4oZOZkaJ6jdnta1IRppfQVsdTX/txl
eLDm56nAJIeRFSvzYeGNZ0+7VECDGiLOtalJj9HndngfC8y2NBn9yHi1hhhjCOzdhFOckKmCq7fg
EShOnMWsmLG/Ry7fhqvaKqBatLdtvpJj3/BFJs36xqdKmPv049aRBvrDEozI50CakdFUl4Y9Ry3l
YIKlIokYJt4SLixC5I/Z4SA+eDyJcSWT8S4iBNnkWJR/ET6MvS19I04sAXJAwMkO4+Gja9dWjuJm
PR1WfvGSyvpMNCDRt01vOwBggrwdrgQrOnoCD3m3jNqYrtYZ4tAQmRjwWfY98ccW5hliCskblNma
puP14uL2heH2SUAm1PcKe2rRDx5huIe4H1hLUuza49Li1dxHS+k4zJK4bpOJyGMXZiVlL4MSTimF
GxX74o70lZwPHALrApWGD6xYPiCnDnrhHKuk1NrCzTStw1HU/ZxiuZY9ULNtUAscxbYR3EQ2msag
vvD1xAJt2sFEgVF96FVZf3ZtIxlTWq7T4VKTru1GiS+k//l5vqzQznOdfIB90egKAMxsBkYBG1NQ
IeHYpukN6wSZLEJxYd4eCngWiX4RFQw0+ZjNpfH34G4mbOS9DiNTjl2wplbZtCuSKAp/YPQ/jjdy
DQJAkv8u7gN8ivM+GSaK90fHE5CImRLW7mhsXa6xEnMAHhsOU8/XmApbpVyrpo9AOZXq7MpIRHvB
I9+6Nn8ikB/THaHSj+nGMjPzqlnTGP96NLYhc8Ufx6EI+weTd2JLD9RC6BEMTCqtfjzQSzM58zJU
DpeXy1FCKRom2iSRZbrLlmu8csRrpLjWgXqh3CPIRNLNQALPPETG26Aza3XugC2xiABHp6JNPyLE
SscvsBhwdjbpjRYoZQ87sByzqH30hjlB3Y30dKgVal/OSQ3iiKokDYdv9Bof0vWBf/7Zy6z0gEdA
QG+21k6YnL69r+Kitdqt6eRKhq/m8E7seyQOWvSLMcjocVnjfhgWcJRD49cxU3scVIkpLKAR0LRi
jPONf20svajBdf/e3YloFJHvo9H0ofrFoC/JTepJqBw9p3aWaKDiX4YBK9pszxHHjxBkv6/YmToV
akJM7UAn2221zRwlVRuVxQua/lZMUEdrRg4tgn/ZDL56pfFWO1ecyzpvO1AKpRs2lD0LtGq+Pam/
s5hqWOfCll8xqavmqf5f2zrLiZs4xit8REDcdr47VCSP1nTWxthxuPH84Dnzlm9FTOYRdmC1HqkM
/EIYCY+vsl9ms9g6lVoi4V7OgZUcZNnqChDyzxVh7O3AmTVQ/PJY0PlbrPVwFtA8r1zNLg7N/oF9
NrY3O25+U7006Fqfw6DJB3J5ZRWL6zJdabF0FMbZsQ8Q5Ti//fHcgdc1owTqHczRrmamBs+FNMUg
xgDirOBOchkFLDINpdNypPS8Fi6BraXgtLUJIjI/z4V1sGOhYqO4iNpauWpMnPPbmM62yJkJeB1a
aA9Qp2DRK7JNkdSaj4TH8rqLZvFg+Din1/mrvNeLI5iuyMVOunwlXXUilt/rIhHyAECiMJxsgRf5
aDVXG+959C4nT5Hxg/gmT1gpGvmsHFo8o6ENujMo9Ab8KhpTXrfrlRfHIujoSR3NO7aLlinE3xdb
dA2yf0l4ty4NwaSVjDjcc+OUj500JJJ57gBzHFPScENmzD4s1KdYj3Gfgn4cXP1ut8giYgTKVz8u
rWZgUAURfM3EeDxYDQ3XrVk4Bb8P3YSAWwK3DbGaW0AEduj87qxyocSxiS9CBCzGsPftgNHmHhlw
tSaSatN1SOIGP/DTG09Eii2fU8ymYWmiv3zCTAyx91H1mqxFdthRcq2Zp1z+xzAP42iL7YWLvx5C
b4wwZZnd2+srdlMzm6X9G9NmRnN+MrYMUn2lo7jo0rHlQ+rl53nNQm6C3hSyyxr3NVTwPE+80chD
3Jp/29VS6G1omBqJaYY9FBMUxfbwKkumwHjTlM8l7Y2wR+d/2uzuUgkMAMVM9s1spKU1IaBI/gDR
bMkoDw5UE0TSLfGNOvfevgMNgywXwAGlDN3EoIBAJgbqn7+1Erul0LkC+T41SSeSpnmVg/A21Xql
kir3X+Ht+3lA/959Uk7YD71D6Wm2aUCXRFK9ZRzcpb5/6OgIZnui4O2qnhBxWTTBKBtEg6CrAYHe
1Vpq1BOKYoUH6Z1Tq208KDGoHD21pHMyS6wgJMu4qAZkWBzLJtaFr3M81UYQkc4ZDvCmadUi6p7B
Dp1aRIPVTSazv+lmudEMS73je3p3rkwijKmnM7ehnA82lV4GJ72oEi7hRfVF1v/ZVuQM5ROOJ3sQ
VjyRKHctsGZyyX6CXALe9e1GM82Zsc+Pio+AQNz2CLW01/28HQmiW+fAea0pHXblDhho3J2BGOUJ
4KprGRDro9hZMOECGz/LhqxJgaqGDLHT7FiycLyUQlslizNums0gkdkK8VheJ4SeMBcIK59SKqpG
9nqfqZ4eNA5FL3s9zbmmuhCgsVijbulGc5tqKxYdC/HIoLhMrQJSnRyXMGsswwdGtOUi1//GGRLy
9GJ9N9hgEbQwPx18ncsimy9XZsx1Tw4gwb212aN4fll5VmKbMX8CQULJt6ZAzaOi0Gbf61lvi1zJ
9i47CFdjfhtcPwG/WjfZ8KvStM5QmchJGImb6gZ657v0ZsBMVfOIKfoy6Wnoae6s+ZTxwCbxMSpg
W8C3ujzQmTzjxi6V2JXE9CVf8ycinvKscnWdUi8wm5oi74lAD9qN7WdI6NfYS7/IwOwc46etUGFV
oYdz28QndIriptVP5WVflU8WcLlRdQUERoTu5ed+PycSEYvBifeqkfQnw9XRdKFeI6+M1GWQ2kQ2
zsrJqofRSUa9mlLGXJJYer7N8V/VBSGVhgbaQOwU+zHP5Z4MMRGEAVoC3lWcFvbjcKsdx4MCCH5Y
QKyLXJw/tbRIvf0zBpSwwIMOhwQeOr4cBG2EJUo+eoKx2wm9ylCe+o3QkjRGAi/RJj4ggPZga0zb
+1w0apeoGH6z03pbhBh/E1Bgyweahm2ktTNICC0fZqfEbDREwaRV2uSToEHiyRMJgRl6X0xfHMSC
yBIGpF6i2jKyb8kW4IM5+F8lRoE3LSUUc9rqP4B7hW2+vJQpmFhmKWL/i7eiqqgQnKz2tyHO/Xwt
skpwXYGf/yuz3pxvjyjYPkL6YiIJEKXO3lt3eedGsWVq07chqgrntkV/YKlRWRa854NyUdtmBNAW
ca5Jz1RkQmSXcgku2RhSgqqAtDKpvkimn9B7f8+pu2Cfyqz3j2l6lyFTPBBLWamg+QEMfeBeFySA
GT9ojNpYHXMub+JLEyZ5WtRxra7AoKaanFiZol/E7B/GvkbYpn2bBIJBSwP/eyZP7HgRlcL015wY
xYJ04cXS3sy6VYKAxKSMKw+WzZEsQkO93Oedq105ccAeGqccPq27CQ0mtQMGJqJWZy59G5G7ONYw
Q/2DTmQ0Iovs7j45eLex5P+rJXyJ6HNzhjhqXNfgF6RVBLQ7zeYgQ7kus+K9PnmwWPzCNNCCm3mN
0y2WEBHbyiqpRL83WyrFDMp4I+sKm8mlox5y6+mUtYrTomut96WhzYsMu/MDwvLF+AN+4GbA9VNL
HJwAN3cLLbYjnFaYzJ7TBI6Oa9p7rQabi24cWxipVFhp0hjnPe5UD/MKuaeX/8+O9zJH1jES8InF
+N+LxxfjIO+d4B4ee+osL48jT8zZVQgv2Jo44t2Gf5Na2dEUe3Bz2OIyVIjQCbo6g7lADObBz+8I
HftZi3fkJubWRzLBiMa4PWmS9VAnxZ+ZfZoDFBfP4OOSmbB5j6IfVz0yElMRidJUAoqmv0mt7nkz
n3X8G5G3HvjzRiQ/O/5R7ZrdwbR22vsE3WKKyrXPxzatlLd90tplogfdHRKoR9iJ1K56QCK0Jz6K
PNG8ArX2f2LFQAvVDE2NgSnAllnG+1WApaOnaco7LfQsXNVbgA3CmfkAsuq2fKbWLNcupNK/GM/V
9JvTRidpxFSMbTLda48qdJGyHn1f0AUnHrjZmeiIRs43+J7y9FSoLtJtnnZR+KJZb4Y4hRMwxJGQ
nDwqNHXCaDT0mPr3G5lCNxROe/0Um66c6nG/4DlhEHI6cV1rZnS1NkdS+P5oMK+cbCnFhfXI2ftz
5i9Qghd08AQS1Bw1cYRBjFIc8YXKVrLojeX9zh/JOYKHj6RgtE3kuNwHK8a05rdD15+uEBqxeCmg
gUzC1rAK5gnTs4l3T4wgFmLMO5l/Aye04idC6w9oQUXI1jbUvRXV92rTEhRieXH0P6Qf9142sX0R
8/o2S0Tzy0ppht3jMyV7Xmpa3PVauXYHiXb8gQ5NSHC4+lw+xvjzUthZyoat1hvZge6xJUMYPVkB
0q9SMQz5GTmkSoi9MDZf132Y8UdR6KTwm03+x5tppULA/JBchXwDHD9BLBDmhP97vW50eg/Ndmlh
Cm5YQHPj6r4Rv/QP6YqkawPsINEqSmhUvpWM4sM7RNzABoZIubBbGaUX4oG//pcdKlW/2UspIAPB
sVOt0ChwE9IBYX+ePGoyQJMZS3o3bhUvixG14hU/bQ8q4FTOiOYHjYYzUPokNDLgHCEfnDq1nDD1
eTEKU6RGyGYZp/+M+angIgKWJ7GeD98AKxD99+4rG+O00gIkiCDu9GRExbCXVUUKr2dg2JC+Jy5K
/gz3MdTEhX19ol/9SRaCbuMf7p7IE+AMLfMLeeLRKiNF7vB9q2kcpHdIUltNTTyrovmgAsOkIbUG
mGHp4vAjEgFlpAZmmDaEd/Bgl1dN6UidfWs337YJrq5kG9G23h/Ny08kKvvzm6MteeYPqS2hBVHY
zbLJ5NGpjZLeWsqX+20tIZQ0WACPiCPeTho6sfarLIEvrWKqh0AH/CmqEDrhEn7DJZuotDVa+4cq
VflmFCt9klgAcp7g2YmJSUKyTJRxCP2IwVd08ZOEwhYgv5NX1QsVhYDWwD0VuIf7midOAuOsok4m
Hau1mF6ck3SsiksLlEFnn50VNv76rCLc5pDxiJObDQ9bR1epgX7zxRDlXe9vPcHrLS5mkBc0yOXM
8POHr5GZE/8NoujeDbqdnFpi6NyUZGRe6bQJ6WPI3LxsTALX7OllpYNaLHTi97hIaEaVGZ0mxMPo
dJminj93MgssUJOwOSGphu2jXAsZ/E3l4uRrahh8OM+9x25+3HO/tEwDBbadei4r94psF3vu2FPX
Rb5PMVWc4sUExpeuK7z+ABRNLjhhExXZEmCs2qYH6SrVIUMA2lVwnFaMLOxV62T3o4eLFAwlAl8i
n1A0mYMI1UfEwlnxwFUyxktl8gHPl9/S82DaK64DAiMTvwahLq3HAfVz4FkHRPaP/eMS75b2TNaQ
yf8G0vN1nH7G6wGcHUlWPHPfLusgjkvdrQLUcwJnGUM7lxCuuPGG5lPLevoX6n+XP6Pp0r9ykK+s
8rN22As+z2xBOV1TYYax/HKMfaySmFlSCBnguc0czqB1SrlzDXrQJcTgpD4U03d1mfVWE1Sgda2E
kgKdorUfg96R0+dUKTl2jVtZojlj7MctlcX1R/SX0k4f9ex/sDnIglOfgffjIFzv52AtWoV+gUr2
1bW1D8oRu2v1GZF0ScCj8O+YUpIg8/lRjK6fB3+lNocmtVyHN4Kg+e7jtniDdud1M0vL0tISJKj8
l3/nMA/d0GGQwm8fN/OG+vKBmKLHCLzdlJnfAxUOHUDgm5O2dBfOE7Go3+Y686JJ0UlZlhohu3IK
92T5CWd5x52Bp4w9AseSAe5Iy3xnGKfPIbcXrroAnf7M9QU2g3r97/B/UgUqKLYGcS8qdZfaWjYg
t2hG9Ua1y9+wyg2g0tTxdJ3G0X6p38oDzOShXFHjKV+EXEGQpb3U314OJ+gT3+8KdY/Ie7SlYa+f
4H3GdmdlXu0wdfKm0l1spb1zI8vWyLG1DReVX4DtjQ1+9aXpyFsubKwqPk99//j/Xfu/vQgSFfIZ
tEdBSusJhH6fNIenUiItT6XcDv1vPAwdmOU9Vp1J1ZYEY0SdmHxg/S2+7jZcUod24AA54EVFAp5H
KPExKp7ti9nGf8wT8KXWh/Fy5HDQYz3M5QGCL2IJCM/5zpnGxYFYsIC+aJ9dYgb4BYv6Z6Ai6o4D
dImHnIcKq2V1NRAzb6L8lOsvQlXYy79B1T0YtlcAtGs6Orxb1Lor4UjLdbyEHA3TyH3kxOM15VCu
TwBo+stL2Z/4qy/OSQto8HQfTh7Q2xnzwXNHO6he+TNEy2Wc6nOQUBCJ+P3mmA8JZyLtpN13osRh
HVNIiYPTzfZ6G7Jv8ZCfYpO5lKbQPeFYohoXgq+lYU8/KN+LUeymCH6LE/ZMqIRoCBKrIj85Kdvx
Tlxbt1crDLfGJpjgBACCb2osSnaZMRlD1Glqp27SzY8rsUvFpab/6DQS3SNc4nd3a4LT9/J14tIE
zWJ3kCgVR6W+1E8gNSkaoxR7JVvBVPPgy+QdY3fYSLvzUTmlhPUypPysLG8uuaoGFKa5iiH8bn0q
rzLmdi0P51zx65vW15Ys7ukvInLT9wSFosSU+JykXKYwO9PvSenlrbpEg4z6dREQhgbCDToxPsya
QNkwwnH/xpjBpWMwA8PMSMiG00si3/B+IOWX13S9ENeYBQglL3AJWIuN05BBetMUM78pSJQznSMs
AsE1Lp+MS71x4VxpjcHLDMUV5aGFZ+QQiG4VA1VHKcqvTs94UStECuUY+na8viFGK+oHUkWF93q6
saSVno7qfBSKRzRlkLfVklRWzqPC5hELfxLKO9ksEZpqcm95h7zek29vib+eten/6dwpRGCf4G3c
+MMXTwv68eIMeEXf6lgkARHKZH/ls0q7t3yEnNQaU6nJw61rHkwYbCZsXDC57zDrUzgVQQINlq6f
CmLOvM1phQY/mAsMqAz7SSNwBTsVp/VZ3AE5yGlMfEquB2kaPIyH1FXHzDx/3xz+hBJrq5+6eqqj
k93thEdKSby8hxSa0AZ02tY1CyP/EpIaKlvKTpemkIMoSLbteKtWOQOlJfqDAvNSoA+n8AJQRIkn
DLYnzB2LASIexCQRF2eHWCZTAMj51zDHHz1GaQ+dnYkAdyJJj9lYmtExrOm5ul7sB5FGhVYG8zqn
4RExv3vokWK5lRQL71UfPCSMcQMy3xvl1dfuYx+6GVr7nj9qo+fKTP5G7C6EWTlM48aXad8Or/aW
yhc1g/+8wEmgIxM6e0tQXRVX4QqBibVGHSdkDGMJHKI1tWvbBUqy+ZZRG8yHflSIfIl+Lvi5EaRM
fMrB44fu0sLVyg95iNfcc5hHjjfmRtwfLpdLgmIBZnSPzl3EVhePBQXNzCwNDEGx6NPwpr8UIiv9
+xy/4LRhqvUgRc6wnCMmH3NQdatoVR9UmqoCXDfa36mIGcIUz7CbE1mVhqzjQgCDpc9It8MXwigj
YvCg+jcLVRffpat/+KpXEzAIV9uXm8uVYQ9YB45iPvNoiBw8fodhSk9RHwKMFigdEgu7q4HRgYvS
pE8rDaNGB2nPMXqWf/xmdEt1G/BujBDt6rBVdzJpsq3P9DfsOEl6/6h+8LX/re+aZVXPNqYM4iUN
IGLFzg7oGbOPKVzkBDd38H3u8i8vM8EB7uSCLwB4JNA/rtqEQ41MiIkYfQToHScxiK2eGelLYLna
tkSUmdTshY00nzIlCNwAW2vtuuICRpw8I8+y4Nu21iMTjPvAD7pK+ukAXf+UUejS/4MIXs2t2WWK
FDsIMinSO3MMUnjp+xLuJrAkzZczVE/DCloqPK2TsNWj3ckhMWfVBr12TBXSqPf+UD+m+nFBXzaN
7JGnvQGzIOaj32L22ELyP4AuOMMD8WfOSzkqgQJIn9PROBLkDrYdlWqDaoGufDbUuxEzbzNdCuY7
CFRPMMR8y2Z8v8DMzC3o9mF7Ee9+P3gZ4B8fHUlsnhr4vEiA0ZsHZPGD4OD5bVUIsxJFAS5yBWJJ
OOPyyIeWFYShxQuwjVCom/UuHDGBHCgSzxPd9LyhXq3ztDk9CPsOVu55eF3yCznpqsY4GDbS/AEI
fq+Jm5EPP0nrJd5vVqpi5nMHXJrrQ0LN1xUM5YwUx6W0oJ7DFAyhcFEMhlDdL+bSYDQA8RPUt5dk
JkMcBtRCpxF5UIbjwEaJWjoiQ/1+IETjDjntUwRixFkF3lyeIgHN4gP7RDdkgsOFHRHjQC+Lr0Lw
VQZ/d563wSXKPyhzJG4Qi7YyvvfIjJr5oF+Q/2Ryl74WU8m5NFgejpt+lPph48i0BfFt7YqUjrfz
jcvpYUrm894MjBajArLmmoXqEYJrch8VbaeZZz4nvkYNOa3ufquOxvSpwZasJq9OJC91m37553ms
5gua5OVFFN7fFOvMLaxsv7AJ6YAHvAWKtc8T+U2qEu/4W6lh4GywPRZMrVxnLt3uY4OzAIDYufjt
nE8vKVAoecJBAO4X23wvduoxH+5a3X+BPX7T/JIA+jlInr55UeYwc8pmHTFn3ApJJlFfLDys9ikp
kgBM5AlpMtgscnPRRFdRw6PfTsGrcRwvaLrAr6h7lFdEwDRnSNSFysuJ3bqyhV6zjaemcRSs8kD8
Zs0r6zxSsLILGWuT1xuVxW5NWtPCg0sdHg4ERnX3hXtBSBMUi/IVMoJubyyXasVnVKXdgfjK434u
bRT9Kh4RVQqNlAXmx0MJabATUvAYpEO6Mdx1nU5LdCP0sw2JmY7xLjuxg3xyKF//WQlBz6YYDm8E
BWAicyQPDv/wRF3XkhSPKD/EzWLmvHdYvoK9tSDYwU5O5StWFBFgfFCwiXRKMEs9SzmcTLZJIMoK
3d0dRm+FGHEqAwENkLs51OrKPhQmdcOigPU9vx7sw3wQLoc/aO/cHvbhOwwAsTfYw/A2W0j2r2rf
r+voKZOmXy2kn+lJ9HtIOlcMNxZc563RFMshjbrJGTN4E2OyZfCkELelsapXXd5lpus1jTPTi+FQ
d4tnQf2eevkWJ3w40w/TNEOuboev5fCn5hAbVK3+BKEZz+F0qAqwL4/NKtRupAKGXJhKDvMjyhzF
EHSDMEPwFUuzkV5yWT+GF6PrcE5mwFRoJnxwOYih4e/CryJMJGa4zKfXl4aPHoyjfivznJhEiV/A
bREGhLaRrH5XoYmrUPjoQ6QOm+SM385dtq0tYUk7xmDRZLdRxQsx9e9anR2Tfv7dl++wjAqz2yMn
xhQQxdEC0aP1WNtIAOR2PVToj/TzG8GQUXWBqDmhR/MwVhjXu1QYc1kzKzgHq+Os9MW8WCIPTFSw
e4D6sN57ziuU8JukFt/BvrQDw+mTO47DwRej82P7ZbUtMXSittwT8S6oFl4xJ/sIW6MWG+Bz0RIf
FAcDNBxHzrov0SxGDHY+KSCkDFNElqsEu+dT026mw3jUwMiC+cNl8ZUNXIZouvWtWlGAHFepGtHZ
LrNg/MosfphA8PFGIGk2Pasl+lQj8b5RTou8BYl5SPPvAGL7g5xp4zPKLoYxvZuHaOStZN0/vFcq
yT5sIfB3hURRwrCjDgMI2ALmPjEGEcoLcVAIN240C2AYIKHd/oN4RsoM+y5BHmHzK8oGW3jdMwnW
vWAOe/bB7NN2XXLFiL/U4N0YLMBAR0zbWSIIkROr4yBl9PUHKQhm0pxzvGlHFDd54dyO5y7qhruz
8ztLjpS/C7r4wHJwk/npHlD14xweBTWAYgtifEXtzSilKHZMu7RIwFwIhYf6Z7aTXBud7DbTuQru
mrPAkHS7J8GJaN4ySCdGN3uPbeeyqyvRXNJPpeWUiv4fct6q6rXI95ftuAX3/MFiQm4qGh11p72E
IpoSPcIxT6gBHfCPqN8e+Fq8fLSZw7v/zy7rVmNsQ2eCbJzFpfnWez8iTqJWJyZw+y3G2UplvOwn
J6N1ajMEfHiLvV8s8OSKVFCmgy82WJbL0TY/kP5SrAYkefW/Dm4Oht0WNspYwHzKHs5V0LmUHYbU
d6dv72So8UCeRBjP1A8pl3KNHlKvaw8idWhYSCuj0dsXCl7Q72avxLacENs99ysYk64aoJ9YH0cL
pYyjgMEjPbuZIK7t30A3qCx3Bx2WqdpsWNznBvEght/6Y+tonQbbZG6hH82xmz+5ZdDX/FI7AOig
IE6SNFbRpfZKh71w21xA2pzAUTMcR0JaC8y6MbU6hqlhh2I8xKSWM/x+yjlcxc7NQreqIGs6iBC6
gzdU6jlvxYl43BJGtlv4Pc39EpSgiRY1sXLPAit8b5KlUb7/EsTG+snMaEjTt5l0m6bmm5ice/n8
jEYM2gaKdUW+lm0dGWXlq8+TRuhLIVR00vCvrDE2kw8FE1wqEV7KvORUKYkooFFf0cU5MMuIKlSk
W7MOinp6p5Gd3e+BEGzzMMNUjzzxhta0esbLQOfxKljKaYmI5M7/qqRmMyBV8H8pcRDH9KKKjTmp
6ayOXwNoZQU9iV5Jb2Ps9vfE4Iv+q1ldZOCwRE3M1IFm2y39aAXt/j22R7IvjdFRImBxQTWtpHhN
4M36HKHEoXkIAxEJnuKSAvRmQX2WtpoXG9WJ6S+lvgbSy4HQwD7my2EzSXFpqOxeO7eO4/p2TH1G
POL0aVdOAXpe7njfTb8yjIJytRm0VIwAgYigZBqWtMTsYgapN3ioZ+L4/FNxV7gjoJbL+c88mIg1
mtjWZk2HssO/YvVlAykUPQfjYLNOZsN5WJjZDWKL9i+vUHmcWTYhnKqvcy1YMqUN10JiDeaNkiBt
7/0Jj6vyL93azVi9ywm3shbz5daAorX+fg+U8DSWU/JPeWBDVIm5rKss4y+KG9B/Hadnt5cKgd0L
bBjBR9FBR65IGoZUVD+0OSnQ5p0bblhbbwk7r9hH0on7jyQP15L8Cz1/Tv/QWWsUTsQ1pF4kJJNs
x0Kmzdp/0DTxadICxKFuINGg8PDeX4fC35p7yZ4e4zt9F4eMlx0OWDLvhZkqRyWMvVazfX9w1lSz
yYPceQjxXA4KbD2ie8xtVidfv2ZabBLY3b3POKgGOVGdBvviMVAluXf/gTHOzWvMECKrNFuOFzZF
12x+CrpHC2uxPoHv+8qvMrusV5zGN43YOXRzW87aPq+mG0D+hKBPFLEKY5CFS2w0owQ1+H4+tu3R
yduflUY09N6xiTnr/V2J4uFPH+RlbB0gX8KfXcudRQSTsCGFgDry62ApyQu26fKA6kFNgZT82+KL
w2Dy5xtqrYHAYPZSz4kK5XW7id4RywoPbnAHNM4r/NJaQX2c/twzGfcWH6AWrTmUmP7TPkK2Lz/I
ppJAaCJ4l+VbkGYbIqsYPe8wD+HP+ZwDHiM3SQKl2RzXO/8ITwXuOAQ+mhLO87R2Rtn4duP2fBOd
iL20pOlFQ0ilRuJDXXROaYwt5daLGDe+P/L3KRiGQVTBEhOf/espHpF/Cs0H/KAk1/FhdOcEj/bQ
A3wOeKZPP5IF6ptQ3ytBv3hBajwCy3mrjyVMxlD7BzubQry36FRn56wAD88ZSZo7VdGsG8ib6lLy
4VyJEpOnJcZlMNRA9/qTEme+OBqmRBRCAKDCDEweCByKwmBnsk6XK/JapYxbG5xvCdNWhJo9JT13
NB/DGHxiyNZzY5TS0ErZWAYzirIg2YatpmHdE1sny/fX39c56JVCvpZbt3FIexv6o9hJv1oujQQl
vk23alLjVIBBsqHOSBy3NAUA0nPpzgWm/GngOjTfx7CvMuCtO8m2lYYc2s3p2nmmlpjH7zsJ5zRj
N2WeRKqbMrFnzqncr3XLMe/xzP4Jhe3Bk0fgS+UI+w3q8cdu9aIVOtAKLHOnkr36Rvd1dfJW24Wm
Izchz0usmJCeNCHrNbuhUz+/i4V+j+eM4PciAjcSPsEygyLsMa9pl5pECWcauo1V9yQTooSlVo8H
VfAtYOmEUuyostDUsBJ7vOV+BE7Finzd0Xw5P6yLTo0zjaj40NhT6darCVt+lLF3ODCATwpiqpbA
nexCaXxnkN0VtUjZuQUFmFrVMELcVJorIiQC4825Y5XcDteKq3ZrYea5JW1dEPTer4f4C3sDassy
Gd+bhXu1nQlSIeFtfXY0xiSpZXLuIkRYmG5yt3l1Z8UtcpKqRTPGgnBeeRLw+kTQ9B0Ewd33x4J9
zxemquBtkugfN3B5atF+p5s7/ThVvbXqIxz01ELFtxeCpMy5cnC6TnqmlaUrHCb7NX/htdeC5pDN
R8DLGijdP2ET+2xmkm0DNeBl6KB+Xc8FMBKRKSbliVrzflMSrs/jK0G6Jl9IYmQR98eqieqzWKmv
oudqmxDL7HZzBaNPxrIK/bGsjSwlLHdtQKjfi9opOco0X5TV2HHH1LvrWvK6DuNaqqJ+QzS+D5Tg
eUul+HFq2OfyUVgzp+eTPapJAhO6AW6tfy51alr6FJ10aDsE952qcs/vJqgJhR/G/9SAKLH/gnca
oEk1poeTZV2SAdpGN71ujTzet18QdHmUz0Uen/+68xPO2GUtow05MpZ9OBdDxlL4cBtKJHjM0vr1
tczqLx4JPlwM5ZJqzzmikAY7u8n7K3q8MUJl1e/q+pkVcdiRRq7FHBvBkl/3+JizEddqVi9cCx35
fQVzr96qgNMGbTqCi/oPx2KJYVbKunZeJKyuWdLIJvd0vl53FhhSKaqyTubmn30wv23zBe8njBLM
GM1A+9ZU8upA2v0ki6mFx/DNQFyLvBBQl2CRpM4VzgcQKaafLhVA01XxUDIPacAxzneBmmZSa0/J
Y8wP/siuOk0TqHv86+0V9bN2mYPqnuedzB1I0KiXYsIJDj6igumIS730oZA8U+u/4hSVtmmXOtNR
aCzvB+JKZi8o0KMj3xc7D8XjkRCo0iyY7DtBFbJaKQCVIgNyO57Iqqv6oZmQuaANs2Xn9IK9KtXN
y1WcoC4DHSv+cqHfRPULcrPxA3BYUDDhb1g6HqUkYKGPabtn++55hG3DV+UiF5oUfhCnU53iRgoo
B52RqQ0DjJGGAN84ujEefyAkTng703MaFywpWJ72WySSfcgrs2Aki7CtZatdqq7hV5mLb4gOnNJt
BV1r2byucjPk4uLCKkArMyB3D88WkJs1GT+yQLMWoigK5iWvogno6HlfLYjRx2/jHgXUpeXaFrtT
caGAmSnACrIORntDjYCerZNkW0brIKNfDU+BIfFG6nbWFPJSOSS91Me/vgJM+REZDLlsono3hC/0
16FT2ghxOQxdwT9FBKivvaNcqLXWvSRLxOc3ONE2Uiw1DvLY7PhtT7WzXatqKXHRzfYvg9C812pl
N87l1ZOkmLNKSH58l2BTic0b/TJjeigebCcbKtN53gxh6B6J76KwW6adWJJupaoez+8Vb4zHZu8W
Gft3EJOV4bjwZAdxVKKexpZkx04AMfDlA+rJpx1k/vd9h96Y/pVtdRcVVFCB5RFs5l3P8rBEyVYj
zxeVzHaDfd7MFpRKFkG66XIDnWvMpKCOr3T6OffT9aVE07uCExFjYS/t3Kf0MFFOwTC5x++E1Qx+
Zd63XWrHfr5ZQPtC/Vk0oqjMXekgr69K2Gkkp9Yv8da33+S5noJ7rv8A5k+awB+bdJBq/mPX0BDF
/XDgBHNmS48ItAGOjYKu+GfXfLYwaj9zqf3p0hb6BJhjZUcu3FMtJz5KCa9hxs7SRZNaYghE5g39
Cwp0xMrhFC2OXOKKIDaBQ4UxtrZ+7t1OhZkIwRE7e+giHH8fdDrfW6NpVRqjagFf4eHK5stuIniA
fbDB0XmLjux5tDbz1H5MleCI4KOJ6mDv/e1H36iYflhVna/gG17QtLINUV4qNgpyS+OrBbZjnvhl
uqI5Rfz2XAjN4HsWQ5KIOOkWdnltd3n/RQc0cKw/AEuaIE/I6+PbuB3eJXopENGH1MLmGU7FbP5s
RTPAQmU3hku36YIlxMZNL5N11dM6gg7uI9Le8sCnb0Y9EkyrzjWjiMpJhGTR4aJzv1FiL2Xtd1b/
PLiC2sBFRM3cKR6OSFo5gdMBfJBuDtz62OTlfDDeeo+vk9J6ekVL8z3kxUkS47/wDk7rtvHVThZJ
oXjmi9X0abUF1bhljayG5zNmHg4VLTCUi1SK4iK3P+oIlLEXbDIrbyCcuGBlqp8hTD9RSM2VQpM5
ZjduTHcBsIHdbLfDiF/A5sgTDig0q2woJc73VBGKD7b4zYZ//6xSiti7RoByP4hPhl8Y3v3OpRyO
+3w3YXMEQCuElxnOCh+A+iFyvkxtzO/xcPw10Yi/AmlUpxo6JWCGc3xIHeoqqL4m/FIPBK9H/rwO
ZEfY8i7HwuNRaHpeCtBWjetAvU+7weKlA/qQZgq7V9EV7KPpVZ/PQqlW/TPRwVWVK7l88qYtaSq9
nHzi1QWOZ4dffFWykN3uT4+83kqYoFGvsXk/gaAXO+GzruK3x7GEOAsjoMDF62ECr9qMyfQrTQoQ
OozKUeJAXnkn9nVCmJSj5cy3pc59EjZuckoVMjszH0mtjRxKNpTDdq5Rm7p+Ii6O4ow7Ba51bVEU
3KscFYmSMUao2aMeqPT5CNUuSiYSWqmND/TKH4T+MjzzrYQAHHF5iHjn1xLjQXvMXHMMqUT2eHrX
EkvuYC1cEEQaAXLiSJi3KLk5Xje0voWM4j1RBKFfoRlRy3HQ2IM5DxouW1ZKkoHQCTILwCiztKJf
yItawJ7Y8mZMBSWU6gKBXdwRAp4UC891GP0/9B8K16PnV9ejEasoGc2Z8HW4YRe6ammwnatPC0zW
WHBokMQnG0SvTzbP+JBmWoc6hU8IpmuOC+BzO1aeQ8OaV0Ui66D72AV861OSqPJ2DIeusy4vg6m5
X33QZLQxQDbZrs/tcoN3mZkLJGIz/y9/OkSoXKnlYZLcmEfM7BCgTLreFjlsry6kLzATWoL6jNf6
PBIOk6zZsOY4E2KNyuM3BYCOaubbG981Q2RPQlxQZWjyYpkpNnInmzxJS2iLPXHKKUCFxOFSdx9E
m7+ldH2jZeXok5jBo3E1e0ldrk0uwj3CLMuGMZFrOWiDTculuZ0eTKwmd9QM2jVXK7pyReLOHiTR
GwlR91olCwqu5BLIjiz+a6/n9yDlIsJn4NV6dKOolqhp8n7uBsw+ovwJj7H4xmACJdVuZF3T+x21
/Bq+NAHBzj554gpzpwb6Ehl85LcAOHu1mjvNlZ8z1KoOMT2bYAAlEDCVG2AMjxvLVvWyn23NbDfA
lHnr886Uuh/mSgTP3L4RB67LlOs734dTNadnf4FQhPTPjw4QllP0yd8vu7rZgmmvzpWTVMSb+q5A
bdDNWBYTY2XOZFX82CXEY9EP1dfUJ/oHRPn7SlvUP8IQYixT32pJEjXQmxlU5LLj/GCX71DXaPJH
gP9HaTktUXBKXnLm+vlKoJffxWK7QZqNK81QY+WO4ABPCxQoEIF9X4+tKD8O+IGeCOSciINlfWay
hDbzJ6QA+JklTc9odwQ5NitbrgjGOzjxIW8cIhYdplxF1l5ChuEQdE53nZvNWNpSaZUXAShC8fWO
4ESsKHQBQtijT7GWMEHo8V3A15fLdbLSgQGGbBK6HNFjRVte2knQT+f+7JZ9PZnmY7YXVkM0QiL9
1652TvBvBZqc9F3S5H1JtMOgNdo6veh11nWV0cpJ2PbuON83G6vYI+UAUUaV78/Y5pelc1TTuIbk
77hk5HF2WOJehtv2XS1wea6sd+WRXDdT5srxrCb4foBo1Tq5IdiWSTw5jG/wckwueqwQe3/vkEZ7
VZd2KBfsBj3bZcofrGA51rRXB7pEuqXrl6gyFszmL90f1UP4rFwj25Cye60H0lbhcgM9NalINicc
5a/74SImwCaduDi627hxoIxj9e8C2jI1gdBzw3kb7D/fZ7liBtpX4UQSZD06uPQCW7nX0PDC7o8/
pYNqRDpTRP9ZW4CRyMv0fv0ct+QiOL1PeitSRjGNzOpOE/3mJjmq3hun2TeK+9pASZDL/8HJgDrp
rFV/lsHU7wl1YfKgq85PT2/QVYFVhn1GLok74FG7FaZ+toMkAeKMZiwHPxePm/qVjipfQt8pagp6
OIEz7R6Toex///FhmaleYcjoBqIqnh1hPocmUURZn6Ds2zgxzcnRmfZZnGYRflcccOhAvzRw2c0m
zreMbw+aRYOa89ydDJ15OwS4Ycign7DNiDxQZe1/UXLBtTIbvOPp3bUh/vIeM84I0BMG6WXkNhjc
+HUjZuPsfQgB/4Wu7WsDp61CzYTQtXyA2suerewzZ0clk0MT5KZAR/El++v+58H1RMQQ8BjQ4xZy
VYagp7/0VFf113e1OiqQVk+taiFUfs3WHx/PmR3dSadj1N4xmmo437joVVfG3GEkpO0ChB9ITpTH
W/HYDpiIWMowQD41dsixovdXZu7wsNivdTTHW6d5k4Rq9IGW43KnHWeO2qswoXKcc15Dummd6qch
9sAwhS3W+1JNGJj3nQcpB4pTzqZSzBXlYIobUg+yxV32JPsozIeUgtbKMKgeNNfZmxZvqNPmSnAK
KSo2FIPy1nx5FElvGvaryLsygiWVIYzshuJuDQSak/wkA7hNIl3QIqTqMkoitPNp0uw7eqZDxk+p
DACrBsmL3eOFL5oKuOIH8SKkdZ2q24X6a4J9AjwR1m3aQFi3n67zDw3bwYypVbCheLGsKnZZfpFe
EfsXT7iPsxPwB2U3W6PE8qxdMb87ypAfb0cksRpl8K64iVmMtmDu/abb1mH3tZ7rZwNKcMvag8Bb
oBfjLo50ZyA9iJ1w+qz2qprhMDlqXip2mUqrMGs9OZJBZPSFJ6ijYfzAabUTgviAZeMebPBXBErV
8ao4WJuXAp8xCGVY3A6yHWXGlurt+ixoDK5H5yx2W2QWKyqk6Z/GZVh7iVJJLzT2f2pZd8Zwwxh8
ZIzuLjl5ZzMstg1j+izMLkEwffApNqEwlEXqSS4JZE+I6G+wREe8CwcmbiBwcPXb7L5WF5lSMKjv
mD6Ow4+UGptK9GL7QmjyQ79j7uR3d8GB9uuag3KOK+Pux1VmaQ3jFyOVHYDOhkUde+Fd233SaTBW
8W3DvTqQen6fDeimvPEiS1n/hAM7fqVdvOoRNUHdAxDo6MKNJI5foK+Q7KtKK6y925kxrADwC5BM
2B6vZIAtvrN+oS6Yx/k7ao9Z5ax6wZXmJSHNquTDD4FNUdZNsWTy6ptPLWJCYDb/yQw8+Gso5O7e
5VzuDQHKtMfqe0RHtErhtIX0g5GpqhIEYY4x0v788HTOuWcxtz7coZr0kg/elF7V1z5RzgKSQdUm
L46R/ZUV/jwN1fYFGZrPs7UqiYRe7JwN3Eonlls8npG33DdFKoJETmjsua9QbSlwSztc6HDIdks8
Jc2PwtgBim0Ufj53OYeOMqWSkzlqlKg/7z0sfua1/kdo8KSTu9RJHW4FUNXY30sefhK3CbXSiee5
QJmiz88oyISeCjBB3JuN+jPY+OPnMtYW+1IzHzVT5ont1fI0/lJJFsTY/YZx6SNxRG8HM+h39dpx
+HjNxoccCOOhqd88rIhIDjrZw0KsjlAgcVpxwoY54WDdrS56RKP/XidxLo429W0+CkEismb/aiTM
vPR+CBEiX0ygdjQoyN98nhEa4kK0FVUUbdT415xMGX6CDxTVM0ztdcLz7xVdF/naFqudo5rn+T7j
utTePPd3VYUujy0lmMh1PAy7ac/Yh+2WQbpWHqC1jWR2rlV6YYnF1mnL3GFuiQhKm6OBAW+XuDII
C6q92YZJefSYBlJQHVNoQMK8kCEQ3O7uSKP2pb1smXXD7VYaMAzo6ugDLxf+pzxmxQZMNky4hokU
tGR+YxVVM8YmnRs0Dt+4AQMcxpEzXgnujczOhZCEMjdWn6dTku/tgCUJBUIFhZmmAnZ/fhfznrjg
IyU2D5h7poHuItmSLxk3PGLCQAjbYVLJvCuNS7NoeUGHgYUeQZ+7Bz1lzZ+w/+s8fhaYOJjSpjk9
G4fTEidbfueMxoKwi8ZwyWOf2ZtSNzWMs6IehSleAwyFWGYBDPzdOhGQRP4kpJzXaceKHj0VGQPu
J4k+fyp5D7AXLkn9Ip/zufJlO/p4pG5h/kSlHAOrO7DIlXTtUh7RSzHJhZ4isPNS89fUf/Mtj6LF
FnR2o+9KfF8oVcLcQoJTP+OemMu2tOAMa5SDpQNNg4Ss/l1MEK68IaJM/gwav9vxmZUXzcWDx/WP
FO8bXyAiW7x50AZEuAJHKv2rJYxGt+E7Yn6eOlWMFzKusAByE+GPJfyG+AgtmqY+gnfqIEDepkKd
DEXrMWYTdUEoqXPH2cXag8JL4wiVlzvKDbnDFAO8nBy1NfpSNishP++t+7UBOEU/xCKdjQ93xefE
W1JYga1itq08fSk3hZ/gjxgn5Ah8VPIT0YPfD9hfQ47Gh3zZviIJ+BSC4apRUwyMTXQdy6aIt07/
zCCe16CidOh/KS/W9V8vdPdFLUTHFBhVEXHIKjtEjw6551LfRINYuX0NNMS/vEIWTFk7LpcnQMfP
Iav4kA40UE+zrtpwei4V+FzFkVmHma2z+tXba+7ZmAJblNwW52xzAsxQRU82VPu9NwLtm4ht1v/Z
kIe5Bn26fP15DX0Q6JYLTksfdSTUOoA0eyj/aHdSaInnyChovF5jCBEQrOX6+L+MQlBGfjVUufer
B0DXg8VHisjnKEWs+ZwqCu/FjdfvGF8A8zcOFP5G6fbemDJUaZ9/xLXi1aHSOlJrTDhqYs2mQ6Tq
I/ZspyPs0vmh3eD0FkLO7/f4EEPzidDbB/xDt7+W9wQWoXyKIerC3BKYXUmOZ4osiL27hxYLJbpJ
worS4r9tqlas2En0/xL6DVHcKZC8hhmmnCI8T8my2T8odGewRMcEN+aNaqeuoZgjZTHDdqoSsygM
AfEMUmpregl9shDVx+1Q2w6Qn8K43szzrVyzyXUQOwNqPHbYI9US/RlzktwVh2gj+RsCsMGfdxnL
LRdYfjClLOmmgTey2GVKw7VH/k1h6Z1y7iMygUQJR8y35L8rZ8vYuibTOgokAwPpTuDQUFIfCZg5
fRSHZjH69UCQr6/TVuJCdypz4F6fhL6pWP18xWN1rq4OS7dLuGD/A1klFlK772/aDq2D5vtbERbF
1lnT3Cd7MclscPyH8pl26DgFJAql3Yeknu16kyYH4wNbx0fMNf1BIKZuAgHpAZyQnODl+li3C6Ku
E9cub5KKO+7YHCYIFX3rhZ4PYu+nJwsbSARRbT05pDEU2PRKI1XCbl7CSvAnmzZHlQ9RgQoR+01I
oy82ozXlRgp9xu7K1Ow+1sIxs6x1h5DIU9ZJG7RrI3ocGjxr6Y2tZS2rMGJauEYtYuuAtFGonZDB
qh1uoQbG0axR3igvMIfAax7tJ8MjwdjAMrBrtyM++OMARYuzUm1CnTqKGnRrFcb304APof3sa0DA
64/f4l/2ko4C3D49aH+pIbKZKzZuo3bFTbWSKQr7xkzveILHztsVOPgLh6sJcL66SNrMrJKOkVOQ
+71d7O+aUIZK1nTw4ErBL3njqwKmpAkYCTJS04Cb3OiP6p1SLuDjptgG+3xQLJF1wniq1zBH3isa
jklODyXMqPMAJmS7+hlud3IEFxaEswRvZRmC17HgpUIm82P7GBOkN2DVRBwB7v8/fUGa1mEtnsUG
2uxqBAtRY6h/G8AVo+qxYEXIqI/u3GgxgLVnjX/ydUNXlLxdoB1aRXvDx5dCzUL/flDSo9dx9KP3
MFiIOnruYlEeVpcyjOHAUoQGOnK5+VLSS/bcffa7g2jXhQ2Q0hTKvlx+wwoFn6HsUlIISVhe0A4s
Pf2jloeyQzt6I0GXQo3OMtUg3DAalE/ZrgNjEYhPym3+aC33f9ajX30tZJP4hPoMxz3Z3PXAOUPI
T4PsTq7gjEx/YRJSZ1vOTN9X+IyjvE1I/nAPrAAb+rbLEMrPSRxQUPKlWPJCBNZ/OI4gIIMOvVlQ
6lq9eiiUg66roM/ec+OcVtLdSx60lPFZkQx6uImYefRWy/XqpgCe+KiEaex+/xH9LNckX2w+Q9nF
t1sK8TYIZn3TGFfz2ZLZQuT5D3LGwcBYnzgv97+JgxtOXjo7N23ePXzgQ/udNG7eBG+lPLh7nJc0
o87JXuMlmArLESzyPjvT/eLJbhAtuB+bbjhHSPRT2wkDrNKdq17A0LXfbcoxvDk3dF6NADZR0HUf
qpjcITLWNxZ9voduJFuI//XqTb0YcnE12M/qrdBUtCE37+ZF+HlE+bMLDJUzycN+xWdZFpG+LYvB
8eI1tEBAgFLrbYinWqZfwLFLPRU/EymjvWaUGKW4y72S3cZNa2Xpzj1FZeT24+TcewME5m4V23+B
4K1ZF2xHlMVSGS8a5Xn/g0qDrAcRpc3bRnjJvVMFgv3V4ZpmmEOIxH9kzrbsrp7FHm6pK4MyzGcT
lfscuvmybvh1jdmEmP5YPkZb1TBqd1B5725RyAyteKeKwugpwwS1ufhAt8KZLwrbzIvlxvf2GJEq
TAV+IofwTYsnK0AbWYCTcVMv28sAPsDoSZvX5mfjn6cWjaZhZovpRbNs8eSzGXGBErlD+mYF1oqa
zV9WrTYbDcW/NvmEfnNPMKUUYpo7KFYCw/Rb6zoPmjOUMeQBKa6g9UMC9cIjTTy+7Wv8HKkJZSpN
1HWfGWE4meg+oMzHDkFDerTQZlusP2tjxtfUoN3Ga6FpQrKtiazFJrWmTwdTO4LNztIKjG9hEN8D
5VPIglGJ41202z8NCwjCKspH5W50BKQLHoUAf7fGrxv0Q6Yr+RzJhilS5bX6MTYy3zL5dYlKZ9+z
YnKbRtB/uB3HsFHU44NOVbLMzrNGWKt22vBx3UEaiTQkAl+XkEvEWKJ1GGo6JofjVHzbRRZHGZNd
qD+b2JStDfvAT4FsvRp+1x5Mk3VnrKQgbmo+V4GwLfYf984MSCxlKMfpEF4fad+7VXTP0GyIepYD
k+rxI4SzvFIILxvgFFVGAbZRSnaZsG2ba4xzXeAJ79uPFE0ZQ3HtNAXQiS4goge9IR8Qt0or23cU
TMiABtvZ/f473VnjNnsBdYaUGpYraOSH3jBJ/gmU/Z6AJh0RxS6fKVUqOR8L325ih+SOxjRTOX7L
As4f7vuaxRf6HTyKhhSATzWyAXw+f4Bh0w/BiFcJO2nwjmGQWF88Olhnf5RIRAfVdXr/YgAsrmU9
8dRnzTeCCRzPuSVFoHG6Z3YSz7FUlrez5C5Hz0vD9rqA2k1WQfXZoOUXJ8eUt9Kj/hYwc+cnlOrr
8Q/L3ywvw/BnqxyVzyDAGGhljXHE/vtZ3cajAfLCNk3QaK3pIEYRFtVQSejV+jaM11C7ZDNPLssf
Z/tqXzB76zEiA/nNsJkt3X6pk7esh806vfpIukB81+w4JB3A0I74L4Gc7k2p0lIU5qif4ex5dR1G
Q3AT+/A0GidLITMKJeoPnKW5NDOc6j1ulD9TebS+NLIbZDGDwNDeTVm4kX6LgAjXRYpzkeiswDk3
ICOjmEvPk55L1Ni9iVin0kHbVbkqVL0LBLmfZRPooC7tE7denAo/Zm0MXG4E/3uMhoZEqNO8GVR2
FKsIM275qE1F8QOoLDnVrmJpGlqF0qJ5UTE6aqKfDhgPi43Tfs50jQ5xNjO0WyJ3auxyF9tkaH07
zFU7TDsy7RG4ocDhmync7ZQCWw/+apL2DqA2eGdzt5TbhJFH0EvDwFCchZPWrQtXC98g2LUK6z9f
QjwRF6tSuWom+p91Gtp638c4+t5MInn9weYuLFol8Xjclqp5I5ATopfBMikiQ+qMwbO5qXVuTNPd
NHvf8HsEM9ycw8gmMXiY3Dq4jQJM5oVH+Zt0mZRNMwc3pZTWTyoXt24cmzKFtv+SfXSlCfQ3caS6
u43KhMxCScWBJqqB+apv00nYj79X0qLuSW0t6IFBnrRcpWqhSvYKMbrSxCo864PmtIPrXRQbgQao
9QmE8F9WyHCMTsPBWp1r2LwNDtDMGX4GpeK5EdkMq8zWVFoF6XworPA0tQMzYm5V53lC83cxc7rS
yVhBUlj1SFtlWyyG1SUqaeJ8fZiX7EDaicBhXWHlbX7qpx8AWWAyWqkc4syQvCq0yka7y9RE2+cS
LkG199G3GieR/BK0yu+YGRUBwBntuK0R6WLRmXTSF7EeOGsuWj1EUGW//k6DhEn94sOeoMilrAOc
shbMJh0cGuhLq4o7LrU6MvnEF7lQtClZzw18Pd3pOn4ioo1syZ2PC7SID1TJ5ejL5/SxDOqOblt5
2sV3mVleg4SxIDykffCppFUVhVYmLRTUsxlALfn0pLI4ungogFINN0ne0UhVwUuTTDCWI5mNboM2
YLyZAYReEkPNN1g7H/Gm5Uy9Efd5yLZ2XJtqLLsTspUECn8+eFI3h1OfK8YXKuPJBwp1lJhz60uY
iEzAqE6TxohSBx01k/26Sozds4+nm9Skl798E1sH3ITv/Xs+rRKJNFy5HGA1hQyJXBhOv66zhnY4
8rVHgOOY0nIrScVi7Rv0bDdH3iMaGZwvvqDVyb9U8MqfthPzIZL8Y9o2JlLDNAErW2Ev6mdV64J6
1zwgrMs+9lrzMAuyed/C86K9J0YlzWbyzpS8DAI2MYK2oO1JTrMGzoVxKBHEy0vUcKLUffxZWDKg
klZaUk8F405n1Vfcv9sia0SaZae7LO7PYTptczaUkAyrtJxocV/DFC+FP+h27NCmdm+jw3B1/n+K
EuFqb5feBgYdFoJV60wgjEitcdCIzbcrX7UUhSvPPiOG1xZHGfmJyhs5t29TXrV+jn+i6fB5SgSe
eD29tTLcyAOGob8dy2uPeKF8gPp2uvQvPN0N6X5t1NurmQ3tPZu5kTEzoxyXEpTnbEbwqffRMW2R
l4vyGv0XmvkVCEsO/nAEgT+RonfukuQsjK8m2oyQ8rdtisX/qYlJRYP+J4zcmapLHNXBXX6Jqnpj
wshqsbTKKv/NyCp1Jtwr6QtJBkCkP1duGBkDPktdy9PMNFkU/liZ3dtn3w1HPVQbQcf46iYmPvQz
T7ukM3LTclCguu3XmZCD2WSjLYqEFrwCBGeg5E9eWRqKNAKLTUTMPOARhMAKMwk+WQ1zHl9tD+pI
pqxAH1Qcmja/LtQrJMTSklokKikRLyxoHxilY4EOqlaBiLb1bpjLZjGIRQO6b0aDFs6YG1tlQjgg
M4jkpj9gTgBNBzBIWBJa1WFELZXqzVwZQ5ZnOAALXbxuD3NpepqkCPQqtCpDwZJx7HETYfQkbIFN
6VP8PpWS3KknWbJJ5tvM3fMmKvKMCUceOlpCQdlaemmFGfnBt99RGrZ89v1qVwHDV+h2fxH5aaQE
mJul82GMqDIH3Qx29OIbRiJMDCvk/pqsbEeSc3IlGCzbHu/B4flXcxvT+YfXliJG3QPaY+OU/jDp
PpXvWuDMgVzNfLoT6oyHtm58xu1Dvb41rztsRoDb4oK4WsyafxF2Acv+tGLBxC4+RKWj3eHmHVNx
Xw6dAen3M7lbBrVPtG3bNU+S9o8CCO4EDn4UzDpSC9JDveBt4JarpyMITVW9Q6TK/ZpTkdv9kbO9
XAYRJVAi2BgY6Okg2rLvVw9DQ+KmE3HxFr3AXKOMjaw9iJoPJMNj4FpfoHzRtcJF4L1TYxPGBR1g
d0Ivg/G7m2RGxtdf2NUtWxRlPEuezvWT40IdVgAHQNYzi1535dE2AVSAbE2mSUn8FXhL8CidDbXz
on7NUC0YVaMPd/HXDiThJUyIiF+a/Lp6b+wca6et+onpdL6U2NqXP65EnORDQ4IMmsEl4RmiCZqD
ADo9ZyVRMuQUR+KchLGx3qiJDEtm2tgmYQ5QUASyCgSjMu79FXZTdyGMDmkYo73+PKS9JPcFUn6Y
qqLlt8it/KKkW3VWMYDc/ECZQzSWyPxdumXo+E3xvZ9urP9etmTJxnW+dh0f9esvfv+nHmpOhQSO
eKzDssjeDJl8d6UjjpuP+PZ27fbJkYiEnpLTo8iONAYL0PSoqtRR2NUSjSeJLYOtSn/9mkxO4a73
s/5le4xhJr7tWiInjvF38NP6kdm34G7Fl1wa0KrvshO8sS8G3uIjAjR51xXHrb1gVS5TmD3AFkrb
KeHltQpPx7KbG4T/ev1L5Ei86iN4vAxd2Fgce3gkSgqjBlH8O3BWVQ8VYXIBqeFqgH75LhZjcd+e
D3d2+E9bXWpDMLmwrzzJs19z4+cFk5SrbUYi0C/lDrt93CdhF2GVLKjyJ+Y7UL/2nUBk10SMePkB
Xh83TU/3cnLRV6Qx7dLlkJ0Z+UYvkHxG2X9wXXwH08dHrJkyOWpXFgOR/B4bzE+zNXSushuA3dxa
1P+KE2WtpfqmUiQoK2JoTLzbNgS2MgwoNqxb9XwZLOEnxBiUsZa0X5O8eAXVJWMuFKSEEvY2iFWe
2G/FVtstRNmSVZaGgx1uvviwQky87kWJrKZo+KtxG6JtZ67GpTWOvjS5oIV2eS0P9jlIkziqFvRp
MWPStafN8OeyJKO8k8C7BpY9uxcezwkpdvF7rAk4TUvaMDcGwPdFUKgv5oPfDnSVPK0v0RYpxFii
bLa4lu2k16bcMv8931VuFfzrmFPQC5YlS0uGB6bPqacB0O9bXdQNaj2L6JzxlH8Chx/I8q3znRYO
CtF6dVhiktO8M5alIFUtsKO2eA+LTwKVNF+jZRtkJBMDATogdwFuhQefKEpLm1poAv41AoBA6G2C
I4A/9EvUz67YSd3RRcl0/vuArvkC0sw7XrmFEK4XXjz11tRPH3/6eebfDpwkqCxFFCaYCigoVl0v
Tfgdvne+GpEDyHyqcixh4DkznibZi/j6l2B+YTROxtueknVeD3C8Qt23t0dnsU/GG+MH6cKtKOe8
VDUhglCee+uVlDyCjrJOJg875EbfcPajQ7z/oRvpCW/ccs451L9wtumkmYC1apwR3qF/KlDJwwws
we3EUFANYsTSZBx64ur9REF1md1ez/EoT+jEVOM226Sw4QZ+j1/+ofxJiU7pRCa/ybDSrXKfLYot
mUkvqiDxMHJlIKnpPvrZ1wqXgKPNKVHo4c75zR0oRkHJA6Wf0heKniZ0eUNtkmuT91pBzp63NDok
HO/nFfLGA8hu6+aL8hl2GYfMS+iDZH3KFc6r3hj+iPEeVm8iBLazGV9xfMeR0uKBAV7U1JnC4Ieu
5qf4OuebytyNr15KpYL/sRWHibSXxedDKjPCxmvFdnUWGv07SpJ25BMl63hLihMOe9AK7qJac3oW
wvq+4T4WA7AtQyE3IWGOADTcjWHuUQHLLmAqSBtSV/EzvGdRBRBb0VkHO9MIsUK/SnZ1TAeRG5PA
7gDTbGzEGI+/PcKfIa38b4DJ6JnAZo2HMv5M6UeYfUkKY8miKA+meH/zLXhpz+ekVdonznQ7TG3g
t8B1/pic+WxJB2xeaptafs3GHWTWZPy4tLtpzGcJ0ig4y/J2tUds+ktdKpucpEpyOUyiXz8GWw7X
g2SD/Zmi5yltV/R2KyWmHqzqaqLeguzdlQAsuFSzo0tYJPkpsaJavQVwStrqDzIVNaiouKzpcZxk
JRFw6lUY3rGHN6iOKScfcPbq2vrcetkySTqrmvYeqNhSMHuGz+ksyu4OZpHkWUnW5jHcbanqqS4F
jq01+j15bqhH4W/KdgVMJx77NJYNmR/+fdzualN5/LKApJCI4Usqaitw2O/klfg8DM3+EH4kPCQP
OkkMxT0BruiBtVqbceCdcgtAuaI/iJ2E3lQx21Nh4KT2iH6lm9HNdkfWWO6uZTweuEv4B/y766Hk
472WGW1baG0XU6/yoxPyzdohkumYQmxhBsc1H6aFqGO2KvpztSUpOeB08qCFgRNHtHrqxwGe64bE
shMeqpvOq5t1JOi85NiYfkgs4y64nrstduj/ab1ajWHRsSBlMUOZfSSfnZhm/GW+nxS1b0Ss0E3n
v4fW5czZ1AXZ+LkBRQ1waIYagYpRmQ4AJKQfRzOsqbSg7mpwOqY0FwwBhrSlgaespR/unK9ZCpIe
QRDEo6TOO1eOxcQNSu7vN3W1+P2xGde3c0G5swHM0/Kr0IYtFKuNB3ZRcxP+6VCnqG2TmrMb90Xp
JdyKUOLVG781PfnbMXn9N3sP4K7uDWuvxynFa1dqrx7zt8RL9yfqRHspvuNySrtBMzpxGmQ06wJT
OwvePVW0FdO94InWSxU7ciu9O7FgyV5HrnfkG0XvsV01mSSkd4QHuwnpT1REbKTcJmjeyawGft3G
F+hoGMXegKKXnzPBNn8RyyTpwOCIgGlGIaMinv6zYs0cwrWA5vJwat+KKmnR7pie2Vj2CexQm7OE
YDCl9jG7CLDjjMXUU56mzaFuMcM9/r9vqO75w30VsBfM4wOA+HEqWN+P/jfeMm7kwwbOx+Xsb1G3
fEXAM8yKM3pdRvMROOsbX0CDfFIM+GxYpNHq0+UQlUpsv4jjKxMF2VdKJIuHq3G6Yq6sbKLufwSZ
aTPtkFPGpnUqVypPr04tFmB/Rwlu6dh+MwFjsjkbuuQ0pHp3gNLk5Yl0bK8yL9j4aHj2G8YlBhRH
s2Dgp6oHX5C+3ELg/gtAe3B8f4i4gV7RvdS+qkE+fKth1OfVted7caCUSINVbfeyb6PMMiLvHg1J
UOVncexjRfIrDu9B9S3MOL4dLN9wNkmI4oEhbRI+PoXSsT3FLpMAkOkvmL+hVF49Xe+OpX/w0Ho6
joVZg+QnupoleEDQL1UjhyDRPNDpgxcYhsttfBxv6Skn86td6j8M5/tQtoM2dzRa2PJwEqjtnRwu
TiAUZ9U7Kw+ztkjg3dsWKk94h3P2xskzGgINO/83EoQ5Cx12xKSgp324lLtUzHFP21ekQLDOlsD0
QsKfwC9/+g0nhIdpgJVCjasegyeodR+NX25Z58swOWh+fQyzCC0WGXF6S6qsGjWKGnp6tYcHiCm9
RRBYcnGB5TlsUs31scnCfLdja6yFFLS+fYTDNSKgLCE59FGu1NCvPHB0FT3xhhR72SuNocq86+fz
KoCPDdQVD1fm9YqzK1VJ8d+hhuJ+ZsRz2jZXTtokYbfNJUjId5OEPLp18rD1cxP/t4FkNQNlW8hi
XOTK0S40zrhAmbxTtHAwbQXllQIsMOmCRg/rfe1UkVQ87oU+3QfhGO2Z94bcz/JvgAdFx0JT0q8h
XuNgVHlElQbfBsKsNX5EC96KamFeeB/sYAawAYkQNI0+YH3c85uHlmlZDgyj7SrR2UKtXi33CgAZ
3dm7bVuBTW3KHa8efP4o/1cRWtpOFwSg2dbfn4QR9vfWCBTQWWj00X29m6wrrhkNP8PxWPBvhKH1
Vgab6keWxg0DC5uppwkPLqLVeFj5fhuS9liJKnA5jCi3kp+pMGNR88EfjJW9eKgHwTA2Etp5t75J
Ccd+w03/8zCUAxJih7+HTjUBCn7uJtPBXhxE2C4xJ0PNrvhrqoTYWc2XTbNn0gS0J7hwCDL58Iu2
HB5C3yTOuGFgU5wLXHztfx4kDNYjle5+ZuACQiI28ThJ2PmuA5Yo5wROslmu+Jv4JP1tCcOiFUbA
b3JgnDGzxOR44bTZtLJrx6kBrDbHjnZkqbpTb77i3/U7Hh3tVyjHDqyXuMFplUWMsfiAABeX3aes
juaCC4ulgooLC8PPn2HTc+4gkERQle7x6Gt3KHYceMH42QsMVmuoYNlra66d6mA5gG4GSaIMWwDl
oW0ThKIS7JeTM4jwltGgEOZpDANUbKvifzDi+sI9JaLK0e78BVwzyVLEvLuH3swJTpgtq2MFzI2X
yjih+uVbTTw5XfkK196aRDkIgC/FVkY2tfzyEAH2zo+0JtRuO3GGmJSAvG6TbzJpvbLfrCGYyPqe
Vd8zdyjcstDH/QbbmLOcFZfEBt7my34EdnJ5BmRQu0sz9dKj3IoHihngRGZDHaThc03XNDO/T7cZ
xdR6joBWWEzCqmyvUERFngm7/zGL8SJw+bmh+fkl+uk/x7gDmbVLypVZzkiO0ia+FUWKnlxB9btS
rBEf219E2GLgIxRgZdVUa1aLjXuMQabdLHXMos7c7HoOXCuiTCT49r/gehnP6oLlB98TIsoEypmB
FhW8lVaMeZhY0VYS+QTbXOZs76jJbao9DCnAOOZIVcJjDJDEQzqwQ/8RLQRRtl1jvOp9iN1yQ3NE
/q7UOo90eHNWvjmwXaaThTVEnVMJTrzCUjM5m2VAOl1cdxROLSRdL3hkv2F398QIlRdMsP3L73Ay
LELYTyqsiuYXLemtqlQuvQbSVCInL6CWHPh+CrL7Uw5XSzW4VHC+X+JQDEonSagNN5lAgN9JUWY8
JPRKRhioNJyeJEEXnYmRCOPmQZeLdSXAtxn37uUUBGbN4R2MborhVr5ssYt0oWh1odENKsakYfTN
PgjPNxpvg4o/ADPet6xuo7xjwRd86F/5IknDoUSQTgT5GcMq1hZBenW2v7ez/QL3eVTGZet31uyk
gfnGJJf4Zx7MaMstNDGQtDfQqWPu9a8pFkdX5XClHH58CbYKGrqvy1lcRi59jL06YdV6YpCPla3U
UBPs9EHL4N+7Xjr3/LgYvqA/rCLJhuEbiOuCdlVljDCokAzxBa5jstAYcq+ah8dYsJp48OMfOHEX
dsmm5srIHhdKezOY7I6srqoCxKvEnDRdiB0ufdr0UJIB37nOl23RW3J/NP8FItfe0QQ4q6h1Qet0
fW98HTSOMdX6XV2VoAUUAIC8t/ASgsOZXqqXgaGadnV+Q0Tag2wyYSKhhQgjZ684dTRsOJLfpngP
dspN1DnHuFXtjbELRuH4Z/zD74MM4QqCeElnDjqcxnaiuI7d43vhi682xI/uPgp7LZ32ys1YLH3L
9pWSvMn+hxPzzxW/dTIs17HJ1WAhI/fiXPB2entE2O2NFpUbBZJubqmWUHQfC8j5xG5tKhPE8nM/
zQ2fe/tAxvUfFCDV/vNE6NL4Hz8q1jw4YzBacj2J610FbdHcJh1RgngyUVVCf221LYs7XJMYV+MO
70HYX+As5M+bfrflG3dcTU4Xrwgwxo2yoOcKtHD65b3d3IGShd/bQbABWqazX+R975JbG8CQfxR1
rH8xAIp6Ok9DsRXUsDCZaQZvBtYQ8Fd1hg1rmQalbU/CdQ90+39YiDiGuQePgv2VB2ITFmDuRV/C
uN/O/wjvZkBQB/FzG2kMm00glcnlp5LEhKVKCkEfUeNATZq3lJpdcHdb3FNl+bFfcV2V8bBqzBUM
f0QV1deMBeoPiVxfPBqEVrS9s6PKimVKnCKLubtlIRPZL15EDETlkWytJC1+ZpQ03SEFyj2D/DNM
qb5DWhzlLFSD/6FkAU5SHdv/arPhDAAVbDdZccUDEhLAjjIWN9W9GUQYtXcqfgPaUNSFhQcWIbzW
ISTjF0fwv3EVADvj5MsNFuEoTNAJgX7yIkJ5gBpgEV4hgbj9vMabgQjAV3jWhW1X3oaQWIoOy7Kv
Q+HVBJVvupyAhHg+L39TI+03S9jSA2Y3/vgxxd83qqljPpBdev4gVNdh6//gdorr9ii+Wy+vaAjL
0myaY8/6yA3AcX6194cdrlyzwttOALf3gv0/vkSWCh0rfHhM8m4u8FmITH8MC9ZR0/OrJ4OtBiep
d2qJOkFfQpAovkz3+gnNX/W15z4ZCxdgrly2keVW9OgSqKrsVfThqO4CduC0mT3S7tYGwJfgtISS
f3YWB0FnfRtR+ARJ3aHghmJ+kWIw1AQ4NJQ7ZbwxxOcn+Vd/5YlqJOTRTqfjUTSnQNXbITUseIyD
ox/piRPzJnGrFKc4OfQ35oNo3fjVDgySw0WFM62056sW0IK87lYf33sdv/W8tOCGj49JsPMlCYvj
i16KG1Hw8r6zui5V//Zu4T71y22tzF+jyLybQBaW7k9BUV4boJ+5S7tnUi+FfSHhv/toDomX6yyG
07Gi7KdRAYkGIb9vEMOs2bkwkXRNfAAqbRyGn6ejAnT3IHyunA3VG1S7T6zWQ9cRnz1C7pM8R+OA
/+a+ddRhHkTAk3Uuq07BodmnpQxxpTVL5DOxT5aQN/1EeGBMAANFUkbJveOurddfgy7eYYxIevgp
m62P3Fe9LheDgOEFJxf+LYo8TOAbHDle5oPSp7m8TGPXqFpASzi2tNhHzy+0HIAXEvqJY1rJoa6D
sYGh+TdYcS9VClnuaHfZQ5ykHOsLHkh8GrXPBpKZIfgN4mWR8HmO0sGyOEyFAVkbd1bH+DqNnQWe
uS+qEuoslwKtwPMHDeL4reM4AOn2EPm9R784Q36lcu4nckjeLOn/okry6VV4FCmd4l4U4Z1wJIpK
i41nfgSWsTQe1xMGlJuLjdA/xjLD0SS5l9uFyjxOMXEWIJJDRY+j/p7yFbqevvVPVtndBhzoyLHj
bsHMJVgk/7ylRmtV6Wgg42hv74LrA+ZSO9gAuSBb+7g7OAoqHtsP+9lhVAGkVv3l/A67bNckck7b
qNw/xcPKCxJFTCuLpjKsA7yqqK0V8B76KSfm0TiVjeBnsA5BCp1LovFopBBDVvi0A3B4iDC2WpXI
EYznaxCoDCemevgN2qBaXWYsRh+Qznq6P2DQc3ylJ4aFsnTlmwnucVKNG9b0gamIzsNaYWuoBCyh
adVDj5I9ZecvH0Bj9JVk53FG6S98pj8wnHdIhfaQ1KW2abr7CI1ukD/jWVBGf1KNQ4SJO+ocu+50
YD7TW2/LE2T/gs+VhTnJ+wc1f8rkGgvSgxKioERGMIs/Tlz9XhkTCpErHQngaFxsRsfv6uFoN3ZW
dySgiQ+MtJc2HgypZvzl7bCwdZaFbNubWGV34bi8WFf77WSfgNv5yUu7lt9GAMHjuewr6cYoIyG7
GqoaQ4N3aJCDVL4OhYhpvkNAjF0dDmVuwoZowGsV1KMSpOIEnCODx84vSlN2RC+7MlxOB7Nttnz+
8Vp5VtI6F8bsQmK2RYTxawyXUVDj826Lj/FrtohICeinB0CkZCqZuK9m/tRgFPB2fbhNhaxj0Dy1
sQEUSiL+eeZ+w4jb8TIAqvD4w0FWMr59uUEjFeYJCziSUA84iFezebRcVeHcJ8C18n/rtaPQMBX/
6W1q9vrwU/Y96Dy4GuZJiKe6NBa0ljmLC2aEAaMulQaqKS9+Td6cIcvym4DeM2tf827B2qYSqL6L
CEearOv9j1d2KVqEGIoICbg4HfouiDc5syalkuLIALQPiJX24Fk3+53Wu6hFibgfFUoozzWXzL9z
gfOkr4Zo8wHg4tmVDFV9XhSuO/LP0/DpiliEuABID9tya/bLysiCMJy/+kDSC0hELXHO7Bjn9XrG
38gDIIUU7vNyvHv5Aa3ZCZ4Gqwrj9SLOqTkMAwU+NQfpRHcdih2jht9ffZk+i08/ODLPXBeTaTc5
OMjLKIfFFBqUpAnpud5UFJYxuNX12CagUCjipMBtkh9BcP41jDlKp8GJgrMm1vJ5e5Zv/ZL3oEKz
+2rOYJ9ha1ijW3Ng27XpOnRI/8EOLSNwZt9LehT5dYcH0L9d7Jv3d+TMBMzHgzWs8d9EMHLU6PN4
ryi3sltxQ6EtBgeJX5QUjb8RmUwPSWI2rfc6/AkfTUaDkQLq7C3EGDZaxyGh0RVq/OhIgcXp96Kh
65bkWMCqkTHdkGe8ss3l4oDnn9N2YoOQOUQumybwiSogKv9cu68fm/Jneq0YqeKKOB4KhXhDPHty
crgRosCZod6JpYrqS3VUw+BYgAjuAtBwdqgzm1zRXMeZGk7p9MU+/EdsYavobGRVdCtEBwXhl9mw
DmXJVBsjniz3CGc91WrkBDYBHL/Rm2Q9qAliLyWfnhsXMF6wN5DV8rGGO9Wb5Eb/h6ddyoCR/9zR
wNqZlqhsG1VSMucy2xMlWYpN0fnXLRatBUXbktQjPyMKeQ7UsFYD+AoKt8YvkdXki9BLHU04PonB
qMM8p5D5YR4P0M38nzt6jszLlS6BdpmnivLEGgZbQrmtNEkLaMsvWlYBN2zTsZKPaUC+UZTB1p7Z
ebafJ3v2wPZbrhDMUeHYrcIZfn5xZ1zqayPOP1DpdXRhNxcDfnAOi445DgGED3dw5L7L7V7Z+RQk
Py1AnJP/NBDLWAruLrc84qKHhzdJFm5tEXdS09wq/2ZAINNDvaJt8F+W+Vi66KI3t3juT9FWhJ10
BKKB4mP1A6v4mjPObA+2Ib+kuB/HSkyAMGQTeOB9CEQf+5ENL4V2+s20ioX06w7t+qcci4/P5R4e
RNF8v6KkLCnxJMHb495FmA0++pKJjzQBJrKusw/ot6MKlEac3cOjHiy58RVojvwG2ST9Uj/AkXmh
KldwKzc4oTN4QqXPWc6Fp1pG1CNztWA8uW2nW10tseW5KxXiNvq3LQNvBO8mls+RtgzjXZwwl66U
XTMVJNrsJXYm1apItoYu96iXdSrbCNzLysxwUXB4MUUihLLIhyBvQ3KPBX7aPx7/YmcF5MfsgPTm
sahRMnivcXbbBNyenb+j59kU2uYk/jBS6LCb/Kghtvz0O19hDKxWHgcAWI4nxEQkvn4991jBlUEv
Y9eD9VZpn7UhniwrY7dC9Bmpuh97A92RVDsn+vp+wiy68dpj1UEGaVBwpmJ4pat9TMlfRoVp/olL
gunbgqpkW28n300U6WDmQQvTZ//iK8a1gnawJfplM4bNLb3G7l0wlM978kTqzV8l0f81eWAZyMHl
YDBiPK1iIWwmqHhhg8fxH7IB0cNwYuOSJA6Ps+Idbceska+PS/5/XvnGalWkuPYfsNHk9017Q97w
NdX5jVuucdVk3+K23rWZPgK8AG/OrxX51ZTdLWik4OTQi3TRf6qC82UJpdY9sbLgRpW0/h3DNez7
SLmCy8rEduf06pAnqAbyzma0blWxAbYPtkUeCUS2D9FcZ69THvumncXlpD2lmwtsEX7800E7hKhR
2VtfU/VaEKD4ZfU2kbtpvkIepXrGqnbwya2auWZi1a7TVZw3lst1ad5n9q2vvcjm+Gw4562Yt06N
EG+EVsqHJQM9TbYQ+aSOYHbOh2/btBrxEo7EpYjXj6Fii2UuG8oY+yAfmtt46GME23XBpe9ZQIz+
rJp4q8p+ltq/8PY6Fe86wHruUIwO7iqZqUCG1iGuIFxXmh/wB0N06/kQuWqEdlaoWKSlbw/CrtKO
7XctCI+kCVvoYb2AqbQ4CZeANKmahyNUTOSRgR1Y4p+nGfiFvaCTcPt4d1TO+XO48JQKhGShsm9P
HPzMgrHJ0aDZEuSwZ57axRJN3xy7iWtIfcYJE4l5KBMGh7nzm0KDMw5EJctcm2BGb8ad3arzGP1k
g9Xk/aNHe4KuzkBtnGWo+j71YlAma8Xk/h4IY3t36oxF5eEN2cwL0ZUNwF+s/wN8ShKS8PvP/VS7
SVTvTcfSUrU9CXhEpwqOaooktl9P18xZ4pCVvOuQPTRGuOxg0AByGwOJbQma05fP3nVeLHeD/Bp5
GlDHlZ/XUav0zA8Wc+HnjrCYstTFSi8ANKmitV2iz9j71nr430cSWk/ToGbSWn0qeuXIILZTmvzD
yGe3uTKjMbSqb0xC6yx1IkUpnWadQQYw0LFKnAEtAdnJojHq3584WmNrXfDPvsrn2SZfknIi4Wb/
bX0r1fM/UvEMbCREjerE2nF40QpqymcvRInXIwoUkKmluFtl3rxdRQP95SMHlqH5Lqol/UgNsQW3
7fV6ES/P4eKaN0crtJBwd7/ylPHFAB9zRrrz9CpfWx6w0rTF61a2XULDQlisTTf3GmvBrVxd4cL/
dbFJA86pMzRHmAUSAZvWJSc6W4RFUI1DjZB9ZuuixEVONKHYcna09GGUOMorOJF2f0gAYQvJBaq9
luz3rerWMRTv+MQXMXPAk5h9DWm1JTaraOUwk5GdTRlLZRTFdGHeJDnRPiYYRSJlltByn4bhk5VR
LbweQkNhvuP9ajZe7BXhVU+CIVkpaZh0j11/7JY8CeDCBL+KPhHIYGXrFyXqOefXZY2EW+Uv6lxh
mkotEf/xE7195+Z/x9v5Yq6Yg9fj6m2eKF9k6M1zub4aS4GTYn+MBgFbWB7lBifESJI06vh2vps2
SSXlz8YDYbkSMxjuthSP7HbyfcKchQwLbekyhuXg1Ko9YIozzSRBIhToZ9HSbJ3m4ofNirSV/Wl0
II16b94eLt804H+fd7MQZbVGvdhMu1A7Plded1cUC/57uP0zen4qHe20z7R8mywWEJCnFy9nNnYF
GTRkpIxZpsW/+ZM4vrhxJmE9dlCQqZn4LMFGWVfeAYNmK+SCpzggM2p5ik0M9BAxIebi1p+p6fil
zQKIpNEo4d0Ix8zcvVbvwkend09H0w16wlXufv1XU9u5g1A8K0TbQ01f5qX3X7uV/PJg8RX3JjXz
wEEn8RDi+j2HcRbj8jnv7qJAH3n0hJK3ZSzXiS9O88zIyqGC+da5PiXxSOGBD1RYiC8lrc7+SqCK
6FnyDZ9lon4BGZ2P/egWwoQ2zYE3be1LfTmR2XaBMDAn1Jv8zXE3eCug3c5WItGRUHypZ8Bt6ouC
4ORUEH3O5g8lQ93M0MoE7SrD1wiEH/LpVJVzYkCjsvHEHn55YxZeTS1leCH0O/fo1BJijOnbA244
t9xYHo45XX5i9XhuYrVcX/gD7/g7Nb+11oSN1wxa1K3JU7LGOgDQ5pU/I5ljlsBwLJXAndpc6zjT
MPHr1yC3wnSOd9Y0AUV5HrEyvSllHD07fzeBTDrgQQgAJcyN7n47w6qYZWbPp7xUPO9DQ7aUsUgg
7TDj9I4CPIocs2d3vgj/7oybEFlsLlp1mtCaoiU8UWm/6CMwdJGWC1Z54d6P7f+MKHl8+WLGC6g2
XOZZxcmJXS/zgRMWxYm5q1SqF0+4HpxDhocySkMHZ9zUYB7e7saNEXpDVXd4TQiGOQEtPYf2g71P
VHzcSrooRIVOuPWr2YUDrOmfqml7XSqEWMITx4ry8ZtRsr75/w1YSG7EPCK9gLBQqWi15ONd5yT+
NMr0PHaWOSoobuybYeRH2G3GKqaLmaJ3QPn2YnNR8E1djL64b76pBLL1NMvi/ljRdTEehG4kr0xC
mYKocizrP3i0jPV8ukL4QdT6JRYWOG2X7hh2rOnIGKPuGaKJhMIiTKcVVNL+/szRUqe6vXWvv3FA
D2Oc+rJFcFTSq+oZIzx/Ujko0ldNpuKEcl0+xnf+SI8si0G5psG56DB1GkGsRrhJOOVdw6gt9RAS
2B7iWg2WGVI51ilBKbytYzPMbrP2VAWF0AqvMMNruzSxdnAMNY8wdZqG7YJ3j47Ccqk0ntLbsTUf
K95cP+DGHvdJDJP6wRcbriAANW0+J+WhwdMfC/vXPaflMg7DbqjDhnqlpJMZGfFAVdYsJ4R0b13y
vyfUlQLcMcGSmRs2JmWm/Jfmg3EEnYg7w1TXjPy8bwg9cf+b7j+C3ZFZy5kUupPa3otj1A5pUOFs
Gf0+k23mmlrEA/sDUO0hZ1FAKGH93xe/WoYMu9NaWvarqtcA6ys07Z7Z0mXY2ZSnqLcN7gIG1+uR
9ddATTrycupZXZSkiv/mgoyWA0PJGJx4K4x6uEyzPhfSS4EUz2OSsn3052BkPZOgUkUmDDo3pY+B
cw9sZm6hWuLkMs7Wa8Y28F+jYzWVGPPk6tY+4+oX9I997OYq5Rp7Wzc9h6LjJUoD4me5rbSvDy3J
sxLWLG1NKMhYKd/EJJs8YDiJ2F32DpUmEvwB1RLtgLRFDgfnu196g9dHsw47TCBEWO+yMe/GmNSL
AZ3j3iL7SvuC+0ytB3MPNvdN72VuX1wxbiY5YtM6IPmXmSMVSZy6WZ1WpuviYJOyIiA2VkrCNFL8
vHjwjK9BePD/eVTumGmPdLJvpkZuWfZA24J2iEdPphnDXmugdGFGwOf13Y1cv0A+N0rYHjbX+a6F
EAHejSoBlxK54exoOvpDXx9NxnffT3/8aBj43quKrp/ZiOqidWGgjz4dKX4IvZI8DdV5LFxHK6kp
X9w3pBP4SVusFXW1HeTrgwCCwfORZVwjSTD9iWxVPkhrOlksckMpcDS1bR8bvqdikuO7iKQw5crJ
PKnCQw9dOjm9CK6+3YpCRxFwqhlt8eoE4ITAZYNGVnfuaPR0kah1s5YbfCxXBkKS3fTwg/feN2um
kDCSXva9JDb2FMnukg3OQZWKr8WzEEt1+alkbaHq01CD/5pTzXtetqj99BOufJlNLX4dyEI0bmJT
F/srzs1dRN40w4d4zn51RuwlVvEqlgScZVyaa1SJ3XOFGCKfBFhEwzInrB80UoGvvqk2kqoejHzz
3cfu9rK+iNMTM+8jSSRHk1VFr0T33I7Z2DvRnjc07QB/xIaBABt7I2Po0+cQAWKxTiPHGNRMzQBL
HSPSrSXXzWxWpREjGnPSQkTWr9fiuUgp6+2JSyR7P+8NAn9aklRKt5tWLvWNJYy7thRDwCtBuvAs
RJNcX1hRvINtfNZiPED5d1bt4mdmbxAlI4eRuoN3gGtlpnVWkhb3lQv8EvndMlz3sXib5RatRNaA
n9R4LuF16P3eHP/T4gNNPMMRjsxG/pfRTAXJlB+rYGYa29i6kb4Ny/H2OyddqcCtIFjzPHdjcyWU
6Eyx9+3fSap43knpEUgtAXmrTrHH07zpFHZxKirJI6nTKDe59REKTVZWtvMRrrHojxelECwkWUjz
20XiMjIwruy/r0WwezNjZGe9rhKo4yFe9xGsALAqBe3Oilx34I3bqVsLrsa8Z+eztPOYg62UTqTb
J+mfW8i3hp7R5f7exOcy8R+fVQrk2DPf3nXcAYJdgQKvXGa41FJZhb/qaJxu/2TzV1thjOhkZpub
EaxE2oxNUCV28BC8e/CGk/wgw3Z8xEHLrADNFxOxjiUOYVi11NU5/UkAbnbxFkMJG6vl2r48DeKI
QSF1Pm2GIe2L2xTRG6s78qgQWvst5iatlpo2C/vDKrFi+1417ckwWE68iHw7w7RsuVknhVk2tOo1
zL4PkBTHJns9V1MJJLHZcUEMCvrA+77FSLQrrUiflk8xRurcFb7Kee0+n9AWRKcMeVfpbGvEUrmd
r86bbp3cJm0Md0kEjaNvVoE0pUNAN6gbGAJG2/0FDJyhqePaQhVNEGB6U9DZBARSLsGkFLWu1bcC
BPelIPj9nyrPAe120fSIeNRxHH0gBA6ZaV33HpMVEemzabgjYlXqWEBtD3Bp81ovhZIHWq5Rq7PT
cTjLEz2ldaNOTExITcb5naqKWQW5YNHcGbE0ivikiJWlVQsGcnAeXlWXgzKO/37CzuGcX9/4GprJ
VjQ+5GECQkmPd2LB3CcqVXcSHemJ5DhWADPbFPKZKp27ilwstVfNaDqKt2UB6A6IQopj1MASP0Wt
hzZ2FiJzaD9W62REbYseVtUEaCvgNYzE+rUp8NKcfuqdq9jqoGavH3uI6EP1pfLFLHVxtwsRYBib
BkzWVb9/Pr0E7+tlABLjHFkHsgkUxOD+ivyTs5GBTzG4ICPTSLViqKtypmHdZt+Hn4SHoilLlJ0m
Y8cxpcSKDHlpfMbFUBC1T+wOrvDuinq6JRcgreq0yCDWG9CUtjP9PFCo245AOWFqiM7e4KWhND7u
Vi9Y2GEUdDmEJA+LRP9JV4Xp7LVcHlnwLKvoEH77bAkT0pXOfxR/PidF32av9NVPg5/fwUwmTvDB
s/ZWTPTFYf+MFRmeBx712MckVxcU9++Gk6hEZXjTDK3jxJ76lozFKhhz5pcKReVeSLPzftTkOSpQ
cJyS03yclT6qUViuMtmF9kRk9dhnpWmW0fC/gNXm6kf4XkRTN3mJrjLEWJAUDKfELY1C8iCrC8Nd
XxzAcpBdVWIPDdHDD6Ol2VxIKf+MufMgNghLQDhenGqGdS1vg3JNP2cG6AwjGbMX02yULEEChjIr
/a6cFoNdC9FrkzCFmjrWj7+Vq9AWg/mQTxE5HWaQtM9eFmMwg6X/1r18Ekc2h97gFHqmSQcFu4BG
CpIf5JlTZufBgoj31qrBK3+L2c0/j1HQio6ccnzvuzz8x6IbziuUK8JsmMU4v92SR73qEWG8XQDS
/qCBdBGBHP9QsPZvKcy3AND42RQGnQTn6i7O/pWMpTYDVK+lsldiX5p166ZdYd+Ibr9ygifvrajm
VFnu6mPOnapO6xni15J9O9eqOCFOCOxTk4RA7mS182cKY57n7C4DiN2JQoaMy39mQ+MvfKdfyScE
FYgGoPwIHLsvlRffm3jhcZ+QPuH05s9ZiN49JAxR7ph/+o9kL78lLffUoMM2Van9kcvgYtW1AyDO
zpkCIiAiaewhgYaihcN5yfUWxxq580tIJvZ1CWcZl0k1h/REVhv13WHcTH+IyjZ6XBfJQ4YrHtvp
YfdXrEyEUgpKrt3EbDsVQS2eMzDiZSiMqQisSSJ1Bt5SQWIPz2w88L0l9g5msPZ22zsdQ1UaB7zs
mKornMQzUmoBrzByJdS/9UMgmMK8e6+4OaZpHPGMc8CjbI5lDICSI041S6ra8VT3MLDnQJFDGUaX
iJv9HxTaFpD2nGvo9d5Zanlx0f43e2IAMkssFrSSEju4vzGLkOP5/8pvLWC3ntu3nN44HGJlY7AB
C+pzPM2K2a/1K0SFomoqCJp02Y1YkGPlYELoSpR5FkQlW8DmIbHk6dBqHSmxM1/zMFMpN7pKXyFT
tjntOAWSWAwOsEVX531q9yu2zSkLevXgPSlEMW2T6igWcpjNEhnqAY1n0h0S1KfIUC/bNVz6/2MZ
U6sfYYoBRPwkgIaH9DczSSV5pdpViB1LYZuyPI8ZU37B9epfXS0WMEXAN6TsAl0KT1VMUguUebKd
jkkHutenHTkQt84jh/Uh+gikjlDPSF7oXmADjvAYqx0EFdk6Wl/+xQcJf5zDRItxQ0JHBOcyGJXu
cnBia7YEUbZIUTyIO6FfyvWg7SNTHAaMRnyzuniezGbojUcjHRa4ekFADGr8WxH3Aswk4ZkgZYAs
YBZqZdYa/QaieWOxxwaq9hjLMm2wUZwtFrlOtwYpKc0iGoVK6EVk/nDxrbY3fCLlFotclugKkpgI
+1IqohxPl7akya5BD48ZahYBBXA0cLaTU0zkHvJ2ALP8NlSeJlBnl4VdXnZ6ei7znuD4YSHu70HZ
MqHHWfLtGpQzTTdKcWsRsrCWkkszZqBhKh3nXGIfuvZ0nFWMqPZOqyRtsqMbKvuLjLhRCpC+yAn7
nOEVyOAT0qPPH7Kiw1/zbvsFfEsJSG3BNb8cVYLtQZFx8U6iGeYq3HHlhGvSQWrO22VyVEUCsdZV
3MG7yzv/JjPEMdV2or9sezk56I53SD+PFfm9GjfX3SZULXA+XcCCahshgm/WlqVCR1rfBuIQaYWR
jAfqy8bzg/cIpoeGoStq/X6Olw7N0dDpgZ/n0gspooj0csE8X7iPjdX7I7JKGkxqehaOeDRgyj7t
Z5TDnUH/TRJnMdrsULeqYQG9OQPBtZViJkd5+9A1DTOtAfrdhKEHfmpXhSW38klzRfRx4yLznmvW
NfmprLwGpKwhQWjweI3Iz9M/62TptSPGIwvxgrCeVqpRy9DMUwHLz7W7SO3emx+FBfyi0TW1/vDi
t61UlEJUPIbWK1QoUPzADgGGfsm8IfZbCJIjFDT4Q/rSEECr79g16XVHi3Bnt2Lh+lAbwUsKSKlZ
QwBVnPXufwN+dSshpNYlmFB5zbc6cOLKS/Y+A5UR6c8icUYFWoytqBloGkol+O8DLCuHQtW6kyCx
RdtpXNSrehULrueLGAbllQ4LWIO0rHoIyohgbnt9Kx+e/wpfG26TeBOMuPZaUGMvFA0VzYwTCCav
cU/tSUBjF67FMHPz3U6ISqxKT8L7qu0EDn8ur76EHJZd73ZPeGzUpg0YCOoi9Nytxff+G4jd0pKN
vetZm2017czyDC5HvSCYfcFAxn4DC8naVFn++43dx5yzGlBfc3paDP3zYs3JoUmLtQ/pB8LNFBOl
Cdyn2wz9d4TwSalSYNFwrGZjo7I5bJkEqROu0VsHfsbO2EVoLZ1m9lXy5DSsTbeLc8e3fjyQTn9r
cy8qqGt6++UW4AvAwg7Bhm4S4xgttoUmin8dFFem0nkug8CPOLVmDb9IEvYeZC/uxZK8ogTmofZJ
z6yh4ua9yx1TBDA+J9d/BNwkUf3H5lhBhiY9fWPwr1FvfZpT0nLg2nGtQix4zZ9gnYaqD8XwQrqm
AsPaQG+kRJbtutdAi/HtWQe1MO23CFVg7n2wiaIUUTqAjaHGomb9epPGdDyx/2x6lEQ1r6Iv1uI3
sLolQnKIknZp5uxzcqXaE9XT2nWNlRedHk6eTsL+xuVi/90uTnegDSreMVyVKvl0JnUYE2LaDJC8
mhEf0I8ByMylQUvMc6TSpxEqrH9XTkz/TZR6Zo7TflfmtKKMZZgwlCOtOPhcaBOtNQZk3qsYgkGm
1H+S0H18kmT4MAAD12h1HgfJ4d/8tI3TShRsfT6JI29nvzWVW6bqXLz9C3oK0Sw/fxujlLBpSyaY
q60bAY1GsGgrXD4F/ZAGX3MiZ6cR/4yCOmer82QMmNmNUORRixqEE/N6Ktzz1YZdJM1F6dLe4BD7
Y1N2WkyLJ0qost4f/yDzp6W5mPyEofLHhIaqjp9R3HQtV1sniO6yFkWDcTNN/er1n49UJ4VqwXIK
XjR8K7JRMb/ULqJXVXhHTuTsuPQRLbMTcgJ6ZkMFv6/Pfq0G/YC2C/6XCjcvXV9rvkKgdJhOqCnh
9aziugSNh1JsvmIj7azIzS0LDQx7Uy6SZ0eKQKyaiapF+UOXBXzFHGfRwx0p1GMeuEotwX9IZ62+
UvlmAErUWOwvMLqubtrV28j8lZJPLsv2JTGaY3BWEan/iQHkA+JKiRDjR5hJ+BzmpQiZJcR1VLd5
fbg66FxLUJCPzvIU1g1pCHJs2YgkWPjSetm61TahKHl1iz6ZSrHyUlYvJI/sspjf/l9M4f2xJIud
ko4PP63KGhnaYjyfdSg5OeKlbBPi1V/Yed/e7+dVqKOGHpDrQuIG2dG04q5DR+6yFso9Lc0HbZXp
169Qfa6QAbjyaLVALq2NGTid8n0WzDgCIAtjizWrBEXeNfK0YQgKFSVfaRUAlBbFp64UdZcdTKWn
NtLCNIO7wHJmyIFaAHDxY8am7j/+qeLCRpTt8F/rpnkl+T8mJMp5zN6cPlZ+TYJgV0Nw4s1gXHfC
IXj8lFpUKFZTp6hx8BX6/0oIUDg2uIy5pOdYiThwUnKScoVi992kGzSMFVMumstNh2ORaRI5ndxs
cNjub8UogePcWA9bMIbptKtKi0stfmejwi+HQjBxkzClsG81xnc64MDWQbsxHVl35UuHiDdZb2tq
jkCoSFcykY/m3jiJwwGYzI6Ew2LrDx0KXuWjJ0MftslQy+m571YrkOf86zxNlZWuZnjXa4Pie50X
rXm7OP7KJeRVKLMb0Sqtl5WE1xupPGwoi68fS//UdDvU+IUFLsvw7fqNf6EWXEtDovlE8lD4SI4p
5UN/vCGqkrmOT/+95QvZRCjJtl7lhs8n1NGYhunJnG8DmuaETawjgDR4rhZu2VWILroz5i0p8mv8
qQIE+xjL5S4iihHpmLkhxj7PqGieK5xMJhETuJsDJGhttsQK6qbOEw9WXiU142bcXTAtBQ6A7dUF
ZSCVEys9g4a+GbbVwK+O2h8viobiulpdzqFcJz7CFeX5vWmjqrc7OqZKM4FAK5F9s6YjktD+xEd1
f8CuAKC1DzvMTKuGEo3tfwQKFo53zuV1Cr+8an7fh23lFY0FOIeL+V6kCOa+fE5YvI6wLaMEaCIs
BAyDvSDomxBW/IVMjLv+gMK2rVHb/YYHTZ/pKP5NvP5DsNNk2ciSyjyrELMhXW0rDAcQjo9XJfC1
EqM5y8yzbo77Xs3k5VdMC52s+HeQIm2HZQmmpkSlCck+eFlZe+zQT8Q6vVUL6ShEyQpUzrqQfKHc
/SVVqcWRwNwyC025VJR6OSCH7VjnU7X4WBdWPnVdkpT1gd2Zrlm5ekvJwd32BkFI7RIfOAzc8a6J
2xpFK5xhm7EEYIYWqSYJ2Itjsfkaw9x5e/I00/aYvFxEFShuYiQWBvVEu0dn0GgGXPt2M43bfCtd
uw3lznwbzDxcHw4YNbBATVzslEgnkM9ddoiowY43hAYqOuj9Hihzk7Wet9LmjndRmpqoO7NEZHKw
i6YlHz7sXj9gKZzEzd4NtX4o33pXzkx4swV2uBrZzvspirPhhnOZcsDasoJo1DItz4+A2UbCl9g6
dUwb0M+RWAmpuSdZHkAY4LlO1Wv+J/6pngWIrxupkcxktDnNhAwexWSTAXddOsI0rClZ9EMoDNyT
1WRCM+PPpHI/2RLAHtS7kdTGAzaAWMYITeChvsiRTUMc5xvTKN12f2yiGXMFf3gcgVXVrtRL4ADx
Ovhztsft/y7advaKo67Gcs3lYFngu1Iflz39xR5a8DBBAjQ5jRS5iCZ0o7hjvyEMhIxUpietKrak
vd4obaFWN2jiJilraezjUeGf39/ryyFG3qVfBavNlSmGAb/ejZ6DsjpDbY95xM+JQHLkjeBCn5zZ
CFaqBSRR6XvjBpXREQsSzOFXj3W8TAIcTFqZCmaB8d6O/d9Y47xkt5jq7LyQFabXiyp0dJOkFUh/
7RvfH4/BEfPQLOoFQKolbsigd/pKgA6LSJuzuZrZ553xe8suR2YYApS4waWaZZ4iIi/vl37Vjx8b
QgTTtFSnA+C+THKn28T7pyYwzaMlYlCvEUAmm+o7VqBKGbc4jRjxck8FZhYaa6XJhvcoQKd9Q1Gb
8H3oiGLdRzjibOjpUoiaTJK0zoIBQiG74XoIqUcti2MeuwUJj6mLbrIKeV2BK9fmIGVqPBSTPF7n
5VbTJSCsPJZv8JK30SCUlXSFdU7wDZ4ShfFbaiBMmifDQXG6tvFHV4nvJFCYzkl0HSaRS3vPTrnR
GhWD/kRd8kgqZsmZROxolDQRp033c3PKVtauZV+XyVPVCADljeKobNVPZGwkQKP6izXfI5tH2v+2
8N/aY9PpfIFdOqbtTfu9n6zg/TP3s2GtQx0syLtwL0k5DpZQuy/A6MBKnJU06cUMA5asJPOIqX/L
BPB0FWhFJYHsmZ0f7QPmnsB/sF97kyi4Za7ztad6wajV1nPRlH1xLDKPrGDwaRsxgsgjoGB4n8xr
cAjfIrTEvJ9bplTuwy5jcUCAbBLTxWs7BoAJ/AulBSXFXhmjc8RMw8WO4Iv1OC/ZmkbNp/xKH/YV
2T2ux/6lVNOtKwautSJWgtjbNPJY5979KwoztP8g1BE2z7SPJZQ4ov6C4Ldz8XMBRSihdA56ZdB0
CAHq1Ykx6iHAQqzKfMp7kBW6SSGinCK63pmTw8TCnDWvup6Yu9we1Bns+sx7BblkQUki5MMW1T77
upY2n+bJkYLEVebA7LVfyJY7aej4yKKIx68/TDHH43kQP7GMcEIX2PnEG798bNmJnBGpwUXnk+Iv
mV2zYJyiQL/QN6p6T0jIM0s070WtCrjt/KglEWSfCt52vooUQ/tLo55FL9OUD4GMF+5qqvgRU4gu
nzjjpx0BwM4WJ2PuiGPxW4mwCR2YMj4ORE/44G3ukTzOPg62Yo07r+ikQs+v5XobZS7mV2Fux42d
mwNTlJ/eWEjsv9ZzwNmiEUZgtQdbBFImUhRY8FgJMvk1rMV+z/Gs8L/AQf/YBaVLnpDCIGDhLEo+
1ZX0NW4d8HZQG42itOHy5kaJ06HSDnLsD1sj/agiiMzua9ZHB1qg7plL07Kq8u7DasiopANivI3y
pf5nKy/5F6XX9JbV9hTWvCccy6rpBkr8e8xLVb+UgPawWLQXHUj4WGBg4WpLVtEI1MTLn/08FCao
hejT9CgI4mcPqCpVUcevFfYdVNyBxZq8cDP3Til4/f3k0s6gbML7jkxTmxFBQli3CMDHsfxziOWM
TiNNG1pUgH18QpaAIaD/608k4yt+vQgqbQ7T0uYN39XUrZqrwvSosonZyCop/K+RqtyBhLLF7Rab
ElLnqJ+krpdNP1znr7+diy7Uxl4wUWS2gRzfmM5QCUCFEfwdPhKkpimcKIAlfUAYzgvV/K+2YVi0
CzVawwzWtuhp4FJxvMrd9mIO+ihGHB9opUFqFgbPOXPK8F/Zc8mZwgg664qkkPflDB9zAtYAw0Ru
RQupl1YkN7Mhs4wFR3n1fKbR59Mq7ztX4T2V39cHICJpEolQnlxtgYj8Tl2LJqhpKdoAWNxxtl7K
aef9HP95AQDV7560BdPOPQt2UfpsjngXB5GhVl+TbG4T0dp3bgm6FP2Tol6cb0RGkU8o16bD224t
lqJBth/x8z0fHEr9NC56fEksEm58GYVKyd7XEXFuGh/zciZJukNRLMwkknAXZQo74IQLRRXotpjY
ZsKPyneCp9pDxwiTsXE9AOnZzwNpD5yWNGJzYkAOWyCVRyWP8xwSvLmI++0lkhjqriGaJ/kazROB
pakvmYgBG1Li+f59OVTcEn9bObru6S8AXlW4AGaC8I5sC4bneO6i6KNBlvivYsm72RSLg8M+r1bO
Lc/OqHrd6Ffgguyczwh2yJh9t8n1rg2KGWf0lxUYs4laoG0dQRgS1jMzCWWreh4govj7o6ZIX8kd
XGonVw+zEUwRBncZAte4+YRZIm/K4D/zn0LO411o0Prci2lVPS9ZB8DIILNUgueZJq21tt8HGnNG
16dAJLuPSx3eWIrkfad9GFI2r6XOeAfgbTq3Tld4eumYiWrdCQJC31VG/S5eGY3jHufmr8HIcsrg
XGg7O4YjCeas0fgKgQ/j/D5ZsNZaLn7zB89gIdnezmLvl9vX0qlSGezuqi8+ugdEiZLtN8bpQ09w
ZxThpxuhYDj+g76F92xw5Z9edKVnEU9zDqgJ2fnLpxbS/FnN/1K66WDUTRCUYvj/GrHou71g3Uee
EDmBl0/gxspac+Icb+HhPN3XxuNCTI4rM3FyweTjPVk23U0zYTXGTMVbFx2FHfSShFTlv5mpwWtC
kysdLOnUlbXNV9S4JprY1/rw2EP33/ienzCw2xb60y3iUiQFQ8YmPx519GHWTRg4pI1bqrFSBP/C
74pEClcju7D6GJ6k7TRMIgRMPWxLg5PKcb4LE/nuO12EuBDC5oIMvCT9Vl0oQ+lWjsl2+HSlKLIe
qbqkUTO8DL5QYvZ+/3yFUwiAF6rIGAoyt5TjQ9RaN2W11cLOz+krTLzvWz1mmah2VoMmIr/oxWi4
7dwmwhBvlTE9hU2FL3Nt3EP/lLioJUZf5eIjjmTtIvvJHekkZoW7cboANQA/ai/ZQPdjyIwuWKnI
4MljkF0qX7RWL+ILR8RLsqckI075AKaqDa6fzWqeTwIzXz8Sy/G/H4V2z+bI8sIiH8L+D/3dzf8k
n+LhttMpm1g1IbPjKDSLc6n5IMG6jTLs85/WluvmGgAoOBv/SBnvx7iTpTdeyrXqta60QXbqZd7I
6wgJ7S2OE1qjsWNJIPRry9FWpSmvKd87PWNTeCmlrP+whm3k4dM6QoVaaMt6gNAXQK49qja0AHEs
RJn9lubxFhC1jokxS+Yua7GT3L2i/5w4xZ7iBXwZngRJwKNl7A1ZK1oRLY4AXmYUUYkaSJBDUGFr
aYUmuke7bDiurfC5ltBS7oa4A0GsS7n7A57wYE+xbWozDfoL7t0lqVc2JSjhauWVM8GfsafMrMJa
gjYr4RMMWM4z7NeZoLNjBMHZi5sdrN8FMZKwXBWA4P/rMujU+P5yzH4/yBYCFLPpLem4IXZQYKrZ
/Xe0qJ3omBIUwroAM/9AQWRfCG1CXXOoWZWf79fo2LL4UCjEnbnGMzZtyuGog+4UwJcc+n1Vsh2/
dW3stjh4CKrMDpnxhNtyDbXVdA0tZBsIpeGls8QEfCiG3FWSfdoeY1B+vWFVMVv3vObm4AN30Oba
6aHQ+GsJ6XdEnmV73/om4Hv8HWMhOr1M424cKKMBv7DV20U4XOKoh4ITsWUONPjXlUYe1myfKwXS
szBoce8vMZpwD4Zy+XCm1URuM40p/qGyef/JeMfk8suTkX8xmcBkgvikF255xQ1ydJ0G0aVwI9Z5
7+xV5OKpsSY6JaVsg15QBqjF5o+VFQPKUQGrmoj4nCuuu3fnrfe8FrB3AP/UDRUg0jECsXub7dSl
6UmL5KPnrGsGkECZt3xsMhUn9/ytYMX3cRLi+38LSjvBKLqO8WYCKUFjQS2eEaHDyd3JIej8nCbN
QrPC6wLdor1po16/XidU8riMoLu0P0b56fY9nprw0XDV5m2cbMNv2fL2fHyfsnh3LgkbFzHC7X/w
ZLs2vKm8ezFKyLX78jxd+oX0ResKn9pWYRgvf3P4ALEDFTLrzyRdUyk3F70ToBQf6e+Gqhrh2Ith
sAn7+Fuy3KnlHxNNKL8BBbOiCc10c692EMop+/hO60sldJRr7SNmUFlW1bKvRVKvW/hUHLpx16Fz
wZHbwZWjDssTwp7a4N96PQ4EI92214lrO5k4kxxH9UkM0mQkiK3zla5nQE1xbmXsSVnYDkggBniw
dPqJmq3gz0RP56+/zHoyhZQoeUww+84rC/qmmWjEuNwzGXUsimrg2ZQn8sQxB3Xhfb0F+tlydlw5
VfRPDjR+u2vAEZ40UzlYx0jQJUayU6qBm180ECigZ61Ozl1fd5vgqkNC+Qd8U/zA/QpgzPebhJtD
EyeyFwlwnSU2vuyQ+jXnQKxg1nqeTpDqjSg4pZhyypQIkhhsDg/C/mgf21XinKmJXBBuEYsmoqTi
efGK1nFXvOh1y0p4GTpdXG3rdvp1ZZHfSl5lkDneSsx+zbopqGkDGIkBtHVBHb+YrV0UpFL/F2fF
+uSUeW6GENi3OkkKZ8nC10VjEv5ey6mJnP2vyKf1+KRDybkIfVVS4/AsL6VDJ300Wi23nSh76dY1
OvYPUL/kPy4WnBv/g7B6d+YDNZc4nCGXCFLcp5gqRBEhyVdOQOUHQQZSMATDJYpzMqaZebx8DaT/
+hmJ8mn0WpDKO2J+M6nppVHGfpus91l0oM8SuSY4UN+dWstcPTNzJTnGoURqro51CKdJlDLF7gIo
OKMxHyb7+j0FaozT0DYBSdPcvuuS+U8wzxFJo9eP4OoaPDaGNZCLMzUduKj0qHaUbXVbdt+4fIDw
O0Ne9vgfTjHXhegQGfDjWG9gEw6PMa8LLszf/HWHQRMNm/eKsxQEJqz+yYqjsedLlL41HB6hGHY2
e2Jiv5JklxXe874vXjlrmtsW6ZPVLPKvFLTmyvG2+rH0ZSA+3XXjPeA27fVoYok3kFjePsjgCbd/
wwGejM5u6amOWJgTlVbgFXmsMJE48q1uDRT0pCbQaRzevf6FrAUkkG3gmNeM3e/Z5ELqNAUGR432
BIGZngusBHcfiLQEkMj9+ZkEt2r/mbK0ZM8frM6MX8DRnWJ9bI5bf16E0aZHwWYWe8tvTcIAJSSY
A62cHpjxfCnA0mnpAxe8VDqdbXNbfbfNh485IhUerl9ROmNyd/pHurQV1zstopcD1KCCt4UQHfYF
q2jHVS96RwqliDC0lv3g2QcZhQiHNHWMK4Rb1QPOIagMHrAYPlC3mwiOZqSMcdl4nbhgyrUaJA/9
8I78yYSmTCToeA2srPt9Xucmkpp0rhqNZB9xrnqMviXMz5DqIp6cvMXQZN1Q53Dc6OC23SlV4ycZ
D2ZlXjweEbaYfGE0A18TCs1fuQGFWvLTUG6ZAoLtMRR11aDJULd+IlcOFJhaM1wvcgWWIyEobXpZ
hL4icKaaHq5+j7868cjzjWa26LF2yg376kgGPdz8rGMDku377N6zglg2rJZxJyt2AFBDk9QL/QMM
zUx03fnpNhtBZvGrumMD5HToX05vA6CctNa+eH4OMlNN7mM6WPh/vcVOZ7AqrWbL7oCKxF6yQkUM
KRtvAsNffbydkEJqL5eNVblPKKG2P7F+IfLhg5wNvXaCqkoj3Y50qKq82+1jGS+cjCnExchTvbn2
ZjK6yO4T90rpRxulOPbLFCM1vMLJp2jReUyUoJ9ENApmGv69A8D4PEM7CVpUUKj/oIGYxJlZhuPB
g6r4nECutDYElGHl+uDK4gactw2b+yFxDwuMYbFV4BYiW1rvXEm+DPepoXO6qb2JqkrOkRoIOnD7
iE0Am4jOvYQXTuVVMFd50nmSxetsaqC9844O8JFRMDc05gKhcwL8UEbdeSISTzQyqItGFSDsNigb
1Fs4naYMgN0oh6rVAl6D5eQRoyTsTY5J6IHnycLw/lzrg2H0r9gcgiO7noXqHIC0Z4/2glX9zzmO
R5bQFWOYh118s3vZ08VwfiGurUooln+ilQgAXG07Vh97ZRSn7jToW9UsvcVO3mQqiKY81/bBChO6
tIgzBJ0mbnt/VcCw0A8P2TSsqrw2z9cazHCv1oMgh/ezfAlvHb6wh/d7mxwmiSZHMuTTSLhHviHt
/9k5pk0pLFptST7ZlVl5XqvLzxi9z3xsNSIp4DX4bdxZohbc081Da6Ra8lzWxChU5fwMbYGWvc/0
Hiq7UT030pxPKoo8JkY4cWnbZoUGCwK1MVaXNWGzcg9Av+onJx+G09W8tLdVMSAJ8uxbaNaOia+L
5kNtYUzgpO9ZjBNBx3TyroSt0oJZsu8wTEhf/wcUzX5KhP7rbiYE5Ea8p7XH0K1tobIpqMZEsubB
9D8P6kpg6802WAnFRo9m5RmJSOqE6oGKn1mQUgm8vblWh4ewoPfB/2muCYysYh/boNFjQ8xweWvW
p3YZMAYY3hIl+0Ypq0KzXZ1l8/YgSXcJ/OSx7T3/a58NHBehexblMVWE/Z17BCgMa0co3z+67/Hw
K2hCB8E+RJmVxx68VuftycWS/d57nDUBJnB8GY4m05L1a50OwQ1tdxMu2VfE0CktkUgP7ja1LYbO
Gry40d/KfZ7etcfmAb2XlgTBRaGfbWU2HqFI9Pu7aRgfO/HRKtbHuWHPSuAr/dV2hgYOSvG0QcWi
0yDyUGHitusfCW082aP5H0+6f858TUGcfKHbHvA78lL0eizfhySF2g2UyIwBVY1T3HTr4tWy5ek4
GjfO4tPV76HmL6PKMtbfrQsqrrG4uvhWdDWh2YdyQq5XTkkfclslKvooSAZGJdepUdFLuiVpRTxe
s/TJebGh17nFdv4kug+ukuRul+MbO6uQF2UF4f/A5icZmO5WNPjq7oK7oAFwrSytq/ZJs4ioCGNA
dupGsjcRvUaFpK833GEmxMna+EpsmUHZitxtJK4XkT58nciXET/V+MX+3BgsND30jP4bxU/8RXb+
LSWvjsyHPKy5WVteCyS4llwnWNFztz/KJTPv3ffVJ8WyF5P8+d1qAnzYWXR5iT84NVZmaCuMmwav
dgCsqxhBoXl3tE0g8LznGuJXL99ztjIlmsR3rk/1CBuF5bpellURcMA4yIgs2UJxebSvLcE/lvll
cTIa2sfXKISsNVEYMjwxRS5HgTyTDCIBR4G7OYwp5YyCfw0epkCCr1ujXHxBlAjgFpT2RrKGaGJL
mzTg3CqRdEpIjCJvbChDVwIWXQVlfjAykiWq3kwdFxd9D+Gb6UWCLuOfEh8EjvL+g9hLi2wgnVHQ
+wfhHYtpZEPj7nxz5DhtnHhXVNGGo2pXZJPHsSb5RHvd5yFeml9WkEiapV51RKmv3tgvuSGOJacp
jlbzm+pExSEuTm185Zjtbo8PMlrUautmwUiIxs923kdNqaNsq9CEjE8zH9KRWAb7q0SnwDPBQhzi
CHzwyDlyGHOTCPmMIvQPXwuNBBJyGxSsot7XO1iGj2IRDr7NIq6D11LATHHZxAK6E4jAj5R6Rfmo
LPdnafENWGrELU71FZ521RRSR0nky+nUx24b9w07X5Z2Uuo6zYLHgILrWDrm37QCUQy2nDFD4Vj+
V76zj/8Q1tPjA7V/d2+k3pFgvjXYOMVvqyQmnsZUiOq8N6BpWicEXp7qWkeKhlIBCS+xJVQcj78C
i0OpZqKkXTmimpP2uV6jGZbgKAlAtlfYt7Y1VBrMlUaZWLwjOP5XJKuo4DDVG7NU+yErMsQgXMfv
ydGPP1R3qIpih59gW43DgAJWE8QABDI2bk2RWCXfcM3+JJ2iMKk/kz9deh9SRt3BbsnIQcoxo4C+
5Vgno0A8Gx17bbFWt2bbSVJ9SCRU91DcsMgaRmrAPb4G5CYAwN5xt3x0sMx+lpOxjSgqeMIsyC5u
veE0zYORX9Uounf8Vn8McM3ftd0iYIM8NIQxK8VVRiBy0Au3qEncfGrPTujCfgbo61N1E/T7eE+C
JfN51rWNOk+IBygy41OsKgirWx73KUrdKGMZ5AkFPXtFquzQ3KGt9mn+ji0NSKeqI9kbgl0cGyWw
qJFiyEmlDfSguV4S1km0nCB5wmufXYQLyV7uO+dZKlSIK9tsM+hTv1BUQ/8FkfNS54vEDN6//lsF
ZUDwobdQpk3wCushbQzwwCjdBnNwr69pOPLRNkdFb8IHZJT3v8M5D24Dmhk/jacjp4gol6OsD+E8
BPANbPCDZ0/pSL9b+cxBvMVBd2QELAdRZ1Oy7LupJJVDDRwmyf5Tx83S12V5PhyXyq598+rW6gbo
e0aDkMVvrV5hqe24GajTeEGBn5eaz3aAz6nRlqO1D7lj3XVQSgcEgSLde6grM5VF8UL600Y7pFkV
ETeLDjueZRV/MOAO+jP02pwg50U8EaHnhX7vwtH5adbbyhhpT8OgspfmJABAPHOxRPW4aZ0kfqwA
Yn/ozQHV+Cc7UHC9YWYR5SnOz7FLPNJTbpwWxnFCDXYzBdAdiAE28734vMjt0X32qBSTGPUc3dJM
GoxbaBdUYJ0KWCEBiLjKjpTPg3WeNkKfmVzbMpOV3NZp/hgx1OEj+8xfRlWObN67HwwqUe2AJisk
B2H902ZXm3upVgUOKGnLu8tm8y12xJuYUF5daB0tBpXE0R32sob185TCJHJ80VEOVC1wwZphf3b/
7o0ftKdQREgnyw54dQ49RuEVdDos+apmLUPTY4Wzx0hrOa34XMPy/ygw1bfBkxtMMy8ac1UXTYFP
ZBmwo5sWGCMolS/1Pdo8XqPN5eJE5db1MaIVQDM5ata8PKN2mnExiFzwr1A3Hm867Ik4Q4d6+sHh
V6oG/qNFFPmgBbrQXHaUVsvnow6tL54CYJSP04SDvYIcL3LSl7OketkeO0V58KBju99cdNFM+adh
lqHiI09Y46R/U9u3UOC9S6AFNKOaTPG4/HNB25JEN3BQYTOEo+kw/beEzkaHDYzDf8JMCaQukvUR
yujgvRBrBxFpDtz/K7QWhWR7B+zpaLW/DnMp7RQi5eYC+ec6mR4B0vrSBO1UXt7N3zujaLrwYw1c
+ugKUii3zqh47gqf7Aopw6TwCEK+dIS5Y9ra2zcIE5rJhilHIr7Sa7Kp/+nROrl2I76nCXvmI58k
oBT545d7o5R8rq3QrkXZnH3F1ne5YUFHthBtFseXZVTmdKSOQ+K1qNijvxC6zDwmDqDmYLqn1n0m
/NkEGKPftG0y6Mk7qJiKye5J6bRMz0aAYrK0if/zJs/rkEb7jfD+khfVNxHPSD1cO/t7FVE5EI5A
b4u7xFj86Xr+iykWBRjvs0acd0zzT9XihRcbQEiFcsHilE9rksAfsT3zoRFmxtwmRJotQAkvqmNj
MK+gGsSK+qFzTXlAzkYRp58icXP0MIvwzYR9EVbLxUfBhRY9FpFIMik1JQqHwFX7tna0BPApubeL
owTQpfHK3HCiuzfDHE1Q0C9j1lklCt0ly7TTEmWTcJ2amuNOCIe7NTJ0eC45hRyM6xHnNT6XdbUJ
WsJterOZhJRKpvnraP/PLEKvf+VsNRCm/imiIkPPptlY/bAZBOFe5GP+J1nRPOz3Lazv3avSOZCO
R2vUgghiw/JW8LgTDChtJ6dgoIJ0JI7EmnWgy0TKLUsBfwx3DkUwyGOOSwDQz4P1yZZuCn/Krd1W
H9Rv5uOiO9588KXjz3LdI3iw7wxNFLxBwmP2+I9b12WOFR8i5M96o25x6lIe8Po4BxcDSzwmc6+W
Y2nbefif8S9DRV4pPh3tMzN5SsxgKbADLFxEYwOi/swQpDfo2mYLafzn1Ob79DqyJOzoeDb0ZlD6
CnpqZ2p5+hzcr2aZHbEQUvfjQUlXeCtj8y0DNkcOZzflTMUDQDRsVKySGN1yqedjGbSMxQVgjTLV
ju8I9r9vLSmIg4SP52Vre9Jjk29AOhHp4iHuOAcw8vkpviKXYKB8u5GmvxZi1C3Imhb2VZtbPAa3
WAgr4/qiJEeVRw6B9oUxVmrF2DkJgnzdPwHFqG2hTsNOqiM/ECCSsuMUuvpeWcWJr63bSqCu9ojx
VT8D0jyklatX4u+39NSVjWyJSWspX842JfwSIrEipDDFy4Xmhjc/tVGqp1cb90JvivT33TDAm688
MRfA12XwSpFSrRsle7qDuk2fuvVwo7Egj9UE7JGntio0qT0ABv/HiqpJPYuenWYfw7whITrONB3/
uW7M7ndXUb5CaCGA9So3H2zJHE0KgUdGe/Vfytld6Tja4SntH5ywji88yXwqnaZyyunpidQ2j13M
btRGxkrCGStxmZU/dYUsiGR+riv+js7+0ctmZz2qN0SPm1dK6OjuV3mx4COEy5XHV20aFOK0ilfg
baC0ok7nSBE97gkqmGJdTtKwehqzw6My+M7yzZbdKMUNPtQC4fAMuaBPNpcvGBWVNi24q/AOQDvV
OUo4qA42/hit3v3rABbbiNO3fqhM94QueTrLyrh3JzRZH/kekPlZcCZ2/SUgQLcIXQ3uXTSDx+j3
BSh1s+64guBHzZ/9IX/VNExGhm5LnSXppCTZe9gI6E9MTRTbC3QPK85r5U71OMNiVKIA1TVnmucH
fYKbrVgKvGAkrGDtgHC2PMYgUL51k5PKh1xmZFT0paXXon3wN3j4jiBsHzst2LlYm8Be2KxlC9Wc
313xyoB5wDKHoB+3kVXs8D4eOSMh9sQGEkM0N2Kap3fS+VpphIhJJslLKRhB1utnLg6AvR8L+Pf8
iOnCZkgstVgf6NOQXH9UuQTRelFKnGNcNPCbE+Kx+PiXPTAKMR/tXjX3vgasrmMv+4qxiaJPqK2p
fxar6sIN3mejMs24UvbX4Mh+BfGmHO8Hc9Kjov/+nebT1Urbt16WcZGseqLv/wYpxtbz++qOb3As
I9jYnoA0afOL3wQ71LYguFjHSc2Dz32x8IQERRQSVtFi+ArgJ01jh8JhJFZJu96wlEv9wyxJUPQ6
SnEtugVMONBwaHSxo7tp1GE4H+pkYz+izNu7h9g8QdpU7WgkPDBj8YcoJ/x8/N2hYnX+ThLjGNeV
TzEAwbgCOgL1u4V3i/fCm9BjtjEWFIeM3XWx/SvznZMmzWH/Jbhgb98Uu+RZmS720UB3Djk0d0h8
fMmmLd1YbtH5BrQrXGQXJ2rOe1AUbOPxOJiN07m94snjST8sNVUUGqrT8mZyemeenbU93JkrV3V9
TO1Qirba+Gx9K1b0o67fQSdGYh5ttVEzg+iv3XAJeE4hKD1JsOZnvNAJ3tdPE5kaV6v/IySHu8MD
LA5OonICqOYpQu546FVGW2KYjXvuHEy5Nj7/g5ZtTQv5DIqGN4JCdG0QPl4YG5IcKjJ8egSqXzDh
X3gBPprKcM/IslArcw5db2pBSKbbZRlBiPyANVdsibuPK22elQvL/4GU3Cvob8UTYVCyjWdmAaK9
eoJzWRRx6wqVguSEnQ1Y9TvgRcPARZRV4S4N6KUnoZLXGLouvLV3EsBaTrtjpqQi0V8xGGHt/eR5
X8gXuC6gl+v0Q1XzLDeJWYlPt4xEyzIg7hOKS6xJGANF7Kj0Oh8pUPG0P8owQZ2oDxExAh1UFSfk
xhxFfZTW7MnhYdiTeSPNTH3UdiVmISuv9qIA00lPi/k70lPsxUrRSXs+FNABaLPsL8mTX0qqM532
T/cYteDXtRXf1uRmggYk55bOs1v5yYsMqqm1e/QH43INig6um8gc65NQz4cJ0KDla/PHxCx8HVMJ
smeZDKU9au8a5V3Ro6uFxu6aS675p751efxh7EEcPySjkiJ74w8Q0xuYiLdqSTW/6LNrZM7O9Dzy
HLL6ndrlDzuSTumRCoUwevM/YQFjhK34n1qIh0fE9SSVc2BbXp2ln6MZBUGLzniAFfGNPQ0+A8+/
P2XpKwfnHo9dRZmcJHayT4EB+y9nMWBjiRkIDEXSPVmHr6Ggf/YsBoACnu6HKN6zqjCUqOmzDA2t
iwXJdWTllt+bY6Aq3krlr9vx6hTjnFX+oyoC/ekU+K/jBZdil2O1hJQeT21WBQa2x5XRncKu+jLD
yDYVK0EFDXg/6FehOqzARrhyvRa+7yYb1bia4gjAtNaFqKFIf+TcBVDFAEkmoXoJywHd1ChH4AQi
t9WbUff3gFcQXf4wi+XvQIhu6NFWCE8e4d5v/90Aa7cXME+N5RRNOenVeH2+oA0TqyQ/qztBaqZN
Fj8EfJhb/OB7TrUTOvzbPNY2Iw65MSvrrlVLcs/75liauW751RCk5v5IBfEoqFuayL7+S1h+sbnG
LjzMQXhxsYIEALSoUeAVDlfXxFJZ5Q/3S6eIsoCJy48eZIR4WeFKd5LD9b6OxRdTIcUrbrlb/lz1
lYbiVtpMBNLYpZoFgtnlshMvFFaJSDGwKuxKFb1CJAciSMI7zs3DGIYBzCS8+Za6cGS6cyOdXLqj
imbiey+uGEpwVDFf5KdUaoz9SQsYrNnsoqY0KwWeK/XQ5HflVrVpdcesnos62/+de/s7lzlwCQoE
oWmhrHDQnIpIRQAQcNxLUXMe42zgwQT5sMpjzBG6L8xG48QgTTy2xey5ISTUEGsNaxz91iheh8zz
DxSqmGgIyVsZ5Ne5ns4+efWbcwXnAuxS+PkUvx6U0+PsW4LoCc4INVcuF/bZdaeUsHW8w4akVTii
YbDhQsbmyLxDSUocL73nXy5Q4c3iL3LSILMHqtryYEuzeyXaaz+2OD1ECDe14eZPD5YfE0TyZ85n
hIX90MGxywkksGGnJf5YWzka3lVd4ESYKhZiHN3zOSEgwm5zQ7Rr971U6FfQ27LceqVCTFzW2Fk+
U9LPWQHKHRJ0p7rsPnWjz9sd87zHjXm0dax+9Z9AdvbKUjBnBiZ9Ge/kD6wxFuveAgTuJXrL3TLT
ZJJ/5LZxgk/lR2g3/lsFMXoKuTZvIqYBP9lxYArJthVciRwSGUObDgrk6pB3/O0hgzIUnNtSTXQv
LSXVkYsGbGAF6YCcQlGbBy+huz8mQc+BFDVGu0Vmy7C2zW3k/v7BmA4OTHgP4PLKT1bwOa07cj6Q
Ni5ikhSSdb2HKeG8wVjXKDc6uzLLSfh0JvHhtndjbnyVHMqkShSBa4ubzkIXULbHTwuD/Ry2kCWp
fmTzgmC3/gtzEcMNCy+6TySGVy4i1XdO7hiAdAG6hq6RMbAoKX/5TixVguI+ms0Bth5EDyHn2kle
WpZgo8b+5tA6epai1rL7mGPjjFPCHrcgjB1UL7qmAi7aIcmYGs3Mk33jwOf8qo2j0bnITcZpWeN4
aUwPtZTN1LNFXY5AwhhgfBppkXpBn13Y9tWZAs3vPdEY15nhNNsSm2H06Py9ExMUt4l3u173F9am
bz8LL20SJ52ORO3k3c+vt5AbD99B5xDGSJ+ku8hlT2damI4b1b7266PQbLacsCmFnitB6akp7oH3
n2IxHxiAQIvtkkJ49A876n7LMt+DxxRP8HuxkvoldVTwwhisSIBq2bBgJYQPVE6X88cwpzge6PUl
fV47tnKjuaVEpSRE0q513tlBNZE6/NmeEO3KcI37MvDANJbENnrmxr1pBAmNUaZfSX7iWgkQmXvB
fOkWXz7EVqRZZfs+TrjpffcKhIs5AcwgDsFNRaip8dOOHcto+qREaJfY9N8v/sSGpL6gop6BDKXV
//uLx10bn4aciDMFaY+ORpBnTXqEFlG509de7UKMY3uSbA4WpWR8s6hetDJ9zR87eo0LGb2QfJhW
th655CTp3y9v1oLX11Q6kTiiLp8/SLBbT05rAIJZUu/NjMq3ulRTM91N6oXmFvT3drIjeDU3GwBB
UnJDt2tvk8GpHeRVCPgmNnYJwbotl+oWJk3LmWhb6Qmin+W0W6YrgwsQOtlQluYqPfUNICxrNzau
AiUdHD7qCs4Cm5M5Bx9Ruf85VKEMj88ow5dB12U+u7JqMtyPjX3glse72pkXj/7fzqSjmqChFcVw
CZXy3obpRnj+7Knw5/ljaK4qXulfzZXtWK8R3XUasq1rEzBBtDqcwYvJz1DspmC+S4wZSqLvvnAO
9ZOthx6YY4uN52ce0OBN5IyVG/7whW0guGiZjsD+ai759yp1vZyTl7MLt7MoHJVimdiUxMz07eld
GgFDdXZTTNaBeJXa8lww3met7FTmzSRM2bi797CpWORJhH5wZWruSpiRV0mn3kpUrfWff4Loi6FY
oLc/giGhBFUNNPPuVEuyiIO2FD8pFkyUnWOLCx2CF9i8/3qeipfyQVvBsWZmjkcPEEJYqSQoA+6q
c+F6nn31PUuZq8PwMhuQedn50xZsBt7OVEu/iUCe+C78agv+jlv8wdHqIRbLot8fkipJKFyP/rnH
1qOHBY+oPEUKZVOA0Bg9u/krQWOLzD2EcPiNQsb8W4x9EqA97hejHlrW6/BUaRg2SpocmIiyhgB9
gYUNhdQMadXnweupJ6iBlSeJz65lCCm6zYBAzHruY2GJGDh6R4T93RNUlOdE5eJNU11jeqlTHMZd
+ZEGlRjUHFOBa+o50wYzfLxM++G6rdcrZ3qPs26SNi4GKOu1n1ew9IScrftoqP/AYsU4cZa1q2I9
nl9o8amhX1jQx+Z0iU2BrdhBsWFXKFlFMxE7rGVyHRls+2boiofO/FpmaK48vgKDJGKEbnvTGIOt
/YLyj/Iq3d6RNDiiMJ+ObjBkoRSli+0cW/5pMpgaSyYjIGtCPbcPcBM0AiExpD1WPS8ftpo22rLV
ZuQr1KQlO5ddU0hkr0vgxhMTzdh/xFoIPuvicKVtzIONurhpMx+sAWjYVNlw28u1MKDGsK3cYurT
K/xvv/QFeKUNgptr2XZhW02sfsd5LHzSwJRNSO8BR2YtTX5HO65EAKThN05uvfSSCrPbZn7DC1rF
Mkv2AJwHNu+yqCaEBGm35DpDOXqUQ5+gG/wNu2bItRKVnFQeIXubV03XUoEgZm03kys+/GZplKSY
sgmADE4QZzMYcu25BJaeGwxQi6QJU23kCMl7U5r3pRLetKeFiutUOH0e0NDujm+nFlSh4/vqg13f
vjuAPVHOuP1AvireMFr2qjh/nEJHcS2JT2vPMFjT2fSgIQmLwVveYfBj/dUZFg4ATPn26hVQDJuU
Mz/a6VPCtDJVTT6WRT0l5Tn6GP4doDbo1gnl2sJ69i7L3ssMeIgoZ9OpxoSRJNBEQX4zFk9E2T6e
T60fWCwm4RbGAx7MpueceB3CRkfgXeCzgJt3zXWQR4vtBxctUSyAHj3FO5GYN7Lln013IfFYtlWi
nPzE7f8EV8B3ahnSRSUj7G+06mZj1Q5MQmDWP6ndYGYU+HsfJyIrC9DPRBj6nY24Y4WurlV7xJfy
MwLNnku5S/d1wUkwC3qSL+EX4UnHPlohDH/LjBFnCvAalUHgaELzHwkF2zpWnhZtzeDjaAVUARdO
J3lhwp812QfNmuadfWxQhYzT/TWfeP/N+QEjk8aGdjfHXcnww8IgXbHj7YmkJChFO5gCfY29eSBX
VhWsAAcCyOObwY/lU9HBQXm5Hg62NVFB5UWxLjcmv0etSHu7dBTNP6MxgNr2KdFzICSm9aFIvNvg
niy2tF7jAmgrpTHsg0p1r7HQiNlxJWrq5wtIwFxQgaB5zhAJGQI7dR5karASd3gAkD6nmMnAphBe
FAKrNOAahbgE4jyxzuDzInkBKOzRxP/i4X/EQazIr3HoxW6YHwXqKBzZPJBt2Oh4ZYk7AiZfLxdo
Vr/XgdCHAmwvq7+859L64WlS7pcUr1iLoV0Xtx4iMCVxvA1mIJxX4xYSt1DLRhwWU0BeV+UeECep
eTIAJElF+MHs3dSbOGoHZNJ+FeP1Ef1JuSI3a+Vg7WdVTHxr1J0StEqOzMzvl4dEMkIBParjz14n
c4d5yVLPyjLKWt6u11vwmKYxGvsvVRbIIvq5oVyQmwcexPeV2Alom5RLtwGV5+1L6l91uuLX2q2Y
u9vu/GuWbURdQatgz+m7Dm4T0X1sKMqlZz15KuE0HS75NJYOuxhPsfo/yAUBTTBKtDaGU2nhVTkx
EQh7a324abwcV5ms3i7gbPEpUKlNip5H3+zDnr5GBiG7ykBvz54jdWO5kCvSENjUVY3XFNWCCVze
2Lx69RsiNp4ZfgrArGzL+5clPMArp0zLgonHlj67WvcpHkdfgDlfykwYkraH1u8lnhNvS6VrZd14
vBfyc0Mo8SnZKUOqC72dFf5HlZv1g3luUUpwfweyYBNQlCueMDy/nzJNxkwq7p91kqbapNWQ+x8v
7rP6yn9IndmJs+gAAz8VNxHxFbiiaO9oxRelLKlNlIIAEY28DMbCeXleStEhozMMLUvk9tOVE2VB
zi3e0TpfFqepuIt+IPP0XiBjphvwOsE4uSaj5D0iU0T4KXmHhJ5/JrDR6wYVGcli+9yJ9WN+d7OM
QSBQ+fhNa/MsZWgWwgCD04mTxZwssFdqX9YpK5iIPx3/qVZk+hdSyM+VjJfAhMYBUpdKRf6vy34z
ngsNHrdsQ0LNij/KbZZ7Qh4tbPTSlnQFH24VtACiCQF466Wu+tHNMyRQhr+ShwDPILJgI5Bk62ub
njPf3jceoCw9x6YGHgEscOab1wv8+9ZJ8mfDX9p9OPbGJufkkn9T6ogH+q8zWM0jYm3L8QTG8ywL
Sww+DePbSZ0mwSOXquXSvk+w32TB0LVeAjdIyUcXDF1XaBicNt0t/TXg2BAKYX2JBvlXcjPyz/5a
mmZLt7Z3LR1k5tdiXU7M1X9W5vdMemDJ51nBik+kQevOiN3B9qUljT4OLeVnZbDQ/8ouF5YlYWaz
4PO3EnxfVgii+gPfg9P30UkYVWrTiRZsDVa8taOQ7KykbZc0Nuqnfp5RAAPek85LLx7yallYHYbO
L1Q8RAFRpmBs/1x1lp6Zj5nIZurAUJIW5yNu3Fu1vadWjbEMNEwiEywDC+rRu53O424twEqbNvHC
7C3pEwHrWQjCF2kH7qIqyLkmCK7C071mjwMtw2bDI0er6Xns6MbTQXestyEOzBc5jj/O1hCWkYDs
PaKle66EwBAOmUrGv+MYmG6rhUkBAeE3koeyxCA29MNjlmraTaXbHPn4D7CF9Eyu3uTEDie+YS7w
mc3NExHNCkoP7DNChLwNRutHG80PIIsRajuoxT9n1CwY2Aad7i8yEqD9usvqYXsHL0xs9Bv2gHjg
QsMjMIBAAmJuRbKqi9s+GQ/GgLuRloP5fEeoSAzyYxVVuaS7fNZL3JOGpLEU31HILKscbvfgnUfT
AiAGMWp+sAJLO+Aj6i08c5oTGCNSWvt/IXJ2cMbmK0ASKdHhMgJqnm6gtE1L+txD7Ryuo3/4Aovb
outVcu85cu5F/zpykkQKVYAKLs43n8+3TaLg1emNDd79CEdODOQsPSm8HWd7zGCgztRG8OOiV/F9
WDoLasa734lDM63+8JoTWMF/scyn2DWjv1BOPMy76koR7RfQ6QQtnj4QA+OR1Cw0Ur7qDjvxpJYD
cFMvicJyhdqjbHUpCgmaudUuZt6A98EEFnGAHUxYzKOTxkR61e2MjuEaIN26YSqo9oQYIrSs9e+1
TxeM80SBHG2sJ3ZPDgWBF5z64WR3rSOEcux3dtgENXKK9D3o3zR3KE79Wu8P9nTEeiweo+net5dI
M+nXgLmG63Sl2nmp0NfeApTZszDmlcjt9x38tPRj/p2ZITxvLYi4A+heWFcesi6fQ8xGBwnGwU1j
NvjALvbDlESUkCbjxhRC1qC0gJ2ASK05QiGxmXm/Hyph9x5OO0ZbmRKJDcnsHcYtrJtiPC4kQr0O
6WqVEph3UdMFLqtFZzh/CxNrJ0Xv7FqnQxGJvnxW2g+tCA2TSBcmDVssSNrAQkrW+1IF+V6/rHYC
F3EZFwc6xzXJu5wKLaucQzieNHSNjzmZodT+6wSK1t+xLeMKRq5GBDeG3qRTC4KKNDU+zl77AKo/
UmE11bHzua64/eGFlpC0L7zqXZZsG4wtWXwygP+cnGaw/rbHCAYDixMWa0do2+WadQc3tN/Z8LP2
BozY98F2Dbwzxwlq0rzFVaM1yaoNt1hYoMOAZrrxAc6n08SdTZvnxiDq16sFgW0otEY21Ozptp9I
bnmm9hemlELQ4Dp+gs8zhrSvmvFN3VJBor2j/v5LgcIEtp7eCxSsrhNg765834DRkCZ94OzJoSD0
wCjuZJg6X+OviB4kkUElUrNhJEqJesiMN4DXDR+mgAIonlCMYT0kyG3U+yEcUyASW37ErkQ9iqIu
EV0kE5WTbYXXViJ7R+n7QpJYeVyqmAteDHENhO13mWUGknirVgTVoK4LRIwUbljjF4XjuGc0CG0S
MskFfACWeiOyjCRJ8LiUamIeY99EcXbQGnLBvB9NPM5jq84vEba6rhM60EF29hojzvARcIhTafAZ
dT5haGaKw9q2rQ1xCYPXv56ieMpmat9tiN1fJZfoLXQYxLHwhSj+wJX6Gl/vHvV58xemt5mIE32B
5Y+vSDzS6IsM76yDFqM9SfdW5VhOdZmTWzXsfVaWXlgvs45W8BJdMmv1wToJSkrGbP8smgK+qKvf
8o3B5GXx7CylJ45JhzYw/DPq6IN1cE5gfnPBcER87jHwWHYVq4tsd8zU/C0M87JjDJcl6TaRQfrf
zGKLT+PVvkx7bTsi1chMKAzKOadYtgTEcKU9X6RFUFy0XkvsNCtVJW6z/QkSOpFf/4atYU3dfKeL
74cB4Nl/rY4fJeXgV8h8TDDLCpDVvL1xzL/e5ihtmSxz4Na8lSMpfpFAmQz5Fjf1S+8K/9G+hQCA
SHtyk8d1myOKOHowL2vH1hDKJm9EcP1lCb+6KVpDJZzXB7JgjjWo2dbaklyrCYED/8E1aUxMxrgF
lINobBCJIwMwDNNhdyj/nby9CeS7yVxGjE9Bt3GtHlP00R5f7SWbPf6iPkcOP2D0cFRcSgk/zerJ
4BxUFI7xPAgD/MKndl1GImWIHtvuBLVpbwneG3hq2Sck/Bx5vvVYwjLsFSwFsp4vNi2yISNpVtQA
W85uAnBK44K0eOmrXhb9zyRQyg30OJIEVj3OdQf4ccA4DrFZcVHnocsk6tBBzn2q3XSZTfV+qOnJ
LW3eVm8ow71eD5TAk98bQp3aDoDSTdlWSA7Yx5ct5xZfrYZt43B4NniQGnf1CH0zGtehgvJa4Qjr
FfHNHxiMx8NMlF3wzzqZHVj7kGhym1Yes9xN0MI0VCWaYUgmRT4NOpyRaNTNJbq+iKnRZFTzffem
ONSFhHLXoICswEKBlpDCIiPOSmJ3UATikiU8IUt/vF8J9e2P143yV2nHwWlr3Y9MUHpeh7mx90Jg
I4Fo+W8Kr0YCnXmsArKsQw9wseUWT+PUKRMa8haxUkbjktZjVNuDNFm6SehSSQyIBWO2sFwYY4UZ
2YNVj4xQ2/7VPY87354k4E9M4nYF5L2tK/+V4XmP4rNomlsRjsG6VOO6C/NbEhFzUESo0CUqy0PC
1OZI6GIE7VRof9Ww69i6oUYSz05AggpBpjZVViHSop/f4RyOqQ7XRQDoscI7KIvhLwA8nwF5tFKj
9fR9iyuNvI5BAu+44i4qbv6W8z/MtcqEpGO56Ul3xFceOaCzbxzJIbWItzBu6bnE5QTkTtbPT+nv
/DJwEevE3Y8Y0JFRznIeihrQUcEa2rcnCQGrzuTSwL0lVLmpm8c0CfzzJp3CsDI3Ira1lhbZPZ59
fp/jwoBW/AOEXR7ru1SuKdzKf/95XvteI1Mwzg79MJkCjIxgujdhpx48K7yEAjTjPUVHZj/xHEfk
yFOxoJsfc4Qs/bN3ArqNN6E3oJeAQhThdn3KDe0ejCHlh0d3Sbf3sbj5S7kZpFVtBUA3S7FQ2rXz
nLYTkcSUB9IH+7IAZksIQ9eNUPzAmgAETzIcflAdcht1KTMm3SZFpbEOzYDhiZ2AK1dSMHeTkfWz
s9/wRxcNmuEZFodYPeFE7OLfpm9ElSZ93EBIyBE70Y114XpWPG6TXrOA3YGxF/tJQEff/atxyZpG
OEoMHX4DKKN8MsTq6IDvocPo0SyRvNwy3LLfqpOq/w0cyAcAqESUWRMrYZXJTMqcIoarlHHkvPjg
RHvRczhBBLobTGjPE+1pICq29awg2sJCE+seGu5Yutzg6+iaKh3p+wvgIbDNBekymIG2YE7bzZIi
y28P34IYP0ZkJN59fNXvSU780Q5o6D5btLVyoF8vDiagOvb5TElJPWBtfdpHrlj22uyCNnjiwIja
sbqoKDKoYbzWOXQduh8DW44QaqJK+/6E3dFT/Xlz3tCYQrHmYFZcvBymfpGilMIMXroWvNDyskTG
I3RvRVc0IH/KDnFP1m1MxufRhKEDMZdROkf3KZ8nbfy0OZxRD47pke3hgrD0yEdtiB59IPIKgaVJ
LrFJZ2wNQ57ZDWrOXuYduxJ4WjI43Zbsr2jQIT/3qash0wgmOQW6t11v9r3Ge9FqYLqCPfG3cKT1
AbfWMtrY8zvNhNdiZO11sd6qhR8cOveTnzYD94p4V/ACTgID6h/p9MoSYBmSbjh26Voyvit7QQCJ
+++sHOUrAlch3OhMwo5pwkV9yhJCyrpXNT9QM0BMp7pYuD1j3TrsgvdWwgZBWtS7gC6l0siJip3n
koDAJxSFOaaFoPuTiXA/ZHduflFiwLjxTrhz5rmDJARsPuAOO3I2MJkuh9DADem7vYBRYWPv4LcW
pM77yqxfVntQYheK54RXH5I58iJ3qUpqJBK6XGSunAxDU41ancOWwdSIG4AUlaIRhAMatz4lV7sI
CJSn4wvyoDbhKqgBLu9bxDRuOyG14IkcczHz4uPeZbFpSOX4ajxqQFdI/HTC93SLAIwSSnfJFmGK
/MBoTc9OQe3DgkaFAXOeOHtbTZSQ1KakoweB8EY7xHehhQbD7YRCzmU9bFMEbtCo+3ikZeecb/VW
6mgGpJ+U288KxkuYK8e5DnXf3IuFjAMUZpyVpKvlHWMhKwIxvFS8fy2RWFbTIIRvs/HCfAD36g0l
Zpd4f7MFO9+dR3hTGWcl94rmQDDluwbPAijtHInpfYT+zt2HradkAT2n+5CC2GBKfty4+yhCNVaf
B9eMbt8KSki1MG6Tda/QQJRU7xgugd2Okbmgp0GsBSxdgVkXCUBFWbVnNPOc6xSd+cI0aKZBM4xG
Fl/xJEH5pCWoGiTv8ZmP4PKS5wiEi8f4C9N9Y1C46qKN5oe5VVHIeaXq2eqxRgzHn6Jr5zyTgmEV
iD6ZyNDL4Tg8m5UCAYG6WyWe+YbxRTx5TiwcPwN+uJeH+au5qhNrpPIE41C/zIPiImgnGCEAz3/+
9xKYuvIx5JWQ7vmXIKV5Wtx4tKL8DO9rULIcC9abI4dOFoW4BKZkP6gYtjwnd5+cuKnVPwwaS33x
lYUttUdTqs0u2raFtF7Gu9PM7jOUxFcqNr9GnEInC17DvuVH3T9A8ZBXurj4ODJGka+N06QbN2Gy
RLrjil++64e9bT3YoQ8ngOYTm6yhKR/z3+7JJ/Ged0BZ8F6+zNgJZwUeJ2/qeEA/obBcCUFkicl7
/p2cokUrSdI3nb5zppyLahfSQk3OxM7zZ4dYQBj1FDjcfiLm/wa/N+6pIfnzr3ZG1q+PSjhWZttp
K5ZTBehrWWYwwIBhZzznmZJjzJbtcly0QruAjKF7V9t8/TpzjIPy1bRvp1dtYnSxovX8wlw/4Xa2
efwq9dIhWz/9TV2HvEBWQxQXoIf9yvmeHl6tcU0iQkpDAnOujfp2gvz4SFQOjs89X/W7iubHVnHF
ao/po0p5tio70jBfy/6+LXfa5x/T6q75aOmOO7nEPXI2tBPLhz/R9nKvUTGnZO2S9m7MJd8ZYR1u
oZ7BtM3q0g17G4xV6sK86cBL1BSWqu2yR7EZA5Q+xgAJ8rWuhAWE8lvl2NnLby1BWzq+T3wySKtE
gqiibGiUZ6NSBkcByo2YE65M5xazOuRoI5QkPqnCHSBE0+C4vXkUr5KIUmGF6bvMqOJHfY3hGbBQ
t/QJHQ0JS3zRfV59aScmrmxSHmw9hP3D7AFsLDe7+g6KYa2ekDeIEDrWJkEI2zNb6dSs+lllhnqS
7O/sPvnjEoFEDLIOPX1GmAD/1SZj6EgGW/uH0/LlIR9QaZLG6D9jLTQ15LVad7Mw7co1ix1sxvhz
uz2cngEnF9UrewuZ6VApkUh6lu1m6qIJCjEimgVNw6Qi62y9KaQZeJnpIrHOL2W4NQe9gPtbLZ9N
EliceEsg3N5je+85rz/NtnvoaMi1UAWg1K/kH1GVu1GLrj14rG81NStCzNS8dBTKskuVMkqgMDTQ
EzX/bFjVDUIL/25wdqN8wRxVEIBBbCfMWVPwdcTWt/D1np4TFdShPXen0DuS193uJcpJdE4ebU9K
4hevuvUU0rdtVOun9RoDuq5bgamwE4ahobZVZhtygw8MCsF7AjBSLDA2o+TA/RX19Jy4HAj3oSSE
ZfNZ6i0JOBD+PTORXJdiUnMskWQAEIS396COCgPI03WNr7Bz5qQCfhPCZNX7FSEBRMGy21e7iMx+
kiEiThymcEHC5B2iBDeFOM9kkKnR9o6mJAIqzsxyMRYL5GIx6hgb8Kbscp6Dd3xl0LKjTFUY+DVB
NvRSFh1HyUslf86e4MeZ3C3/HLhAI4IGeIdHVqWyV4fr+E3Fu3qInyZF1rMSMnWYT8XSIe/dfS1m
bJdvvL1mrt5fszsjJM1k+Pv1I53q1bCscdkcFUaoRkP0xQteJ9Qf4NG7H6qOgx+bqi/USdJT1NGi
lyTHPa2a79B+njcCy3N3W5F9DWl31pm5Qqrf7o0FPxa2BrIpa8dyoS7Am2ja0y2hHzyVeG0/r7mD
eO04VOCFFRgE9p098FvNSLVM18SbQKg3/Q3GS4XOjrSSBnmyzTaIt/OJufzsw0shh9lkrGqPCpbi
azAphgiOp311lzAaS1Od4OWs+TlhBwdakf39z2D4qgVoGSFlcpX29nQAjN910r6N9aqoGcRnP+tL
eJyj9SKMLY9gFCDHbdnguNVdDAigurcsXGdWTGRl0mZtFrobqlPJ5pSPdOIb5QDxvjps2vVem+Sb
wyw2cX68oBE93iNWwFsuqtyAwvxvp15325XkZXMqNOFxUaiaCy5eox8bSHADvXU61By5yKl4+9vi
2zcKw/zLBugU5a41I9i0FqsBsnaGNrzSNzwj0Fr3FYoD+KGzMtdBSD7jIzKKqSHdwDCtNAAL7pth
R2yl8b0QeIugC7blF3/VFdyAecWvFNv75+4dAnC3BbTcbBRAYYyOhSMgAjCmuAVJymG57Qo0JIE0
ULRbCuEh+gPw9m269jRc2wGV13tpmVc+jtXpAjNzvGWyLC3I60G/bMeemsyaXq5AihbhkIOuJgVh
Fx+sd6286mC9FKhRhblpiqkqAGXVIk9tEIC4pUZZck/Ilmwp9BjmYooiZMQwdK7eed0w95zr5b8I
U+icyxrjBnb3Z9TeKg4hxbrP6IkeDVVLVfdHKixTTlR7hd42kZ/nP5HwUqRIKZeUPFYONbfvu5jL
oG7H017z6Rg7NBrnk6X7IlOejvRDrwx91LSETY+30FZojR3ATK7dcGXjUCt2RI4Q9vt2ZppnUKYD
1+KUXm3bwpVv2qF2sucOEYMz3prxK8vexXQLnRWD6oma29H6+rqeZrPlzki1SCetx6zM7zm4M5YY
U2h3jYMxLpOx3GyM+ebTG7apR094cLFFwb9aFHSuyPK7fKEX0Hk4B4qViAOFIh4kJwuNgeiliFqg
QRXDvRfk3KAL8C0gp5vrwXgIuFrNkjb/2XZVPPvOFEpS+46XXygeLHYBMedEcodv9+2x6U4pIfqO
9jN3C4SArf1zL+sFn9qvtsYAX9SsDNJMdg4VkUoF+Lo9MuNFI25QmEfwvqEbWb0PppXwFFGnDqSe
l/IaZj9HSabIhj7r8ek2+RabPt2ZlOwXFiujPlY1VzCvDTpQRfe/hNvITeoCkHzS/XdGfjbxKaJ4
+OJPFzwE7Zf12GeJcN6yqb3rDPYH3CIVA7hlz09BDXHdtBqwZfNil5XtuuBRBKw5JcTN7RfLJZQ/
usnKxMRS0Tq2Z4HUrSfPxfJzIsoRWi4KTXF33hJ77pVIdDK2a8r2I5RLMxqXwzqUpMocvb7ybK/m
5MRl3kVgCls5+CLiqEnBxMXhZN9W6Ft8+ClcQupgVqjyHFlVCbCIXOSci8pWXEPpPqj1YQS8V8tN
uFXFL6aAQv9m4qPbBAjIXr2i6acQhGuncEwYV+F5gwXzRzQCmV6B2ccNAlk9FX+M3a0BdjTQSNqo
dMf80byqiIHVxrbu0W/0c3fjyc2quQ2jin6fenM4qFo36ZfAi5Lt2Y3F0X8ABLjbl1tqwI/eSgLe
I+JI/TuXZPskMOAN7EaLf7zPKMRNMFKJ8R29CEl+NC4FZgnT3v9wrYhkhn1jwtsyvQTg0/kI1HA9
L60oWZgClFVqMQl65/3NRI9j2H2UYlFaHdhRYYOMkK+/wRap/TtdmE4Vwiyjw0IIdQZPMbV+x6Ch
TIVw9t/h/CZJ30n9I9K5scUVZq+pgZguEYjD1tsAqawYuSgLg1v0f4HxpXkHerYFQ7QVztxKHUd8
9bmsMvvnvGdDAF46wYHuux5QkimXBtJToLeQiyt/LMuI7FBfSWWUgV/ozwojUVAbPjpkb3dlbdJr
EzXypbSgR/Uc/Kms+OEjzqSGogAPydpJPQTLeW9x9bLC+UfdCCZHgJMTUBYcGt6fxekLQiGyxAWi
bl5krkGJDBjk7zgg/pvgoEMelk72j61JYvpayJdSbvQm28KjaFconTSGo6mxFXFZzOjFC4h2dHY5
m0OQAV35F6e2PpJlT/woFS/EZ+Z+ulCIce3s0r7IVniiO/mj/be+iYTZjjkiTqoigJu9lHNwlgNq
87jhjIu60CMAyX54Ht8TN6fgm8fLNMdd0WSQoAMac1mE4Je7/+RlvlzU1qSdQpcWdmFRK0lbPZc9
PYMCTQMByCS59P9eCapOtEebP+stSjcvhmIFemdKPAqfccjlolV1j5sM3qeVzzOeilVznTwl96tH
UcS58RppzRbYTovn4zc9wyZpcC321AzOnpNnxkDqX37CfHe+gWGwviOT5OoRBeWS0iCLbeOCe9X2
O4R0dirT0rzh/uoCT40LAXyhUw3jDdqJl7owV9TgueOeV/6SPbSPJ5llEGbYS/J1MUAe1+vu491q
ZNMiFJOpy+a0HvruMGfY7PEn9idPDIeWd7kAijcEir6+TQJGNCveKd6p0jINMWoXyIM+fTxs7FwE
zB7056sXk57y+hutofuVoraaES3kpU5gkt7OGDUJZA7Fw3Detq8tD6Yy6F2g2QV/uQNQ8hcZnPZi
DR5JbXtka4vzZOdnXeUpBcM/sY04UB/VCvo2qjIySNrUz6VK2sN8fWaVPc6QdGib2y2UK8RvyoD9
yQjpjn87kdNr6KLzZ7OIdIhIzRfsOTz9dOcrwpvFKOtEzcg555YPFw87gmSrmU0H8nbqOhaVmT0F
Ie7ad92A1KLpxNMRlqtTUulYaejNBlbh5bgaEdzgsUCb1eCOYZK+8mfS3ywYAN7ES13JmWyy7k1P
5z6BR8yLjgcefUi3QE745HAzopOu9T/VxZN9gCXTHdzK8nA9cODuF27OFFaV7JwdExvOcwE1vGRM
/LHweWvgmzMkMrHpJfFrPWnOBdjRlNBjXBfhqqx2yeMy5OA54c7EwF1ibchtE17B1JkaFZHDwkoM
VbUCiWJp26Pyo6W04J/FctyJ0UuTRW4QFKXd6v/afLOjsBDR/f9G1nOkMv1HB1auEigeBmSB3MdB
aoC4njBo246axqf4ZYy4hdaGJgXoPCW24gkAMTGPhPOSwdir5C1E2aV7VmWghSkPaFvURA6RSHQV
XkTALlZPb2FnUw4qk6PyVO4K9mWLA1wo/Ciriv71hTNTZB1Vyxvet/zeFHxOP7j9d45R27S5+Xq2
3mNbXLclhN/Fy5/yIIoYc40tkClhTHI0CbVJxLNytYBxQkLMQvbpiluz0JV3xb4n6eHfrK6pl5po
tCjgeeizyGQqAtoQKLQEhrP4cg0Fv1BGC0I+lcYkT/Ds+w2dAVeHhLppauZ9x4xmy0derjhGr2HM
vWaiq9jh4FJlwb+qiN1O2tLN2+JzsZ8ufxA2qdWF/cI36wcHhtqgYo2w5azpmhdzoKCIkUNnFtIQ
K5HZiJAZgqDPmbUnPD1yYj4yE7800+XR6hgfsYX46ZCD/4gzMuWTL+Uu/CPw16XBrBjaCwH1H8dF
Rv51HAxSuDcSHW6QHcuwcghLXWU544pTXcZweNc9FdFrpZUHHpzINwjK/7MM+NyAnpf+ZiXoUE70
cS7gxPi668vP65a7axlzt23Ds2UqBb9GuX1c4P/8b2LDoanDNA+87vyC6y9bKNvWOztiv6fKmxtl
W57xQ18fKt/3Dun2l5ojNMbUPMS6BDLArXRGtC7Aa6VwWS4MvFFgxmmgjqIHMQFJnO5pjx89Z6JE
rN19LWgRng5ibb8Ue07ixxpWmNRNf5QBcccD1GL3Bqb5+gSonM84X21PkdQYLxI8+bMuVabZfoth
Sl41wQ3knuY9Uq0Ues6yDXlQDgQaVI/bmm/6xsKfttThmbpUKiU5RdWelGbbiY5PNN+91VfWBtaz
yExMCK8XT2LPxr0kdWlhsWPwTD0/S2jGFj9rT3Kdh7gk1V6DNsgkQPSb9tfx23WAwph4puaLi9tv
j3Ux+mRVcysxMceH9RvfJ8kHesMvktg/BvtlV/SG15wIJEUQNCBaCdB+yI97c5GNMgB/4oDqfddM
N89nVFCihMsF8f78Wkd0CTWowEBhOQsg2jPnwoJbCjwkh+QLcJ3YE2hD06VxcTzbFk/oZ62+IZQz
Kd13FLRWArazBSAwkAoJqJWmKFsNMCN+MO7H6wNGf8U1GqT4IURhp/9hHhssODt2CtFdMMS3GCD3
zbFfoy88XOZ0TMngZ2FuhN7Ihs6fI/huMutWp4BQ2d+USWPxNmIpT3MkbG3xqOll2WrNGsPHc23i
/63IViXC7yp8aSR7INPI5pra6OLyqaAZJFZ7HcZ1riQPZmrmF3LVSDCLlBWSwJg3Ih+LJF3QqyX4
lEBsMbMDsrDd00eB6BEHHLnaqq7qOmDEcyfIdf+BonlJ5Y8nLYPLWa2lVntCFDy3LUcYStILpOoz
wGFbVtz8SJr6fqdc48BToL6qZStDQ32lUAIOJi5/LQ08FnHsVsA8HYNApMnzMiLcdo96YMiZY32O
gTjl4myaYBRI+HU6LrCf4l4A1ekX50WKpPcNynVNemto/xwnRKacySmMCPXOx9yaNBOshOyedWsl
RRWSn7BfPQUlZQxCy+kfCZbW2es0mwet8yymi+opompB/xbkY4OJYEdCo00nIgayj4798iP/b5iN
zUuTdaOYw6ZyC/VWLAanJzJGtjK41+DL8kLzDyiqR3E2LAyvOe7FY2Q9TOpShPpLvhsoI+rWa3kY
JfdnC+L0dzD1CtolbBLqJPZrH3noALGI3Vwic+OPlRuajw9UIUdwd7xS2EDWvDFy8k+i+gH12XJ4
k7H9CO11Z5ZrG58iDC8PAZ9H2KIEWAuZ/eB51ft+GrHcDGSu5ZXlK+YMsEksiNLAlW6T+5tizm+a
+fxGmakoN9rSuiG9H14+HxdYB6YtytHLPzUUMyzPr3htQ7oadT6jV2qoej+1ZBAyEDXS0+m9zneV
volFi6l/5hL0b7i35hMBcsRoRMqbzrGqhivxOGPUzzixR1/+DhDhszm/yFY6U0dqGvU27D7dVdX7
MWeGkl7zaP7jnjjcJPIudxsnvDmY9CGdglrLFhanp1s1Bo7uVCyRhXYjTEGlCCwKdYQT3pnseBEX
lW3jQl8tQ++Y8Vf6lvaglyrOn/0bQ+2qFqO4gcExfdLEv6MDG28rlVGEaqb8nS7Zzrg9Jny2I6/j
UDLypTVaZ0oschrdXzfphEIhnhfGh3FBKyBVh6j2AXhdgc1w/klzWIKktZWLzJ+eDvN03bFkoJAh
xjBbDMsvm34z5AaMjz05cSkgpcX2+d0ZpcMxeMHrfBYtzifj/2qMDmvYvsvQtdWBRQ0qoYRjOSLa
LogAeAe4+HzfMQqBwwiE6wIm5epFVD6OZ8siH+ewCbWXcv3HBCFfSM/x1aFESO0pCM9S4Cq3xCI3
usPwjDnQtj9Vu+anfzc7G/rGV53SVQvx10DELc18s+RL9rpnFSWBqcod8FH8QRKV9hy7woXuKC6l
SBA5+xVPx9ebcSETLWLKxi/Xpy3EZmapIe2l2VRD5fJtjwl3BEMLUVmJYIZSD/i2+MN7Kft0IkSl
btO8W/4Q2YTd3rMD65G0JBpcIUbhXXRoZCiCGjXK9f4KgyvmdX+/EKuHDqrFvbYAMr1qP9hqY9nh
AXoKPwYZcwJmXP1x4Q4BQD/6hFrwjnsrmWqXiFaVdzROwS2YgAMJXhAAETN2SZbnmqIQfkbLCY2f
vl71Hol/g/5L9A6aK8LbAk8PrSWx1rdwV7VTtUImhFmqQDNdlB9caGmqH7L7XzE9N0gnDX1KH37V
XdL+If6iLT5V5aCodNlR7bxgX8+B/rKgvntWMUUvvXo1fivK+Md+4hbrw7HF8BAGnIzWD+zsmyKA
fTxQ4DBYcW0QMUQW4sWPtVbFqw5PNUhKT6QVzPR72j9Qc1Eiut/vWM5l2Os2IACDws55daIIFFRp
j0QuT9M9/3vd4QwBRDGS9iNNX1ZH9pZHKBjGpilsBAhQRVYIjeV5/C9y8VjVU7kvgSFJy5qnZMGE
lnELcksUruO/1HvLpp1rya78j2bypfIIhSTtEnp5o+IKwCKClRYC8S0tijYaAHb8dpy2zK1bNoGG
cD/tGYos2iJOQJK4KmBTtIDjUMZEzBltOAdtlCAFJRG15uclqNCAqb2ReZiw7jqnFAdsLclH7vEv
2H3PdCT9PY+mp8TdU1xpcr9aknvmJd7KSXwehLB7ObZnFZgNG3JqN/p9VL1nCoO8F1heXKbuOTh4
1oQaEgGv7tGug62QYNOqj9gAA3whNJC6Dyj9egqERP4pEExiguMyl8ZIFbzB1dwYzUd5MuMW+qLX
t6OlLBFTrbhaaK8wfaz4HsgnmQ5t6Kv5WkV4AslIs5acwF16vtM7UHA3KTPcXScXotBLpPCAPf1W
mK/fRv2S+yW/2If0wVGmb2LcqpFEsxeRQR4+RwJMZ3ciFtNqVYHHrQaOhqwwb5ua5szyNAi/pDIT
fVUV7R6YMnQyBaz025AXQ6+mcSaLROf17xzBt7DLwHePulSSryG13tAbChvGMMjQT37f/qpvFqYj
+sLYxREVrSJgk7epx7OfKVk33xebzmiW4cYiwdm4cuaYchx6rIJvjpKIKUuVySz5OIdL+NcQAHD4
5SB4+1toE5kA3BDQBGe8AZJ2l376E0wtcBmlVO7slI4W5NcGwBBl5Q8NLngPhafFR5QPeUYsUrxj
yn9U/NfjdDRiLh6Vg4j1yR2NE+vllVss73SRsI2FTaUhcPPFu+awVCkpGqId9DSLaU9OHhqIwoS1
B2KHJEi2jSqCZDF9C0T3tCwTG4u3MUu+C9Cb7n1wev1CG6s6yq4Ahw1mcgjlu5LmaLkgvFXD53Si
I3VXwZADDhZ4KgQSZFNMAokioVF2A93lWBvLjNQmx6P9+vZvGaaYagUUwwz/yY2fhEr9nxcMq1dR
OSFSuYWpQCL/nMOU7Cx1SCbQLMENa4XhUjQdQE/3FVFUrqg/VM5D6n8dHXqezw22WUZI90AmIB6A
tdgwnCTm69uOlFaWGYY4hhnSnxWGZgs+tj83ADcKM4Z2WuvnZryDjzE1F04Q5zY9WCgpb4uCPmWH
kSmHEZWgSr6YnObY/xTlvupP/jgmwpiKfEgTFSdAILvQBjrBwtQ88GEZZCXxuf36nZOT7y9WmF4R
aYc79l73ST5o2ilYOkp4po761dU6II4Raua3qZaLDyxarHEEwvnGNxhyVhwbwwVaUFsEfh+XplhV
bwzRxJo9GryJVIk8x9llsfR3XmnOI47BnKazr6sirdSsNIlItOk3tgsNmTCerIpo4vIA5Sf2tDJm
stOizopkpmDamJb3KhSOAyhhJlFs4v9O15VexOX18PGNDOjpncKNmClIOP4F3ulViswO6E6sM3b/
LJyNcY/kjZ3d4ebI6WhAfUCuqyOJJiZsyephmPa9rZCMb3Tk5xkdaHUirIBQL14KMmAQVQK5qtHm
zDHG0YfqpfK/3aow9SwCGCU9mcl+upXh36MKFIeUSfR9Jtlx3JtR8/rlmu7qVoxcDiosL+AAn7Cb
JSToUZW/jdQC/abX49ig1Omwe7fHSPK9I7J2EdiM8/7wT0MYcKBZY15Ca6vGig0aP1EkIojhUCd8
wuvXLb8mLyXbFCOe2c6IdCw/XtFdw45tnSJ8ecfctPkUuJGXVK+cWfLN6F4V1djsU/vPuFrewsOS
mEYq4rO/kFEFBRfOIf7j6PN8T3zbS+q+W8awd5oAET74dr7lQ672UHki7uGaKXTBW/h8niEOU+Nq
nfa3KvUtGQhuC/2phKvzcXHv9wVl5uVhk6VCksiUZkZ3OnJBkpGoSDM3u6rZ2Z64EwCRGNVAnmaR
Ay5qpHNIyUYEjC/MZKTdbHrWiUZ7VDbRnE/iIow9OOMCN1V3CH9ql5QmbLDR3dwFcp83RZ7QPqqR
HMFN2rO8T//VKHZl3Je3GapmIEK10ogDgL1A/aVIZyXZ87Axm6j4FlzbmLGZyH0in5CyNwxXf0WO
W7AAbF/Nl9FgPVgEPzlztMGuMcvddsdM2voOOIlXdhETznmyVMog+MgS/vdu1H4CWJgJIAKAZnPX
0fcgiwVSq53qIfQQV1MZGhmIT6AzCLXoAbDZ2JHK0EBfuLiJfebX1DC4SdFrByPEOACD/rqH/nSO
eSIMCtpT7sURFQ4fVuCxTUo5IKNtfUVAMtZOT+nIdlwAOyPhe07QJS9jaSKFJbFLeAHD1wkrUMkB
GWxQJfpbhPXhFQICj//hBuZZcpEN59WS6ugFO4x8c2IgpKEKh4DL3PA3XiZ1ErEnvqayJ88Byxn7
7Ms49Pk/7wiROawF3zJEtmhs1WkshkhMDaEb4uXnzQcXrRhjAOHhdr+PJlxf7PVj3rNplkdC89hI
hAA8EhaTXxIZ4SwBhOZ/gnMaad66rpsZ6QGUTaBi499PkX1+zfRIa47WXD3y1ernADUOwOwxj3h2
L6pU1V79T4fmg8wvh4VFtLPofvflfKtCZu2JxRvh0MPcP63Q0K2hf9YS3yPlL0TqYeLyS6Q30fcY
JVayNG6IfUruaK/oiuqJ/0xmixAWKn7pLLBConiBfmm9qTYC7Y4LtETJ4ZRLLBZsJFTAK6uDbXx9
SxYEFJZVNceosv3IAuCHGOF0qIukJ6yLipfAKwqkWy8FCrvHQLiv1Wry+p6fizfWoRRynjcga41X
4G08k9frHSHwWmEK0K6ybO2Uaq0wXPiGotgmgUxiDCq4JBDdGjOZVh1+4Yer9ivojzv7U5IzqIFV
JqZUE/Lw+RMYJxMG2zOfrs5LCgvCBJvVREonaSpIvD07NCmPz3fWlCacgaeXSU3U3NheM9QsTiXT
VbutBhKY5p1o37sByvmDV/9iJp0vCw4/ggygs2M11WZmw4pMJPI/pWj0Vee867wluCmGp+9YUQba
Hr5qElTJcAqzv4UEa3PIxeSP4QWBBtbwBV8osrMbG99cqWuBQoVlR73Qp0KaSdIHJIl8VnAKR6ay
e8cr5WOov6yv/TP5Xe6DA74lZcYd5h9eztuZDUOA4cTFA1jJVcjuSHWEs2M2SQ==
`protect end_protected
