`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iX1WH6lCwGPTfoT4q/xNrK1Aj2reaQarfseiUAS/ifZXhEwoB6oE2D6RZAFaF0LKNSam6Ru10gWw
5pLuKoROIQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bARjz+rQAsd4I8CGYLjXNRkBYuWKzzuB9PMbJDCJ04njXAjtXL/+6vyr+nxazh3VyCYSnkr5TJI7
Ve5ZLr6quqhg31JXTykN7hQnYHCd9kyM7r0OxtPDQ1LBVhMXDkYfsb9It5sObCsIyuqLphQn9OPb
TnXAYHH1Blz3OHUzqJg=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uhPlqy3xo1NihYW65X7CDC709m7cEaomoqflzTMuS/8WBbp6sRi4syCpke34NLfAuO5W2qaz0R6K
WEYPH+EiH235nzNLMA8J24xu5dT9joybYah3TPZ0DYhTF75c6itxyHJIMV1xl+556A7yxyTqF8zi
s7XwcSTxQDJDiuMSoCU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Eb4QcmBeu+Cl8swJPx7VDsvjSfEWrnkHhWG4rWRwsc73fhQAQLplR4cWpWgTSreaLZ4C48JupiM9
B2hgDC4DJky8pusJSDf2FgZJphdDMwHLGDGbvr4ojVfULIp5wq91+a0GQnWhNlTKEmY5lBkY/P4n
7kf1Z9mEwremI8vQ2FD1+UlD5xKMI9lLLJVag6NZ1YkXBsVJcDVAo6BFDwhoEk09WbjqU65vcpB7
TL8fY7vF4lLCxbhnxZdd/P8p5EcddQnV5zhwTDPiVunMZ3hX4XFz2AQeYuapAnELVOwngFw/ukl/
7rL9ZrqYTxZjst53Sx3KBWP8KZxhzQUaTCr+vQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CVMWmA316JheGpWyNHL/MR7hELV6yopB7vREjYADDQToPcmx+apIakfQlTn+lUhbK8TYawVFWrMW
8PVl9nMkWkYU6XADi6k34a09IpJNL/zeeeR9RCXkOOAFO6i0pT+HWPb/mM+mAEusd4sZJFgErDAW
5nJsfDAJaDxrOASWGYFYEhQkMoNA7UNtmA6oAGI4jfWX94mAA3Zr5lTvq25xDQ9oyKTdcZCIpiiC
Olb288Irph+QJBryAyW6n8zFiZg9eG8BRH7elDSTqTNXP1pu2v2r6L/uBeSc84gGz+5wZijOYm5p
fh3s11Kcsikk8/7ECM//T89z/v2tqdQKtlsxmA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mTHmFURTiwMZxNH+DQsg+aX9Oa+gLa+goHbf9Wxe/MlyJHwoCuP3Q5v/Q77VpR/j1dlxGRKVGWYa
yxG6QgffcjhepHu/PcrwyyCoKhWjCNM5zi+Ot4+wTUhVBVdEJiP6WaXp4cnaIemA+otZGCMu2sX3
qnsAP9E78Xd/i7bWf42AAREfamnrdHKEIM0h7CWavLUaIZNnqa4lk91Uu7RPd225C5Psd9JD95vP
eu4FnUKLoOlr5PEsChnJwV4j2zhf9hh3PLsVUF/pW0oC6mECK5kHdByNct7cUUWMPn5vvIYimb3+
5AT2S53HD36AKdsgk5tHDf9csmg0fD3RLMSzNw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4032)
`protect data_block
/szp2oV7ktTa9Pb86zLCM3Q9zWV5CmdfEmzwXwgG1w7Yt2gBE/CAlXNOrMC/NiBkJm2Orivp8b3P
cTUkeiWE2t+dK/VR+bg+S5Ch+5soFd9mjwKv0L9QZyw0v4CPGbOzU4lt8RYdyTEPJGq1/VIB9Qld
tuj75igt9YcVgKhsH8ggRfqnghf2fWMilzLKcSACsMOu5JUyGZpceEQQ8icwtSZ//fHIYReZb8LD
ph6/WiUPRjgg85rCPxFJ2N11Wk08dxsDByqnru+yP2D9D8Q+kVyvxmHgRQIAkflppVrHd39dwxmf
bS8BvK2iZ9EDQsuthss90PZi4JvwgxFDLNJDz7H9QMna2L6qQo1IAOKfDITsRWG8KKHEc52rXHmS
j5/FWb9ybK4aTIduvIUCkTG+2uXSfGCSmp5ugLxpvWSYOdjLa87WMlpcxR0WFmCENNmOAvr8/x+U
LzpZO5hXBMoP+g4u9Ih3y7cYY2Fz8ftJAyyN7i/xEC3gPwxPWUDqewSq0iCMdNn2gYDoSZJhiF19
Z8YG6lZcIIzKGxovspYG+nWO1DbceQchk0YBnM+3uY2sUST8R05tBMm7Kvmb5m0ioG1FJ3fH9oBU
WKSqYoQHczCr0Rd69TkwxciU+VyLdhyhC/d0mSfVtO6pkWKUc+2O/E+VjTqma043PzpYOXTbjATJ
TkkiD2q4GmRPtKnKJHGqO20PmLwFJycMIvILa2hjeUsvd9Rnp9dpQVtDW6Rj4FXox7tM/70k010M
3yz8aWjicBWnuC68FXp071/J+BXaPFBhHoc6b0RzXe9ILJOeI6YtGozNeSfBIw+KOz9tt80t0IlI
E0OtSp0dPMYyr7QlzaHTLZ8Ut7AG8ubKrI6ocnpJUbha4mMNOGpbU3wo5jKRySKBeKmF227D8LZf
moGO8T9xLQbM/1siKovu9d5IBjUJOL9uUU/ooHHXPNIQrOntRp4Ci6Mynq8m/cwQVWUddooBofGV
AwbyYSpGrBlT2brY2F8z/x5WVEZ6gmp7Ri6dI8xBX9JzrKLuY+izWJ+Tx9jYjPlbrvG32JVZyajT
i5u61UpaT8PRLu/ph8mpGRJJEIBoetg7V7kXmIDUXSjc39iZiRKkvLbKL/1bQRMx4U0f72YTZgeS
24Ll04sxa7zprL0QTexfDaywXbjWxfp8TmT1P3DOCUKvPkqKjWsOi4jJw5u/5QYRL7Q/xXNhw5wa
pBmXzricvF5C5LKhRTG6EeCng+LiVCpdDXaeugV117XxoKvIF6n06uM7j0ZPB5+MF3ewu1KDPsTg
hBJebYsLe94ygDfEmWhP+eO3580eRFqjbZy+C8MOLOaUIy3Kl5FQsEM1jtVzU/XfTs1QD9DZqTxG
+pSGoWKjgVZ7VEt9VNX/F8gO5mthcRTK8bm4r+f2ebZJp4rqaXq4sBPCqTMI1eJn2JB188f0cfK1
MzSEGPBn81EWC306H3xq9a8BSS0X6i2mCSkou/eRclXmM3/TNr7p1KuDpmAMTRDsyjJGr8afkdI3
bNDBBnnRPfNGzNYwPHzn6mnbcLeeSKa2drCE9fqBo2i0O7owzs4t9EiY+KkdoJ2F7RgztMyFjcdr
KDAcKNbXLaHDMHZUmoXNEXswOYPzXl5rEc428midkOAb6KAslYvkQcRl6wD7udPzclVMvOOfpGKN
pjrMgFQb2wgJqQ0uXBhVeHFy4r/e+r+xzN7lgQRiv+gz0qoVgyUIT6mymI1S2vYkE2jdT3kGdz28
Kl9sFXtxFjs3YRbez85ofJKvVHvgGjmO/Ogb3PKBNKNXqIiVDRRBFpkYA+DtRGTvLZsw82l8tnTZ
zgHWG0DvXVYVoH73+BjL2bv4bv3326N9lLJKYRWSj2LyY3DaUzgifGRr6kWeRtxLHyXGs/Ie49Rd
dWaIF4kfVwbwLWxzJAsI0sBxB9PWHq5EI9E74KZ8B1pVLsx65/8jGetaAp/Xfykfvw5VnCeox4qx
Nyino2Yh+VuRE+RR/8+JcNC2p+hUwRiwD4V+XR/GMrkqxvAuqo0LB74+XPgI4jRzGEAzrk2pxOR3
GBdG80xJ5ZwQ/aCKBIyyvoKtNcjTv19WbBJcpJxK3n9bbcDtxMGWlNhq+Gb/pHLCs0Z7GJne+HOr
z/wyhWQI3Q1J0qw6bVQRbLS60l+bWwtJ7s1PIFO3bnOt4ohRJxWgX06sbAoYb1VSWcaWoVrTRzDK
Kgmw1A0F8YdW/3npQ3Eu/CoFLR4xVU4YYZ5mREJJS+sVE9I/CIfvvUzarB8EZ2qAKCZzEYaD/kjL
JtMnhKdGckrdQwhlC1niHMyyViMG9ke62Kh5AdCnMuiJAAVrsp8ktAmN6lTIi5pwXI6pGCRrKrwQ
v5RnbA9bT675EmePIC/fudAxY5W1QVvLG5r1PVzLO4bwc6b8qm4zkHHF9tJA/pOY4jRYgdpK2PsS
J+VlwscJpfjtr0PMhfIKPG23ITP1PA9jaZwl/Biv4skwEAKBWVzxCHVoOBklicB9uYY96T6qN41/
bJ9LL5O64V36J607DfhAnrCNH7jLuhln1jq5reHPxV/gtUdf3Wy8k/+qKMNdhKgWbC81Ygz5JnPY
fFFTs/HrXjyi9ILtNuoief8MlDHB1lo/NiDyKCCJlW+yYkAzxM3xx0zl65B9sQQfL5nVp/YTlzF6
fMFK4uKSDjezxvh5hJJqHuGqilSUQeX9Trx9SqZELVZqvxpANpG+laqtFMj0Csn8o2cs9dVk2Quk
U3ne/hZNklxZTJ0r4qQYNXvEzcyHlRv4uf5owb3OjIfXnjAFAc2I7ADOGgFkzDLc0by1Kj7+n9Li
HWJ2kluYSZvKSUIPiF3qfMG62cvTx2c20Czpo63jF0CLEfqi2sKYPLb2syl27uNdhLx2US7ppqew
hpb2CkW1TUxLZnHUWi+MemjzoCTPCYtUUDXo+3YlFtuIogDEsE0HzRz+KVF46t5PK3ROKkWZv1IE
sloN8idZmFiagWsz7FKX2MDhX5eQDgW+rITuAGtPEqJJD2l7ohftOR5p1rQVf6OxclFtPpkxsApO
M4fwoTde0GAgW0VDux58ZhiDZ8QP96Y9t7q6RJG5EiiaODgJReo9tnbVtT2sspaP8RMzvIEv7Xen
mhHM52ZW3srt8SLNeM4fDISMlM/w0bLGuQRkp4BtgsbfVsupjyYuxmlAhBkgvIpTE+ajVF0ECqgU
gQi4zDIlWPidGKYMuriD0NAduFRHYWlKAt9fBUVm7+vEEYbcUWg+d+gQow15KMjLL6AVyJXx93fR
MFtsUoBCuaHZ+6/SNB/8tiPnvwNvdj5Eho7zsWlOEdm6tIWhUfDSxjepKOLNKIEeReV/Ha34QM6R
pCy4uLSLyv1vZPLui/y1M3ecJ1ufYmdPrwKdBzLryUVgqDezFyvc2OKR2CwKMq9xi6mQnz5PNrBE
BwrohnNRVkwlCx82NZLEdu80OY18BomVXYofYrzn7FR7JE9zoX6koMnbIeO6TbsBRlirHS+7APmN
pggE6K6RbOgFvmw9SYzCkID8iFpHKgYhyjBpWdB332yBW1eA9Vl2coKWCb8Gd1ceDRBcXQteMGoh
DdZHitmfuc6hA+TQ80ZY12fG1cuOGqEKhLIPPJNdaLFpTAlqgwDHP3HD6S9i0vGbhk/GGPC8J+e8
RGD2Y8ssq5GguuTDNfqTYUij56hNIbyIThB4efQZI4CoYzwM+bNDqHQ1fADEutkzMsI6JnUIxE5j
1OjhR8LGX0hjM+QRmF3msTKj5F6r+EmostCrzPea+HZtyrfS+0o40wKZgodfj5yxIBhctEWDsec5
vuOCUUJZ3e2CsZmZ1+iG7WUiDJDIiVNaZ/phHTKe1Uf9xYc6FnUTwXAqVO1desALCPmcp7aMsaX7
Xk62m6a+WdKIl/Gb2ya+f0vEHxhxupVoUjxuGAfSL+W4MG0oa5Jo8zMfAt+JSKItJhJHjGIvO/ca
ffT24irnvq8SXstc9LiJTIRpyjnwVKpWHspi5G6WoEArVVVtHSeC2Zo/PeI+rROiMv9HeYloVClJ
wnKqEkojI1H9ttdnvrXmH5znoquf0Qc00cacfcQaKKWVDxG8kRTEJ4yKPfUJsSUOCsANrb/8Bo7Y
x9jvwQ+O9AxY9QXNnRKvN2qQo+pMpUvRwc/UHdEcDOKjS5vWHv31ne4dO46dw9dyNS/CDAuwR6AY
NaMbmj+k5S151reMsu4LVm/BYe3UPLGiz82moIwxLXWV9Il9P+pisjCJVRv3eBCmRFpf4JQi77Lf
8gdjaE2GE677DrkuYn/PIYH/Y4DVJI0VVX9xFvRdysIxTRUcdUxvjTRsGsv+A6awBjiIokhzqfqr
W88rCGLbsHFBN15L1BybYgLmfIQ4m+xpRHynavEEu5KirtZzxDlf5Us/TBw5m4z3f6NnEZT+ixfp
1OeLK1bZXrca+5uCiWQo6DOgbQ2qdHqODrrfukspDcTT8ZU6SWHtbtKAVJowrVvnMlJ0pX9NYivn
S+P1jwfFeIOTA2y7IkKyO+gEzEbzP6WhqD+F89qgBbl6lpySc+45fAnYXjZl88AvUPwE3ol20AIp
wgi5mARVMdpPewlixL160A4KeRr7kN4ZcmF8rd4HLDihfJoWpdIt/feAqSiXPxN5MF/lswHbqy7I
BGhf6RagRSJ/I8HXTzERjwks8gDrVIFLdY7Im+TDs4s5b2YJOf4A7PiGmDpjxKxDkHPppG0ugo7q
B2B3z5ZzThh1XkuGYFV+okoKpJ+0eUb4o2tl+iZnLMSm23KCdzCY4O7AlZ8HxNweQHu5+lrhr0QS
tK1oqFvbOeHuuiIFHKw1Lpge19XexXp2KUZ5cW+EAtw7axBEYw4bOeZOoVEdT3cKe9XxrmlW0M6n
VAcz52VHkQh3rP1DdxGZ3yxHXNYnjFRcYxtLMEfLRBCTPShTEZKTNQ43eOrCGlXR7KqbqR6ma2K0
ZvCGvDkN1icHQzCL9LZWI5MHuAqibpfQcxGltkYQG5ZrnJyrBtCo0FdZLFm+7oF2yxM55upD3O4O
pcjkS6l/ZUUFfKzbG/FiyPjQ95/WpoXfE0U6s8ADkqKzVv/mzYvots5dJKRDYCCfhTgI/n4WycJh
s6VecTTqeykQ5dhB0tXvZhS2QYNM6zsF6vK67OYDrjk4wJ5MFS5r7V+U0HAxlKssarY6GJ+ukVfv
cg6vg5OqpqqlF5fLJ9OIdr1P09+97TJoWJZ1H8yIZ4UGZL26B4JC2xZKgsbfLqEo8cDYON2AlTCp
yuMzIDX8PyObFHkcNnud2vNPudIh8uhVSWwLejW1XdGagr+5FLhzZ6eHaxNnSetYOpwTOed2z9lJ
PHEKZGSDwU1T5nUPNw/xFx5ho/Csrt9so9amr/ef8xYHPpYKXjqaBygy
`protect end_protected
